magic
tech sky130B
magscale 1 2
timestamp 1717261043
<< metal1 >>
rect 40494 700952 40500 701004
rect 40552 700992 40558 701004
rect 59262 700992 59268 701004
rect 40552 700964 59268 700992
rect 40552 700952 40558 700964
rect 59262 700952 59268 700964
rect 59320 700952 59326 701004
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 137278 700312 137284 700324
rect 105504 700284 137284 700312
rect 105504 700272 105510 700284
rect 137278 700272 137284 700284
rect 137336 700272 137342 700324
rect 257338 700272 257344 700324
rect 257396 700312 257402 700324
rect 267642 700312 267648 700324
rect 257396 700284 267648 700312
rect 257396 700272 257402 700284
rect 267642 700272 267648 700284
rect 267700 700272 267706 700324
rect 348786 700272 348792 700324
rect 348844 700312 348850 700324
rect 365622 700312 365628 700324
rect 348844 700284 365628 700312
rect 348844 700272 348850 700284
rect 365622 700272 365628 700284
rect 365680 700272 365686 700324
rect 527174 700272 527180 700324
rect 527232 700312 527238 700324
rect 546494 700312 546500 700324
rect 527232 700284 546500 700312
rect 527232 700272 527238 700284
rect 546494 700272 546500 700284
rect 546552 700272 546558 700324
rect 365622 695444 365628 695496
rect 365680 695484 365686 695496
rect 371878 695484 371884 695496
rect 365680 695456 371884 695484
rect 365680 695444 365686 695456
rect 371878 695444 371884 695456
rect 371936 695444 371942 695496
rect 332502 694764 332508 694816
rect 332560 694804 332566 694816
rect 338758 694804 338764 694816
rect 332560 694776 338764 694804
rect 332560 694764 332566 694776
rect 338758 694764 338764 694776
rect 338816 694764 338822 694816
rect 247678 687896 247684 687948
rect 247736 687936 247742 687948
rect 257338 687936 257344 687948
rect 247736 687908 257344 687936
rect 247736 687896 247742 687908
rect 257338 687896 257344 687908
rect 257396 687896 257402 687948
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 55214 683176 55220 683188
rect 3476 683148 55220 683176
rect 3476 683136 3482 683148
rect 55214 683136 55220 683148
rect 55272 683176 55278 683188
rect 144178 683176 144184 683188
rect 55272 683148 144184 683176
rect 55272 683136 55278 683148
rect 144178 683136 144184 683148
rect 144236 683136 144242 683188
rect 338758 682388 338764 682440
rect 338816 682428 338822 682440
rect 358722 682428 358728 682440
rect 338816 682400 358728 682428
rect 338816 682388 338822 682400
rect 358722 682388 358728 682400
rect 358780 682388 358786 682440
rect 358722 680280 358728 680332
rect 358780 680320 358786 680332
rect 366358 680320 366364 680332
rect 358780 680292 366364 680320
rect 358780 680280 358786 680292
rect 366358 680280 366364 680292
rect 366416 680280 366422 680332
rect 244550 676132 244556 676184
rect 244608 676172 244614 676184
rect 247678 676172 247684 676184
rect 244608 676144 247684 676172
rect 244608 676132 244614 676144
rect 247678 676132 247684 676144
rect 247736 676132 247742 676184
rect 507118 670692 507124 670744
rect 507176 670732 507182 670744
rect 580166 670732 580172 670744
rect 507176 670704 580172 670732
rect 507176 670692 507182 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 232498 668584 232504 668636
rect 232556 668624 232562 668636
rect 244550 668624 244556 668636
rect 232556 668596 244556 668624
rect 232556 668584 232562 668596
rect 244550 668584 244556 668596
rect 244608 668584 244614 668636
rect 371878 664436 371884 664488
rect 371936 664476 371942 664488
rect 377398 664476 377404 664488
rect 371936 664448 377404 664476
rect 371936 664436 371942 664448
rect 377398 664436 377404 664448
rect 377456 664436 377462 664488
rect 366358 663008 366364 663060
rect 366416 663048 366422 663060
rect 382274 663048 382280 663060
rect 366416 663020 382280 663048
rect 366416 663008 366422 663020
rect 382274 663008 382280 663020
rect 382332 663008 382338 663060
rect 382274 660288 382280 660340
rect 382332 660328 382338 660340
rect 388438 660328 388444 660340
rect 382332 660300 388444 660328
rect 382332 660288 382338 660300
rect 388438 660288 388444 660300
rect 388496 660288 388502 660340
rect 137278 658180 137284 658232
rect 137336 658220 137342 658232
rect 138014 658220 138020 658232
rect 137336 658192 138020 658220
rect 137336 658180 137342 658192
rect 138014 658180 138020 658192
rect 138072 658180 138078 658232
rect 170306 658180 170312 658232
rect 170364 658220 170370 658232
rect 171134 658220 171140 658232
rect 170364 658192 171140 658220
rect 170364 658180 170370 658192
rect 171134 658180 171140 658192
rect 171192 658220 171198 658232
rect 172422 658220 172428 658232
rect 171192 658192 172428 658220
rect 171192 658180 171198 658192
rect 172422 658180 172428 658192
rect 172480 658180 172486 658232
rect 388438 658180 388444 658232
rect 388496 658220 388502 658232
rect 393958 658220 393964 658232
rect 388496 658192 393964 658220
rect 388496 658180 388502 658192
rect 393958 658180 393964 658192
rect 394016 658180 394022 658232
rect 429838 657704 429844 657756
rect 429896 657744 429902 657756
rect 478874 657744 478880 657756
rect 429896 657716 478880 657744
rect 429896 657704 429902 657716
rect 478874 657704 478880 657716
rect 478932 657704 478938 657756
rect 485590 657704 485596 657756
rect 485648 657744 485654 657756
rect 494790 657744 494796 657756
rect 485648 657716 494796 657744
rect 485648 657704 485654 657716
rect 494790 657704 494796 657716
rect 494848 657744 494854 657756
rect 510062 657744 510068 657756
rect 494848 657716 510068 657744
rect 494848 657704 494854 657716
rect 510062 657704 510068 657716
rect 510120 657704 510126 657756
rect 298738 657636 298744 657688
rect 298796 657676 298802 657688
rect 364978 657676 364984 657688
rect 298796 657648 364984 657676
rect 298796 657636 298802 657648
rect 364978 657636 364984 657648
rect 365036 657676 365042 657688
rect 512822 657676 512828 657688
rect 365036 657648 512828 657676
rect 365036 657636 365042 657648
rect 512822 657636 512828 657648
rect 512880 657636 512886 657688
rect 144178 657568 144184 657620
rect 144236 657608 144242 657620
rect 521102 657608 521108 657620
rect 144236 657580 521108 657608
rect 144236 657568 144242 657580
rect 521102 657568 521108 657580
rect 521160 657568 521166 657620
rect 141418 657500 141424 657552
rect 141476 657540 141482 657552
rect 519722 657540 519728 657552
rect 141476 657512 519728 657540
rect 141476 657500 141482 657512
rect 519722 657500 519728 657512
rect 519780 657500 519786 657552
rect 138014 657228 138020 657280
rect 138072 657268 138078 657280
rect 518342 657268 518348 657280
rect 138072 657240 518348 657268
rect 138072 657228 138078 657240
rect 518342 657228 518348 657240
rect 518400 657228 518406 657280
rect 485682 657160 485688 657212
rect 485740 657200 485746 657212
rect 507118 657200 507124 657212
rect 485740 657172 507124 657200
rect 485740 657160 485746 657172
rect 507118 657160 507124 657172
rect 507176 657160 507182 657212
rect 478874 657092 478880 657144
rect 478932 657132 478938 657144
rect 480162 657132 480168 657144
rect 478932 657104 480168 657132
rect 478932 657092 478938 657104
rect 480162 657092 480168 657104
rect 480220 657132 480226 657144
rect 511442 657132 511448 657144
rect 480220 657104 511448 657132
rect 480220 657092 480226 657104
rect 511442 657092 511448 657104
rect 511500 657092 511506 657144
rect 172422 657024 172428 657076
rect 172480 657064 172486 657076
rect 516962 657064 516968 657076
rect 172480 657036 516968 657064
rect 172480 657024 172486 657036
rect 516962 657024 516968 657036
rect 517020 657024 517026 657076
rect 528002 657024 528008 657076
rect 528060 657064 528066 657076
rect 543826 657064 543832 657076
rect 528060 657036 543832 657064
rect 528060 657024 528066 657036
rect 543826 657024 543832 657036
rect 543884 657024 543890 657076
rect 162118 656956 162124 657008
rect 162176 656996 162182 657008
rect 526622 656996 526628 657008
rect 162176 656968 526628 656996
rect 162176 656956 162182 656968
rect 526622 656956 526628 656968
rect 526680 656956 526686 657008
rect 533522 656956 533528 657008
rect 533580 656996 533586 657008
rect 547874 656996 547880 657008
rect 533580 656968 547880 656996
rect 533580 656956 533586 656968
rect 547874 656956 547880 656968
rect 547932 656956 547938 657008
rect 487062 656888 487068 656940
rect 487120 656928 487126 656940
rect 499022 656928 499028 656940
rect 487120 656900 499028 656928
rect 487120 656888 487126 656900
rect 499022 656888 499028 656900
rect 499080 656888 499086 656940
rect 539042 656888 539048 656940
rect 539100 656928 539106 656940
rect 547966 656928 547972 656940
rect 539100 656900 547972 656928
rect 539100 656888 539106 656900
rect 547966 656888 547972 656900
rect 548024 656888 548030 656940
rect 505922 655664 505928 655716
rect 505980 655704 505986 655716
rect 540330 655704 540336 655716
rect 505980 655676 540336 655704
rect 505980 655664 505986 655676
rect 540330 655664 540336 655676
rect 540388 655664 540394 655716
rect 155218 655596 155224 655648
rect 155276 655636 155282 655648
rect 525242 655636 525248 655648
rect 155276 655608 525248 655636
rect 155276 655596 155282 655608
rect 525242 655596 525248 655608
rect 525300 655596 525306 655648
rect 148318 655528 148324 655580
rect 148376 655568 148382 655580
rect 522482 655568 522488 655580
rect 148376 655540 522488 655568
rect 148376 655528 148382 655540
rect 522482 655528 522488 655540
rect 522540 655528 522546 655580
rect 151078 654440 151084 654492
rect 151136 654480 151142 654492
rect 523494 654480 523500 654492
rect 151136 654452 523500 654480
rect 151136 654440 151142 654452
rect 523494 654440 523500 654452
rect 523552 654440 523558 654492
rect 159358 648592 159364 648644
rect 159416 648632 159422 648644
rect 361942 648632 361948 648644
rect 159416 648604 361948 648632
rect 159416 648592 159422 648604
rect 361942 648592 361948 648604
rect 362000 648592 362006 648644
rect 393958 648524 393964 648576
rect 394016 648564 394022 648576
rect 397362 648564 397368 648576
rect 394016 648536 397368 648564
rect 394016 648524 394022 648536
rect 397362 648524 397368 648536
rect 397420 648524 397426 648576
rect 204898 647436 204904 647488
rect 204956 647476 204962 647488
rect 358078 647476 358084 647488
rect 204956 647448 358084 647476
rect 204956 647436 204962 647448
rect 358078 647436 358084 647448
rect 358136 647436 358142 647488
rect 202782 647368 202788 647420
rect 202840 647408 202846 647420
rect 359366 647408 359372 647420
rect 202840 647380 359372 647408
rect 202840 647368 202846 647380
rect 359366 647368 359372 647380
rect 359424 647368 359430 647420
rect 233142 647300 233148 647352
rect 233200 647340 233206 647352
rect 471238 647340 471244 647352
rect 233200 647312 471244 647340
rect 233200 647300 233206 647312
rect 471238 647300 471244 647312
rect 471296 647300 471302 647352
rect 208394 647232 208400 647284
rect 208452 647272 208458 647284
rect 468478 647272 468484 647284
rect 208452 647244 468484 647272
rect 208452 647232 208458 647244
rect 468478 647232 468484 647244
rect 468536 647232 468542 647284
rect 222838 646484 222844 646536
rect 222896 646524 222902 646536
rect 232498 646524 232504 646536
rect 222896 646496 232504 646524
rect 222896 646484 222902 646496
rect 232498 646484 232504 646496
rect 232556 646484 232562 646536
rect 212442 646008 212448 646060
rect 212500 646048 212506 646060
rect 354214 646048 354220 646060
rect 212500 646020 354220 646048
rect 212500 646008 212506 646020
rect 354214 646008 354220 646020
rect 354272 646008 354278 646060
rect 186590 645940 186596 645992
rect 186648 645980 186654 645992
rect 461762 645980 461768 645992
rect 186648 645952 461768 645980
rect 186648 645940 186654 645952
rect 461762 645940 461768 645952
rect 461820 645940 461826 645992
rect 194318 645872 194324 645924
rect 194376 645912 194382 645924
rect 471330 645912 471336 645924
rect 194376 645884 471336 645912
rect 194376 645872 194382 645884
rect 471330 645872 471336 645884
rect 471388 645872 471394 645924
rect 215294 644920 215300 644972
rect 215352 644960 215358 644972
rect 324590 644960 324596 644972
rect 215352 644932 324596 644960
rect 215352 644920 215358 644932
rect 324590 644920 324596 644932
rect 324648 644920 324654 644972
rect 231762 644852 231768 644904
rect 231820 644892 231826 644904
rect 375466 644892 375472 644904
rect 231820 644864 375472 644892
rect 231820 644852 231826 644864
rect 375466 644852 375472 644864
rect 375524 644852 375530 644904
rect 106182 644784 106188 644836
rect 106240 644824 106246 644836
rect 352926 644824 352932 644836
rect 106240 644796 352932 644824
rect 106240 644784 106246 644796
rect 352926 644784 352932 644796
rect 352984 644784 352990 644836
rect 227714 644716 227720 644768
rect 227772 644756 227778 644768
rect 480346 644756 480352 644768
rect 227772 644728 480352 644756
rect 227772 644716 227778 644728
rect 480346 644716 480352 644728
rect 480404 644716 480410 644768
rect 102134 644648 102140 644700
rect 102192 644688 102198 644700
rect 355502 644688 355508 644700
rect 102192 644660 355508 644688
rect 102192 644648 102198 644660
rect 355502 644648 355508 644660
rect 355560 644648 355566 644700
rect 397362 644648 397368 644700
rect 397420 644688 397426 644700
rect 404354 644688 404360 644700
rect 397420 644660 404360 644688
rect 397420 644648 397426 644660
rect 404354 644648 404360 644660
rect 404412 644648 404418 644700
rect 191742 644580 191748 644632
rect 191800 644620 191806 644632
rect 489362 644620 489368 644632
rect 191800 644592 489368 644620
rect 191800 644580 191806 644592
rect 489362 644580 489368 644592
rect 489420 644580 489426 644632
rect 189166 644512 189172 644564
rect 189224 644552 189230 644564
rect 488074 644552 488080 644564
rect 189224 644524 488080 644552
rect 189224 644512 189230 644524
rect 488074 644512 488080 644524
rect 488132 644512 488138 644564
rect 187878 644444 187884 644496
rect 187936 644484 187942 644496
rect 490098 644484 490104 644496
rect 187936 644456 490104 644484
rect 187936 644444 187942 644456
rect 490098 644444 490104 644456
rect 490156 644444 490162 644496
rect 377398 643696 377404 643748
rect 377456 643736 377462 643748
rect 397454 643736 397460 643748
rect 377456 643708 397460 643736
rect 377456 643696 377462 643708
rect 397454 643696 397460 643708
rect 397512 643696 397518 643748
rect 176654 643560 176660 643612
rect 176712 643600 176718 643612
rect 356790 643600 356796 643612
rect 176712 643572 356796 643600
rect 176712 643560 176718 643572
rect 356790 643560 356796 643572
rect 356848 643560 356854 643612
rect 233878 643492 233884 643544
rect 233936 643532 233942 643544
rect 486694 643532 486700 643544
rect 233936 643504 486700 643532
rect 233936 643492 233942 643504
rect 486694 643492 486700 643504
rect 486752 643492 486758 643544
rect 207014 643424 207020 643476
rect 207072 643464 207078 643476
rect 467190 643464 467196 643476
rect 207072 643436 467196 643464
rect 207072 643424 207078 643436
rect 467190 643424 467196 643436
rect 467248 643424 467254 643476
rect 88978 643356 88984 643408
rect 89036 643396 89042 643408
rect 364518 643396 364524 643408
rect 89036 643368 364524 643396
rect 89036 643356 89042 643368
rect 364518 643356 364524 643368
rect 364576 643356 364582 643408
rect 86862 643288 86868 643340
rect 86920 643328 86926 643340
rect 365806 643328 365812 643340
rect 86920 643300 365812 643328
rect 86920 643288 86926 643300
rect 365806 643288 365812 643300
rect 365864 643288 365870 643340
rect 80054 643220 80060 643272
rect 80112 643260 80118 643272
rect 367094 643260 367100 643272
rect 80112 643232 367100 643260
rect 80112 643220 80118 643232
rect 367094 643220 367100 643232
rect 367152 643220 367158 643272
rect 204162 643152 204168 643204
rect 204220 643192 204226 643204
rect 489914 643192 489920 643204
rect 204220 643164 489920 643192
rect 204220 643152 204226 643164
rect 489914 643152 489920 643164
rect 489972 643152 489978 643204
rect 179322 643084 179328 643136
rect 179380 643124 179386 643136
rect 473998 643124 474004 643136
rect 179380 643096 474004 643124
rect 179380 643084 179386 643096
rect 473998 643084 474004 643096
rect 474056 643084 474062 643136
rect 223482 642200 223488 642252
rect 223540 642240 223546 642252
rect 328454 642240 328460 642252
rect 223540 642212 328460 642240
rect 223540 642200 223546 642212
rect 328454 642200 328460 642212
rect 328512 642200 328518 642252
rect 92474 642132 92480 642184
rect 92532 642172 92538 642184
rect 342622 642172 342628 642184
rect 92532 642144 342628 642172
rect 92532 642132 92538 642144
rect 342622 642132 342628 642144
rect 342680 642132 342686 642184
rect 85482 642064 85488 642116
rect 85540 642104 85546 642116
rect 349062 642104 349068 642116
rect 85540 642076 349068 642104
rect 85540 642064 85546 642076
rect 349062 642064 349068 642076
rect 349120 642064 349126 642116
rect 179322 641996 179328 642048
rect 179380 642036 179386 642048
rect 474090 642036 474096 642048
rect 179380 642008 474096 642036
rect 179380 641996 179386 642008
rect 474090 641996 474096 642008
rect 474148 641996 474154 642048
rect 177942 641928 177948 641980
rect 178000 641968 178006 641980
rect 479426 641968 479432 641980
rect 178000 641940 479432 641968
rect 178000 641928 178006 641940
rect 479426 641928 479432 641940
rect 479484 641928 479490 641980
rect 177758 641860 177764 641912
rect 177816 641900 177822 641912
rect 488534 641900 488540 641912
rect 177816 641872 488540 641900
rect 177816 641860 177822 641872
rect 488534 641860 488540 641872
rect 488592 641860 488598 641912
rect 177850 641792 177856 641844
rect 177908 641832 177914 641844
rect 490006 641832 490012 641844
rect 177908 641804 490012 641832
rect 177908 641792 177914 641804
rect 490006 641792 490012 641804
rect 490064 641792 490070 641844
rect 249702 641724 249708 641776
rect 249760 641764 249766 641776
rect 369670 641764 369676 641776
rect 249760 641736 369676 641764
rect 249760 641724 249766 641736
rect 369670 641724 369676 641736
rect 369728 641724 369734 641776
rect 218054 640840 218060 640892
rect 218112 640880 218118 640892
rect 315574 640880 315580 640892
rect 218112 640852 315580 640880
rect 218112 640840 218118 640852
rect 315574 640840 315580 640852
rect 315632 640840 315638 640892
rect 214558 640772 214564 640824
rect 214616 640812 214622 640824
rect 320726 640812 320732 640824
rect 214616 640784 320732 640812
rect 214616 640772 214622 640784
rect 320726 640772 320732 640784
rect 320784 640772 320790 640824
rect 91094 640704 91100 640756
rect 91152 640744 91158 640756
rect 329742 640744 329748 640756
rect 91152 640716 329748 640744
rect 91152 640704 91158 640716
rect 329742 640704 329748 640716
rect 329800 640704 329806 640756
rect 230382 640636 230388 640688
rect 230440 640676 230446 640688
rect 485866 640676 485872 640688
rect 230440 640648 485872 640676
rect 230440 640636 230446 640648
rect 485866 640636 485872 640648
rect 485924 640636 485930 640688
rect 216766 640568 216772 640620
rect 216824 640608 216830 640620
rect 480438 640608 480444 640620
rect 216824 640580 480444 640608
rect 216824 640568 216830 640580
rect 480438 640568 480444 640580
rect 480496 640568 480502 640620
rect 211062 640500 211068 640552
rect 211120 640540 211126 640552
rect 488810 640540 488816 640552
rect 211120 640512 488816 640540
rect 211120 640500 211126 640512
rect 488810 640500 488816 640512
rect 488868 640500 488874 640552
rect 185670 640432 185676 640484
rect 185728 640472 185734 640484
rect 464430 640472 464436 640484
rect 185728 640444 464436 640472
rect 185728 640432 185734 640444
rect 464430 640432 464436 640444
rect 464488 640432 464494 640484
rect 190730 640364 190736 640416
rect 190788 640404 190794 640416
rect 490190 640404 490196 640416
rect 190788 640376 490196 640404
rect 190788 640364 190794 640376
rect 490190 640364 490196 640376
rect 490248 640364 490254 640416
rect 56502 640296 56508 640348
rect 56560 640336 56566 640348
rect 363230 640336 363236 640348
rect 56560 640308 363236 640336
rect 56560 640296 56566 640308
rect 363230 640296 363236 640308
rect 363288 640296 363294 640348
rect 404354 640296 404360 640348
rect 404412 640336 404418 640348
rect 410518 640336 410524 640348
rect 404412 640308 410524 640336
rect 404412 640296 404418 640308
rect 410518 640296 410524 640308
rect 410576 640296 410582 640348
rect 397454 640228 397460 640280
rect 397512 640268 397518 640280
rect 400858 640268 400864 640280
rect 397512 640240 400864 640268
rect 397512 640228 397518 640240
rect 400858 640228 400864 640240
rect 400916 640228 400922 640280
rect 220722 639548 220728 639600
rect 220780 639588 220786 639600
rect 485774 639588 485780 639600
rect 220780 639560 485780 639588
rect 220780 639548 220786 639560
rect 485774 639548 485780 639560
rect 485832 639548 485838 639600
rect 122742 639412 122748 639464
rect 122800 639452 122806 639464
rect 306558 639452 306564 639464
rect 122800 639424 306564 639452
rect 122800 639412 122806 639424
rect 306558 639412 306564 639424
rect 306616 639412 306622 639464
rect 95142 639344 95148 639396
rect 95200 639384 95206 639396
rect 318150 639384 318156 639396
rect 95200 639356 318156 639384
rect 95200 639344 95206 639356
rect 318150 639344 318156 639356
rect 318208 639344 318214 639396
rect 251082 639276 251088 639328
rect 251140 639316 251146 639328
rect 479334 639316 479340 639328
rect 251140 639288 479340 639316
rect 251140 639276 251146 639288
rect 479334 639276 479340 639288
rect 479392 639276 479398 639328
rect 82814 639208 82820 639260
rect 82872 639248 82878 639260
rect 319438 639248 319444 639260
rect 82872 639220 319444 639248
rect 82872 639208 82878 639220
rect 319438 639208 319444 639220
rect 319496 639208 319502 639260
rect 81434 639140 81440 639192
rect 81492 639180 81498 639192
rect 322014 639180 322020 639192
rect 81492 639152 322020 639180
rect 81492 639140 81498 639152
rect 322014 639140 322020 639152
rect 322072 639140 322078 639192
rect 125594 639072 125600 639124
rect 125652 639112 125658 639124
rect 376846 639112 376852 639124
rect 125652 639084 376852 639112
rect 125652 639072 125658 639084
rect 376846 639072 376852 639084
rect 376904 639072 376910 639124
rect 234614 639004 234620 639056
rect 234672 639044 234678 639056
rect 487246 639044 487252 639056
rect 234672 639016 487252 639044
rect 234672 639004 234678 639016
rect 487246 639004 487252 639016
rect 487304 639004 487310 639056
rect 58618 638936 58624 638988
rect 58676 638976 58682 638988
rect 139026 638976 139032 638988
rect 58676 638948 139032 638976
rect 58676 638936 58682 638948
rect 139026 638936 139032 638948
rect 139084 638936 139090 638988
rect 213822 638936 213828 638988
rect 213880 638976 213886 638988
rect 488626 638976 488632 638988
rect 213880 638948 488632 638976
rect 213880 638936 213886 638948
rect 488626 638936 488632 638948
rect 488684 638936 488690 638988
rect 129734 638392 129740 638444
rect 129792 638432 129798 638444
rect 283742 638432 283748 638444
rect 129792 638404 283748 638432
rect 129792 638392 129798 638404
rect 283742 638392 283748 638404
rect 283800 638392 283806 638444
rect 123478 638324 123484 638376
rect 123536 638364 123542 638376
rect 289078 638364 289084 638376
rect 123536 638336 289084 638364
rect 123536 638324 123542 638336
rect 289078 638324 289084 638336
rect 289136 638324 289142 638376
rect 278130 638256 278136 638308
rect 278188 638296 278194 638308
rect 343910 638296 343916 638308
rect 278188 638268 343916 638296
rect 278188 638256 278194 638268
rect 343910 638256 343916 638268
rect 343968 638256 343974 638308
rect 211062 638188 211068 638240
rect 211120 638228 211126 638240
rect 487154 638228 487160 638240
rect 211120 638200 487160 638228
rect 211120 638188 211126 638200
rect 487154 638188 487160 638200
rect 487212 638188 487218 638240
rect 280890 638120 280896 638172
rect 280948 638160 280954 638172
rect 346486 638160 346492 638172
rect 280948 638132 346492 638160
rect 280948 638120 280954 638132
rect 346486 638120 346492 638132
rect 346544 638120 346550 638172
rect 283558 638052 283564 638104
rect 283616 638092 283622 638104
rect 347774 638092 347780 638104
rect 283616 638064 347780 638092
rect 283616 638052 283622 638064
rect 347774 638052 347780 638064
rect 347832 638052 347838 638104
rect 110322 637984 110328 638036
rect 110380 638024 110386 638036
rect 295978 638024 295984 638036
rect 110380 637996 295984 638024
rect 110380 637984 110386 637996
rect 295978 637984 295984 637996
rect 296036 637984 296042 638036
rect 108298 637916 108304 637968
rect 108356 637956 108362 637968
rect 331030 637956 331036 637968
rect 108356 637928 331036 637956
rect 108356 637916 108362 637928
rect 331030 637916 331036 637928
rect 331088 637916 331094 637968
rect 247494 637848 247500 637900
rect 247552 637888 247558 637900
rect 488534 637888 488540 637900
rect 247552 637860 488540 637888
rect 247552 637848 247558 637860
rect 488534 637848 488540 637860
rect 488592 637848 488598 637900
rect 224218 637780 224224 637832
rect 224276 637820 224282 637832
rect 480254 637820 480260 637832
rect 224276 637792 480260 637820
rect 224276 637780 224282 637792
rect 480254 637780 480260 637792
rect 480312 637780 480318 637832
rect 230382 637712 230388 637764
rect 230440 637752 230446 637764
rect 487430 637752 487436 637764
rect 230440 637724 487436 637752
rect 230440 637712 230446 637724
rect 487430 637712 487436 637724
rect 487488 637712 487494 637764
rect 115474 637644 115480 637696
rect 115532 637684 115538 637696
rect 381538 637684 381544 637696
rect 115532 637656 381544 637684
rect 115532 637644 115538 637656
rect 381538 637644 381544 637656
rect 381596 637644 381602 637696
rect 109034 637576 109040 637628
rect 109092 637616 109098 637628
rect 375558 637616 375564 637628
rect 109092 637588 375564 637616
rect 109092 637576 109098 637588
rect 375558 637576 375564 637588
rect 375616 637576 375622 637628
rect 73154 637032 73160 637084
rect 73212 637072 73218 637084
rect 350350 637072 350356 637084
rect 73212 637044 350356 637072
rect 73212 637032 73218 637044
rect 350350 637032 350356 637044
rect 350408 637032 350414 637084
rect 241054 636964 241060 637016
rect 241112 637004 241118 637016
rect 468570 637004 468576 637016
rect 241112 636976 468576 637004
rect 241112 636964 241118 636976
rect 468570 636964 468576 636976
rect 468628 636964 468634 637016
rect 273990 636896 273996 636948
rect 274048 636936 274054 636948
rect 302694 636936 302700 636948
rect 274048 636908 302700 636936
rect 274048 636896 274054 636908
rect 302694 636896 302700 636908
rect 302752 636896 302758 636948
rect 101306 636828 101312 636880
rect 101364 636868 101370 636880
rect 135990 636868 135996 636880
rect 101364 636840 135996 636868
rect 101364 636828 101370 636840
rect 135990 636828 135996 636840
rect 136048 636828 136054 636880
rect 249610 636828 249616 636880
rect 249668 636868 249674 636880
rect 268378 636868 268384 636880
rect 249668 636840 268384 636868
rect 249668 636828 249674 636840
rect 268378 636828 268384 636840
rect 268436 636828 268442 636880
rect 279694 636828 279700 636880
rect 279752 636868 279758 636880
rect 314286 636868 314292 636880
rect 279752 636840 314292 636868
rect 279752 636828 279758 636840
rect 314286 636828 314292 636840
rect 314344 636828 314350 636880
rect 124214 636760 124220 636812
rect 124272 636800 124278 636812
rect 135898 636800 135904 636812
rect 124272 636772 135904 636800
rect 124272 636760 124278 636772
rect 135898 636760 135904 636772
rect 135956 636760 135962 636812
rect 238386 636760 238392 636812
rect 238444 636800 238450 636812
rect 271230 636800 271236 636812
rect 238444 636772 271236 636800
rect 238444 636760 238450 636772
rect 271230 636760 271236 636772
rect 271288 636760 271294 636812
rect 275370 636760 275376 636812
rect 275428 636800 275434 636812
rect 327166 636800 327172 636812
rect 275428 636772 327172 636800
rect 275428 636760 275434 636772
rect 327166 636760 327172 636772
rect 327224 636760 327230 636812
rect 99374 636692 99380 636744
rect 99432 636732 99438 636744
rect 311710 636732 311716 636744
rect 99432 636704 311716 636732
rect 99432 636692 99438 636704
rect 311710 636692 311716 636704
rect 311768 636692 311774 636744
rect 114186 636624 114192 636676
rect 114244 636664 114250 636676
rect 138658 636664 138664 636676
rect 114244 636636 138664 636664
rect 114244 636624 114250 636636
rect 138658 636624 138664 636636
rect 138716 636624 138722 636676
rect 243630 636624 243636 636676
rect 243688 636664 243694 636676
rect 465810 636664 465816 636676
rect 243688 636636 465816 636664
rect 243688 636624 243694 636636
rect 465810 636624 465816 636636
rect 465868 636624 465874 636676
rect 111610 636556 111616 636608
rect 111668 636596 111674 636608
rect 138750 636596 138756 636608
rect 111668 636568 138756 636596
rect 111668 636556 111674 636568
rect 138750 636556 138756 636568
rect 138808 636556 138814 636608
rect 239674 636556 239680 636608
rect 239732 636596 239738 636608
rect 468662 636596 468668 636608
rect 239732 636568 468668 636596
rect 239732 636556 239738 636568
rect 468662 636556 468668 636568
rect 468720 636556 468726 636608
rect 106458 636488 106464 636540
rect 106516 636528 106522 636540
rect 162302 636528 162308 636540
rect 106516 636500 162308 636528
rect 106516 636488 106522 636500
rect 162302 636488 162308 636500
rect 162360 636488 162366 636540
rect 237098 636488 237104 636540
rect 237156 636528 237162 636540
rect 468754 636528 468760 636540
rect 237156 636500 468760 636528
rect 237156 636488 237162 636500
rect 468754 636488 468760 636500
rect 468812 636488 468818 636540
rect 78582 636420 78588 636472
rect 78640 636460 78646 636472
rect 323302 636460 323308 636472
rect 78640 636432 323308 636460
rect 78640 636420 78646 636432
rect 323302 636420 323308 636432
rect 323360 636420 323366 636472
rect 75822 636352 75828 636404
rect 75880 636392 75886 636404
rect 338758 636392 338764 636404
rect 75880 636364 338764 636392
rect 75880 636352 75886 636364
rect 338758 636352 338764 636364
rect 338816 636352 338822 636404
rect 131114 636284 131120 636336
rect 131172 636324 131178 636336
rect 134702 636324 134708 636336
rect 131172 636296 134708 636324
rect 131172 636284 131178 636296
rect 134702 636284 134708 636296
rect 134760 636284 134766 636336
rect 129642 636216 129648 636268
rect 129700 636256 129706 636268
rect 249702 636256 249708 636268
rect 129700 636228 249708 636256
rect 129700 636216 129706 636228
rect 249702 636216 249708 636228
rect 249760 636216 249766 636268
rect 369670 636216 369676 636268
rect 369728 636256 369734 636268
rect 374546 636256 374552 636268
rect 369728 636228 374552 636256
rect 369728 636216 369734 636228
rect 374546 636216 374552 636228
rect 374604 636216 374610 636268
rect 79318 635672 79324 635724
rect 79376 635712 79382 635724
rect 296714 635712 296720 635724
rect 79376 635684 296720 635712
rect 79376 635672 79382 635684
rect 296714 635672 296720 635684
rect 296772 635672 296778 635724
rect 53834 635604 53840 635656
rect 53892 635644 53898 635656
rect 377030 635644 377036 635656
rect 53892 635616 377036 635644
rect 53892 635604 53898 635616
rect 377030 635604 377036 635616
rect 377088 635604 377094 635656
rect 170398 635536 170404 635588
rect 170456 635576 170462 635588
rect 222838 635576 222844 635588
rect 170456 635548 222844 635576
rect 170456 635536 170462 635548
rect 222838 635536 222844 635548
rect 222896 635536 222902 635588
rect 271138 635536 271144 635588
rect 271196 635576 271202 635588
rect 325878 635576 325884 635588
rect 271196 635548 325884 635576
rect 271196 635536 271202 635548
rect 325878 635536 325884 635548
rect 325936 635536 325942 635588
rect 39942 635468 39948 635520
rect 40000 635508 40006 635520
rect 72970 635508 72976 635520
rect 40000 635480 72976 635508
rect 40000 635468 40006 635480
rect 72970 635468 72976 635480
rect 73028 635468 73034 635520
rect 112898 635468 112904 635520
rect 112956 635508 112962 635520
rect 264238 635508 264244 635520
rect 112956 635480 264244 635508
rect 112956 635468 112962 635480
rect 264238 635468 264244 635480
rect 264296 635468 264302 635520
rect 276842 635468 276848 635520
rect 276900 635508 276906 635520
rect 337470 635508 337476 635520
rect 276900 635480 337476 635508
rect 276900 635468 276906 635480
rect 337470 635468 337476 635480
rect 337528 635468 337534 635520
rect 119982 635400 119988 635452
rect 120040 635440 120046 635452
rect 273898 635440 273904 635452
rect 120040 635412 273904 635440
rect 120040 635400 120046 635412
rect 273898 635400 273904 635412
rect 273956 635400 273962 635452
rect 274082 635400 274088 635452
rect 274140 635440 274146 635452
rect 372246 635440 372252 635452
rect 274140 635412 372252 635440
rect 274140 635400 274146 635412
rect 372246 635400 372252 635412
rect 372304 635400 372310 635452
rect 121362 635332 121368 635384
rect 121420 635372 121426 635384
rect 290458 635372 290464 635384
rect 121420 635344 290464 635372
rect 121420 635332 121426 635344
rect 290458 635332 290464 635344
rect 290516 635332 290522 635384
rect 97902 635264 97908 635316
rect 97960 635304 97966 635316
rect 297542 635304 297548 635316
rect 97960 635276 297548 635304
rect 97960 635264 97966 635276
rect 297542 635264 297548 635276
rect 297600 635264 297606 635316
rect 252462 635196 252468 635248
rect 252520 635236 252526 635248
rect 465718 635236 465724 635248
rect 252520 635208 465724 635236
rect 252520 635196 252526 635208
rect 465718 635196 465724 635208
rect 465776 635196 465782 635248
rect 289170 635128 289176 635180
rect 289228 635168 289234 635180
rect 341334 635168 341340 635180
rect 289228 635140 341340 635168
rect 289228 635128 289234 635140
rect 341334 635128 341340 635140
rect 341392 635128 341398 635180
rect 244274 635060 244280 635112
rect 244332 635100 244338 635112
rect 487338 635100 487344 635112
rect 244332 635072 487344 635100
rect 244332 635060 244338 635072
rect 487338 635060 487344 635072
rect 487396 635060 487402 635112
rect 226334 634992 226340 635044
rect 226392 635032 226398 635044
rect 476758 635032 476764 635044
rect 226392 635004 476764 635032
rect 226392 634992 226398 635004
rect 476758 634992 476764 635004
rect 476816 634992 476822 635044
rect 71866 634924 71872 634976
rect 71924 634964 71930 634976
rect 377214 634964 377220 634976
rect 71924 634936 377220 634964
rect 71924 634924 71930 634936
rect 377214 634924 377220 634936
rect 377272 634924 377278 634976
rect 70578 634856 70584 634908
rect 70636 634896 70642 634908
rect 377122 634896 377128 634908
rect 70636 634868 377128 634896
rect 70636 634856 70642 634868
rect 377122 634856 377128 634868
rect 377180 634856 377186 634908
rect 246114 634788 246120 634840
rect 246172 634828 246178 634840
rect 265618 634828 265624 634840
rect 246172 634800 265624 634828
rect 246172 634788 246178 634800
rect 265618 634788 265624 634800
rect 265676 634788 265682 634840
rect 286410 634584 286416 634636
rect 286468 634624 286474 634636
rect 312630 634624 312636 634636
rect 286468 634596 312636 634624
rect 286468 634584 286474 634596
rect 312630 634584 312636 634596
rect 312688 634584 312694 634636
rect 284938 634516 284944 634568
rect 284996 634556 285002 634568
rect 307662 634556 307668 634568
rect 284996 634528 307668 634556
rect 284996 634516 285002 634528
rect 307662 634516 307668 634528
rect 307720 634516 307726 634568
rect 274174 634448 274180 634500
rect 274232 634488 274238 634500
rect 316494 634488 316500 634500
rect 274232 634460 316500 634488
rect 274232 634448 274238 634460
rect 316494 634448 316500 634460
rect 316552 634448 316558 634500
rect 129826 634380 129832 634432
rect 129884 634420 129890 634432
rect 297174 634420 297180 634432
rect 129884 634392 297180 634420
rect 129884 634380 129890 634392
rect 297174 634380 297180 634392
rect 297232 634380 297238 634432
rect 139026 633360 139032 633412
rect 139084 633400 139090 633412
rect 148318 633400 148324 633412
rect 139084 633372 148324 633400
rect 139084 633360 139090 633372
rect 148318 633360 148324 633372
rect 148376 633360 148382 633412
rect 3418 632680 3424 632732
rect 3476 632720 3482 632732
rect 55582 632720 55588 632732
rect 3476 632692 55588 632720
rect 3476 632680 3482 632692
rect 55582 632680 55588 632692
rect 55640 632680 55646 632732
rect 374546 632680 374552 632732
rect 374604 632720 374610 632732
rect 453298 632720 453304 632732
rect 374604 632692 453304 632720
rect 374604 632680 374610 632692
rect 453298 632680 453304 632692
rect 453356 632680 453362 632732
rect 410518 632000 410524 632052
rect 410576 632040 410582 632052
rect 413278 632040 413284 632052
rect 410576 632012 413284 632040
rect 410576 632000 410582 632012
rect 413278 632000 413284 632012
rect 413336 632000 413342 632052
rect 377674 625540 377680 625592
rect 377732 625580 377738 625592
rect 380986 625580 380992 625592
rect 377732 625552 380992 625580
rect 377732 625540 377738 625552
rect 380986 625540 380992 625552
rect 381044 625540 381050 625592
rect 377674 623772 377680 623824
rect 377732 623812 377738 623824
rect 381078 623812 381084 623824
rect 377732 623784 381084 623812
rect 377732 623772 377738 623784
rect 381078 623772 381084 623784
rect 381136 623772 381142 623824
rect 164970 622412 164976 622464
rect 165028 622452 165034 622464
rect 170398 622452 170404 622464
rect 165028 622424 170404 622452
rect 165028 622412 165034 622424
rect 170398 622412 170404 622424
rect 170456 622412 170462 622464
rect 377766 622412 377772 622464
rect 377824 622452 377830 622464
rect 381170 622452 381176 622464
rect 377824 622424 381176 622452
rect 377824 622412 377830 622424
rect 381170 622412 381176 622424
rect 381228 622412 381234 622464
rect 377030 620984 377036 621036
rect 377088 621024 377094 621036
rect 379514 621024 379520 621036
rect 377088 620996 379520 621024
rect 377088 620984 377094 620996
rect 379514 620984 379520 620996
rect 379572 620984 379578 621036
rect 400858 617516 400864 617568
rect 400916 617556 400922 617568
rect 426342 617556 426348 617568
rect 400916 617528 426348 617556
rect 400916 617516 400922 617528
rect 426342 617516 426348 617528
rect 426400 617516 426406 617568
rect 540330 617516 540336 617568
rect 540388 617556 540394 617568
rect 580166 617556 580172 617568
rect 540388 617528 580172 617556
rect 540388 617516 540394 617528
rect 580166 617516 580172 617528
rect 580224 617516 580230 617568
rect 283650 614116 283656 614168
rect 283708 614156 283714 614168
rect 298002 614156 298008 614168
rect 283708 614128 298008 614156
rect 283708 614116 283714 614128
rect 298002 614116 298008 614128
rect 298060 614116 298066 614168
rect 453298 613368 453304 613420
rect 453356 613408 453362 613420
rect 477494 613408 477500 613420
rect 453356 613380 477500 613408
rect 453356 613368 453362 613380
rect 477494 613368 477500 613380
rect 477552 613368 477558 613420
rect 413278 612756 413284 612808
rect 413336 612796 413342 612808
rect 416038 612796 416044 612808
rect 413336 612768 416044 612796
rect 413336 612756 413342 612768
rect 416038 612756 416044 612768
rect 416096 612756 416102 612808
rect 477494 612756 477500 612808
rect 477552 612796 477558 612808
rect 478782 612796 478788 612808
rect 477552 612768 478788 612796
rect 477552 612756 477558 612768
rect 478782 612756 478788 612768
rect 478840 612796 478846 612808
rect 487154 612796 487160 612808
rect 478840 612768 487160 612796
rect 478840 612756 478846 612768
rect 487154 612756 487160 612768
rect 487212 612756 487218 612808
rect 159542 612008 159548 612060
rect 159600 612048 159606 612060
rect 164970 612048 164976 612060
rect 159600 612020 164976 612048
rect 159600 612008 159606 612020
rect 164970 612008 164976 612020
rect 165028 612008 165034 612060
rect 289354 611328 289360 611380
rect 289412 611368 289418 611380
rect 298002 611368 298008 611380
rect 289412 611340 298008 611368
rect 289412 611328 289418 611340
rect 298002 611328 298008 611340
rect 298060 611328 298066 611380
rect 283834 609968 283840 610020
rect 283892 610008 283898 610020
rect 298002 610008 298008 610020
rect 283892 609980 298008 610008
rect 283892 609968 283898 609980
rect 298002 609968 298008 609980
rect 298060 609968 298066 610020
rect 426342 609220 426348 609272
rect 426400 609260 426406 609272
rect 442258 609260 442264 609272
rect 426400 609232 442264 609260
rect 426400 609220 426406 609232
rect 442258 609220 442264 609232
rect 442316 609220 442322 609272
rect 378042 605820 378048 605872
rect 378100 605860 378106 605872
rect 385034 605860 385040 605872
rect 378100 605832 385040 605860
rect 378100 605820 378106 605832
rect 385034 605820 385040 605832
rect 385092 605820 385098 605872
rect 378042 604528 378048 604580
rect 378100 604568 378106 604580
rect 386414 604568 386420 604580
rect 378100 604540 386420 604568
rect 378100 604528 378106 604540
rect 386414 604528 386420 604540
rect 386472 604528 386478 604580
rect 377950 604460 377956 604512
rect 378008 604500 378014 604512
rect 389174 604500 389180 604512
rect 378008 604472 389180 604500
rect 378008 604460 378014 604472
rect 389174 604460 389180 604472
rect 389232 604460 389238 604512
rect 378042 603236 378048 603288
rect 378100 603276 378106 603288
rect 385126 603276 385132 603288
rect 378100 603248 385132 603276
rect 378100 603236 378106 603248
rect 385126 603236 385132 603248
rect 385184 603236 385190 603288
rect 378042 603100 378048 603152
rect 378100 603140 378106 603152
rect 386598 603140 386604 603152
rect 378100 603112 386604 603140
rect 378100 603100 378106 603112
rect 386598 603100 386604 603112
rect 386656 603100 386662 603152
rect 538582 600584 538588 600636
rect 538640 600624 538646 600636
rect 539318 600624 539324 600636
rect 538640 600596 539324 600624
rect 538640 600584 538646 600596
rect 539318 600584 539324 600596
rect 539376 600584 539382 600636
rect 535730 600244 535736 600296
rect 535788 600284 535794 600296
rect 542630 600284 542636 600296
rect 535788 600256 542636 600284
rect 535788 600244 535794 600256
rect 542630 600244 542636 600256
rect 542688 600244 542694 600296
rect 536834 600176 536840 600228
rect 536892 600216 536898 600228
rect 542722 600216 542728 600228
rect 536892 600188 542728 600216
rect 536892 600176 536898 600188
rect 542722 600176 542728 600188
rect 542780 600176 542786 600228
rect 534718 600108 534724 600160
rect 534776 600148 534782 600160
rect 540330 600148 540336 600160
rect 534776 600120 540336 600148
rect 534776 600108 534782 600120
rect 540330 600108 540336 600120
rect 540388 600108 540394 600160
rect 487062 599700 487068 599752
rect 487120 599740 487126 599752
rect 498194 599740 498200 599752
rect 487120 599712 498200 599740
rect 487120 599700 487126 599712
rect 498194 599700 498200 599712
rect 498252 599700 498258 599752
rect 485590 599632 485596 599684
rect 485648 599672 485654 599684
rect 505094 599672 505100 599684
rect 485648 599644 505100 599672
rect 485648 599632 485654 599644
rect 505094 599632 505100 599644
rect 505152 599632 505158 599684
rect 485682 599564 485688 599616
rect 485740 599604 485746 599616
rect 506474 599604 506480 599616
rect 485740 599576 506480 599604
rect 485740 599564 485746 599576
rect 506474 599564 506480 599576
rect 506532 599564 506538 599616
rect 502978 598204 502984 598256
rect 503036 598244 503042 598256
rect 539042 598244 539048 598256
rect 503036 598216 539048 598244
rect 503036 598204 503042 598216
rect 539042 598204 539048 598216
rect 539100 598204 539106 598256
rect 157058 597456 157064 597508
rect 157116 597496 157122 597508
rect 159542 597496 159548 597508
rect 157116 597468 159548 597496
rect 157116 597456 157122 597468
rect 159542 597456 159548 597468
rect 159600 597456 159606 597508
rect 47946 594804 47952 594856
rect 48004 594844 48010 594856
rect 56962 594844 56968 594856
rect 48004 594816 56968 594844
rect 48004 594804 48010 594816
rect 56962 594804 56968 594816
rect 57020 594804 57026 594856
rect 285306 594804 285312 594856
rect 285364 594844 285370 594856
rect 298002 594844 298008 594856
rect 285364 594816 298008 594844
rect 285364 594804 285370 594816
rect 298002 594804 298008 594816
rect 298060 594804 298066 594856
rect 378042 594804 378048 594856
rect 378100 594844 378106 594856
rect 385218 594844 385224 594856
rect 378100 594816 385224 594844
rect 378100 594804 378106 594816
rect 385218 594804 385224 594816
rect 385276 594804 385282 594856
rect 442258 594804 442264 594856
rect 442316 594844 442322 594856
rect 448514 594844 448520 594856
rect 442316 594816 448520 594844
rect 442316 594804 442322 594816
rect 448514 594804 448520 594816
rect 448572 594804 448578 594856
rect 147398 594056 147404 594108
rect 147456 594096 147462 594108
rect 157058 594096 157064 594108
rect 147456 594068 157064 594096
rect 147456 594056 147462 594068
rect 157058 594056 157064 594068
rect 157116 594056 157122 594108
rect 378042 592084 378048 592136
rect 378100 592124 378106 592136
rect 383654 592124 383660 592136
rect 378100 592096 383660 592124
rect 378100 592084 378106 592096
rect 383654 592084 383660 592096
rect 383712 592084 383718 592136
rect 377950 592016 377956 592068
rect 378008 592056 378014 592068
rect 386690 592056 386696 592068
rect 378008 592028 386696 592056
rect 378008 592016 378014 592028
rect 386690 592016 386696 592028
rect 386748 592016 386754 592068
rect 448514 591268 448520 591320
rect 448572 591308 448578 591320
rect 454678 591308 454684 591320
rect 448572 591280 454684 591308
rect 448572 591268 448578 591280
rect 454678 591268 454684 591280
rect 454736 591268 454742 591320
rect 50614 590656 50620 590708
rect 50672 590696 50678 590708
rect 56962 590696 56968 590708
rect 50672 590668 56968 590696
rect 50672 590656 50678 590668
rect 56962 590656 56968 590668
rect 57020 590656 57026 590708
rect 144270 590656 144276 590708
rect 144328 590696 144334 590708
rect 147398 590696 147404 590708
rect 144328 590668 147404 590696
rect 144328 590656 144334 590668
rect 147398 590656 147404 590668
rect 147456 590656 147462 590708
rect 288158 590656 288164 590708
rect 288216 590696 288222 590708
rect 298002 590696 298008 590708
rect 288216 590668 298008 590696
rect 288216 590656 288222 590668
rect 298002 590656 298008 590668
rect 298060 590656 298066 590708
rect 378042 590656 378048 590708
rect 378100 590696 378106 590708
rect 385402 590696 385408 590708
rect 378100 590668 385408 590696
rect 378100 590656 378106 590668
rect 385402 590656 385408 590668
rect 385460 590656 385466 590708
rect 378042 589636 378048 589688
rect 378100 589676 378106 589688
rect 385310 589676 385316 589688
rect 378100 589648 385316 589676
rect 378100 589636 378106 589648
rect 385310 589636 385316 589648
rect 385368 589636 385374 589688
rect 53374 589500 53380 589552
rect 53432 589540 53438 589552
rect 56962 589540 56968 589552
rect 53432 589512 56968 589540
rect 53432 589500 53438 589512
rect 56962 589500 56968 589512
rect 57020 589500 57026 589552
rect 378042 587936 378048 587988
rect 378100 587976 378106 587988
rect 382642 587976 382648 587988
rect 378100 587948 382648 587976
rect 378100 587936 378106 587948
rect 382642 587936 382648 587948
rect 382700 587936 382706 587988
rect 377030 587868 377036 587920
rect 377088 587908 377094 587920
rect 379790 587908 379796 587920
rect 377088 587880 379796 587908
rect 377088 587868 377094 587880
rect 379790 587868 379796 587880
rect 379848 587868 379854 587920
rect 377858 587052 377864 587104
rect 377916 587092 377922 587104
rect 381446 587092 381452 587104
rect 377916 587064 381452 587092
rect 377916 587052 377922 587064
rect 381446 587052 381452 587064
rect 381504 587052 381510 587104
rect 377858 586644 377864 586696
rect 377916 586684 377922 586696
rect 381354 586684 381360 586696
rect 377916 586656 381360 586684
rect 377916 586644 377922 586656
rect 381354 586644 381360 586656
rect 381412 586644 381418 586696
rect 377214 585216 377220 585268
rect 377272 585256 377278 585268
rect 379974 585256 379980 585268
rect 377272 585228 379980 585256
rect 377272 585216 377278 585228
rect 379974 585216 379980 585228
rect 380032 585216 380038 585268
rect 137554 585148 137560 585200
rect 137612 585188 137618 585200
rect 144270 585188 144276 585200
rect 137612 585160 144276 585188
rect 137612 585148 137618 585160
rect 144270 585148 144276 585160
rect 144328 585148 144334 585200
rect 377030 585148 377036 585200
rect 377088 585188 377094 585200
rect 379698 585188 379704 585200
rect 377088 585160 379704 585188
rect 377088 585148 377094 585160
rect 379698 585148 379704 585160
rect 379756 585148 379762 585200
rect 416038 584740 416044 584792
rect 416096 584780 416102 584792
rect 423582 584780 423588 584792
rect 416096 584752 423588 584780
rect 416096 584740 416102 584752
rect 423582 584740 423588 584752
rect 423640 584740 423646 584792
rect 377766 583720 377772 583772
rect 377824 583760 377830 583772
rect 381262 583760 381268 583772
rect 377824 583732 381268 583760
rect 377824 583720 377830 583732
rect 381262 583720 381268 583732
rect 381320 583720 381326 583772
rect 378042 582768 378048 582820
rect 378100 582808 378106 582820
rect 382366 582808 382372 582820
rect 378100 582780 382372 582808
rect 378100 582768 378106 582780
rect 382366 582768 382372 582780
rect 382424 582768 382430 582820
rect 378042 582428 378048 582480
rect 378100 582468 378106 582480
rect 383930 582468 383936 582480
rect 378100 582440 383936 582468
rect 378100 582428 378106 582440
rect 383930 582428 383936 582440
rect 383988 582428 383994 582480
rect 378042 581000 378048 581052
rect 378100 581040 378106 581052
rect 383746 581040 383752 581052
rect 378100 581012 383752 581040
rect 378100 581000 378106 581012
rect 383746 581000 383752 581012
rect 383804 581000 383810 581052
rect 423582 580252 423588 580304
rect 423640 580292 423646 580304
rect 432598 580292 432604 580304
rect 423640 580264 432604 580292
rect 423640 580252 423646 580264
rect 432598 580252 432604 580264
rect 432656 580252 432662 580304
rect 3418 579640 3424 579692
rect 3476 579680 3482 579692
rect 47578 579680 47584 579692
rect 3476 579652 47584 579680
rect 3476 579640 3482 579652
rect 47578 579640 47584 579652
rect 47636 579640 47642 579692
rect 378042 579640 378048 579692
rect 378100 579680 378106 579692
rect 382458 579680 382464 579692
rect 378100 579652 382464 579680
rect 378100 579640 378106 579652
rect 382458 579640 382464 579652
rect 382516 579640 382522 579692
rect 378042 578280 378048 578332
rect 378100 578320 378106 578332
rect 382550 578320 382556 578332
rect 378100 578292 382556 578320
rect 378100 578280 378106 578292
rect 382550 578280 382556 578292
rect 382608 578280 382614 578332
rect 377030 578212 377036 578264
rect 377088 578252 377094 578264
rect 379882 578252 379888 578264
rect 377088 578224 379888 578252
rect 377088 578212 377094 578224
rect 379882 578212 379888 578224
rect 379940 578212 379946 578264
rect 134702 575492 134708 575544
rect 134760 575532 134766 575544
rect 137554 575532 137560 575544
rect 134760 575504 137560 575532
rect 134760 575492 134766 575504
rect 137554 575492 137560 575504
rect 137612 575492 137618 575544
rect 454678 574744 454684 574796
rect 454736 574784 454742 574796
rect 475378 574784 475384 574796
rect 454736 574756 475384 574784
rect 454736 574744 454742 574756
rect 475378 574744 475384 574756
rect 475436 574744 475442 574796
rect 378042 574064 378048 574116
rect 378100 574104 378106 574116
rect 386782 574104 386788 574116
rect 378100 574076 386788 574104
rect 378100 574064 378106 574076
rect 386782 574064 386788 574076
rect 386840 574064 386846 574116
rect 377582 572704 377588 572756
rect 377640 572744 377646 572756
rect 380894 572744 380900 572756
rect 377640 572716 380900 572744
rect 377640 572704 377646 572716
rect 380894 572704 380900 572716
rect 380952 572704 380958 572756
rect 166626 569780 166632 569832
rect 166684 569820 166690 569832
rect 172238 569820 172244 569832
rect 166684 569792 172244 569820
rect 166684 569780 166690 569792
rect 172238 569780 172244 569792
rect 172296 569780 172302 569832
rect 377950 568556 377956 568608
rect 378008 568596 378014 568608
rect 381630 568596 381636 568608
rect 378008 568568 381636 568596
rect 378008 568556 378014 568568
rect 381630 568556 381636 568568
rect 381688 568556 381694 568608
rect 285030 567196 285036 567248
rect 285088 567236 285094 567248
rect 296714 567236 296720 567248
rect 285088 567208 296720 567236
rect 285088 567196 285094 567208
rect 296714 567196 296720 567208
rect 296772 567196 296778 567248
rect 56962 563184 56968 563236
rect 57020 563224 57026 563236
rect 57514 563224 57520 563236
rect 57020 563196 57520 563224
rect 57020 563184 57026 563196
rect 57514 563184 57520 563196
rect 57572 563184 57578 563236
rect 291930 560872 291936 560924
rect 291988 560912 291994 560924
rect 298002 560912 298008 560924
rect 291988 560884 298008 560912
rect 291988 560872 291994 560884
rect 298002 560872 298008 560884
rect 298060 560872 298066 560924
rect 98730 560600 98736 560652
rect 98788 560640 98794 560652
rect 160830 560640 160836 560652
rect 98788 560612 160836 560640
rect 98788 560600 98794 560612
rect 160830 560600 160836 560612
rect 160888 560600 160894 560652
rect 178586 560600 178592 560652
rect 178644 560640 178650 560652
rect 288158 560640 288164 560652
rect 178644 560612 288164 560640
rect 178644 560600 178650 560612
rect 288158 560600 288164 560612
rect 288216 560600 288222 560652
rect 179414 560532 179420 560584
rect 179472 560572 179478 560584
rect 285306 560572 285312 560584
rect 179472 560544 285312 560572
rect 179472 560532 179478 560544
rect 285306 560532 285312 560544
rect 285364 560532 285370 560584
rect 179230 560328 179236 560380
rect 179288 560368 179294 560380
rect 179506 560368 179512 560380
rect 179288 560340 179512 560368
rect 179288 560328 179294 560340
rect 179506 560328 179512 560340
rect 179564 560328 179570 560380
rect 57330 560260 57336 560312
rect 57388 560300 57394 560312
rect 58066 560300 58072 560312
rect 57388 560272 58072 560300
rect 57388 560260 57394 560272
rect 58066 560260 58072 560272
rect 58124 560260 58130 560312
rect 299750 560260 299756 560312
rect 299808 560300 299814 560312
rect 309778 560300 309784 560312
rect 299808 560272 309784 560300
rect 299808 560260 299814 560272
rect 309778 560260 309784 560272
rect 309836 560260 309842 560312
rect 57606 560192 57612 560244
rect 57664 560232 57670 560244
rect 376110 560232 376116 560244
rect 57664 560204 376116 560232
rect 57664 560192 57670 560204
rect 376110 560192 376116 560204
rect 376168 560192 376174 560244
rect 57330 560124 57336 560176
rect 57388 560164 57394 560176
rect 297818 560164 297824 560176
rect 57388 560136 297824 560164
rect 57388 560124 57394 560136
rect 297818 560124 297824 560136
rect 297876 560124 297882 560176
rect 57514 560056 57520 560108
rect 57572 560096 57578 560108
rect 297634 560096 297640 560108
rect 57572 560068 297640 560096
rect 57572 560056 57578 560068
rect 297634 560056 297640 560068
rect 297692 560056 297698 560108
rect 169386 559988 169392 560040
rect 169444 560028 169450 560040
rect 173066 560028 173072 560040
rect 169444 560000 173072 560028
rect 169444 559988 169450 560000
rect 173066 559988 173072 560000
rect 173124 559988 173130 560040
rect 166810 559920 166816 559972
rect 166868 559960 166874 559972
rect 173802 559960 173808 559972
rect 166868 559932 173808 559960
rect 166868 559920 166874 559932
rect 173802 559920 173808 559932
rect 173860 559920 173866 559972
rect 372062 559852 372068 559904
rect 372120 559892 372126 559904
rect 379974 559892 379980 559904
rect 372120 559864 379980 559892
rect 372120 559852 372126 559864
rect 379974 559852 379980 559864
rect 380032 559852 380038 559904
rect 371878 559784 371884 559836
rect 371936 559824 371942 559836
rect 379790 559824 379796 559836
rect 371936 559796 379796 559824
rect 371936 559784 371942 559796
rect 379790 559784 379796 559796
rect 379848 559784 379854 559836
rect 371970 559716 371976 559768
rect 372028 559756 372034 559768
rect 381262 559756 381268 559768
rect 372028 559728 381268 559756
rect 372028 559716 372034 559728
rect 381262 559716 381268 559728
rect 381320 559716 381326 559768
rect 372154 559648 372160 559700
rect 372212 559688 372218 559700
rect 381446 559688 381452 559700
rect 372212 559660 381452 559688
rect 372212 559648 372218 559660
rect 381446 559648 381452 559660
rect 381504 559648 381510 559700
rect 90910 559580 90916 559632
rect 90968 559620 90974 559632
rect 139578 559620 139584 559632
rect 90968 559592 139584 559620
rect 90968 559580 90974 559592
rect 139578 559580 139584 559592
rect 139636 559580 139642 559632
rect 268378 559580 268384 559632
rect 268436 559620 268442 559632
rect 514754 559620 514760 559632
rect 268436 559592 514760 559620
rect 268436 559580 268442 559592
rect 514754 559580 514760 559592
rect 514812 559580 514818 559632
rect 76006 559512 76012 559564
rect 76064 559552 76070 559564
rect 135162 559552 135168 559564
rect 76064 559524 135168 559552
rect 76064 559512 76070 559524
rect 135162 559512 135168 559524
rect 135220 559512 135226 559564
rect 177206 559512 177212 559564
rect 177264 559552 177270 559564
rect 487154 559552 487160 559564
rect 177264 559524 487160 559552
rect 177264 559512 177270 559524
rect 487154 559512 487160 559524
rect 487212 559512 487218 559564
rect 63770 558900 63776 558952
rect 63828 558940 63834 558952
rect 68278 558940 68284 558952
rect 63828 558912 68284 558940
rect 63828 558900 63834 558912
rect 68278 558900 68284 558912
rect 68336 558900 68342 558952
rect 97810 558900 97816 558952
rect 97868 558940 97874 558952
rect 254578 558940 254584 558952
rect 97868 558912 254584 558940
rect 97868 558900 97874 558912
rect 254578 558900 254584 558912
rect 254636 558900 254642 558952
rect 57606 558832 57612 558884
rect 57664 558872 57670 558884
rect 381354 558872 381360 558884
rect 57664 558844 381360 558872
rect 57664 558832 57670 558844
rect 381354 558832 381360 558844
rect 381412 558832 381418 558884
rect 56502 558764 56508 558816
rect 56560 558804 56566 558816
rect 361206 558804 361212 558816
rect 56560 558776 361212 558804
rect 56560 558764 56566 558776
rect 361206 558764 361212 558776
rect 361264 558764 361270 558816
rect 47946 558696 47952 558748
rect 48004 558736 48010 558748
rect 98730 558736 98736 558748
rect 48004 558708 98736 558736
rect 48004 558696 48010 558708
rect 98730 558696 98736 558708
rect 98788 558696 98794 558748
rect 109126 558696 109132 558748
rect 109184 558736 109190 558748
rect 289354 558736 289360 558748
rect 109184 558708 289360 558736
rect 109184 558696 109190 558708
rect 289354 558696 289360 558708
rect 289412 558696 289418 558748
rect 120074 558628 120080 558680
rect 120132 558668 120138 558680
rect 163866 558668 163872 558680
rect 120132 558640 163872 558668
rect 120132 558628 120138 558640
rect 163866 558628 163872 558640
rect 163924 558628 163930 558680
rect 279786 558424 279792 558476
rect 279844 558464 279850 558476
rect 506658 558464 506664 558476
rect 279844 558436 506664 558464
rect 279844 558424 279850 558436
rect 506658 558424 506664 558436
rect 506716 558424 506722 558476
rect 60458 558356 60464 558408
rect 60516 558396 60522 558408
rect 297542 558396 297548 558408
rect 60516 558368 297548 558396
rect 60516 558356 60522 558368
rect 297542 558356 297548 558368
rect 297600 558356 297606 558408
rect 60550 558288 60556 558340
rect 60608 558328 60614 558340
rect 298738 558328 298744 558340
rect 60608 558300 298744 558328
rect 60608 558288 60614 558300
rect 298738 558288 298744 558300
rect 298796 558288 298802 558340
rect 271230 558220 271236 558272
rect 271288 558260 271294 558272
rect 511994 558260 512000 558272
rect 271288 558232 512000 558260
rect 271288 558220 271294 558232
rect 511994 558220 512000 558232
rect 512052 558220 512058 558272
rect 59630 558152 59636 558204
rect 59688 558192 59694 558204
rect 360194 558192 360200 558204
rect 59688 558164 360200 558192
rect 59688 558152 59694 558164
rect 360194 558152 360200 558164
rect 360252 558152 360258 558204
rect 372614 558152 372620 558204
rect 372672 558192 372678 558204
rect 377122 558192 377128 558204
rect 372672 558164 377128 558192
rect 372672 558152 372678 558164
rect 377122 558152 377128 558164
rect 377180 558152 377186 558204
rect 117958 557676 117964 557728
rect 118016 557716 118022 557728
rect 216122 557716 216128 557728
rect 118016 557688 216128 557716
rect 118016 557676 118022 557688
rect 216122 557676 216128 557688
rect 216180 557676 216186 557728
rect 120166 557608 120172 557660
rect 120224 557648 120230 557660
rect 253290 557648 253296 557660
rect 120224 557620 253296 557648
rect 120224 557608 120230 557620
rect 253290 557608 253296 557620
rect 253348 557608 253354 557660
rect 280154 557608 280160 557660
rect 280212 557648 280218 557660
rect 492766 557648 492772 557660
rect 280212 557620 492772 557648
rect 280212 557608 280218 557620
rect 492766 557608 492772 557620
rect 492824 557608 492830 557660
rect 117774 557540 117780 557592
rect 117832 557580 117838 557592
rect 259822 557580 259828 557592
rect 117832 557552 259828 557580
rect 117832 557540 117838 557552
rect 259822 557540 259828 557552
rect 259880 557540 259886 557592
rect 284202 557540 284208 557592
rect 284260 557580 284266 557592
rect 509418 557580 509424 557592
rect 284260 557552 509424 557580
rect 284260 557540 284266 557552
rect 509418 557540 509424 557552
rect 509476 557540 509482 557592
rect 56502 557472 56508 557524
rect 56560 557512 56566 557524
rect 379698 557512 379704 557524
rect 56560 557484 379704 557512
rect 56560 557472 56566 557484
rect 379698 557472 379704 557484
rect 379756 557472 379762 557524
rect 55858 557404 55864 557456
rect 55916 557444 55922 557456
rect 377030 557444 377036 557456
rect 55916 557416 377036 557444
rect 55916 557404 55922 557416
rect 377030 557404 377036 557416
rect 377088 557404 377094 557456
rect 60090 557336 60096 557388
rect 60148 557376 60154 557388
rect 376018 557376 376024 557388
rect 60148 557348 376024 557376
rect 60148 557336 60154 557348
rect 376018 557336 376024 557348
rect 376076 557336 376082 557388
rect 95142 557268 95148 557320
rect 95200 557308 95206 557320
rect 297910 557308 297916 557320
rect 95200 557280 297916 557308
rect 95200 557268 95206 557280
rect 297910 557268 297916 557280
rect 297968 557268 297974 557320
rect 265618 556860 265624 556912
rect 265676 556900 265682 556912
rect 512086 556900 512092 556912
rect 265676 556872 512092 556900
rect 265676 556860 265682 556872
rect 512086 556860 512092 556872
rect 512144 556860 512150 556912
rect 50614 556792 50620 556844
rect 50672 556832 50678 556844
rect 92382 556832 92388 556844
rect 50672 556804 92388 556832
rect 50672 556792 50678 556804
rect 92382 556792 92388 556804
rect 92440 556832 92446 556844
rect 163774 556832 163780 556844
rect 92440 556804 163780 556832
rect 92440 556792 92446 556804
rect 163774 556792 163780 556804
rect 163832 556792 163838 556844
rect 175090 556792 175096 556844
rect 175148 556832 175154 556844
rect 424042 556832 424048 556844
rect 175148 556804 424048 556832
rect 175148 556792 175154 556804
rect 424042 556792 424048 556804
rect 424100 556792 424106 556844
rect 86954 556180 86960 556232
rect 87012 556220 87018 556232
rect 90910 556220 90916 556232
rect 87012 556192 90916 556220
rect 87012 556180 87018 556192
rect 90910 556180 90916 556192
rect 90968 556180 90974 556232
rect 178034 556180 178040 556232
rect 178092 556220 178098 556232
rect 422478 556220 422484 556232
rect 178092 556192 422484 556220
rect 178092 556180 178098 556192
rect 422478 556180 422484 556192
rect 422536 556180 422542 556232
rect 100754 556112 100760 556164
rect 100812 556152 100818 556164
rect 378686 556152 378692 556164
rect 100812 556124 378692 556152
rect 100812 556112 100818 556124
rect 378686 556112 378692 556124
rect 378744 556112 378750 556164
rect 121454 556044 121460 556096
rect 121512 556084 121518 556096
rect 339954 556084 339960 556096
rect 121512 556056 339960 556084
rect 121512 556044 121518 556056
rect 339954 556044 339960 556056
rect 340012 556044 340018 556096
rect 332594 555568 332600 555620
rect 332652 555608 332658 555620
rect 372614 555608 372620 555620
rect 332652 555580 372620 555608
rect 332652 555568 332658 555580
rect 372614 555568 372620 555580
rect 372672 555568 372678 555620
rect 137278 555500 137284 555552
rect 137336 555540 137342 555552
rect 360838 555540 360844 555552
rect 137336 555512 360844 555540
rect 137336 555500 137342 555512
rect 360838 555500 360844 555512
rect 360896 555500 360902 555552
rect 57146 555432 57152 555484
rect 57204 555472 57210 555484
rect 375926 555472 375932 555484
rect 57204 555444 375932 555472
rect 57204 555432 57210 555444
rect 375926 555432 375932 555444
rect 375984 555432 375990 555484
rect 57698 555160 57704 555212
rect 57756 555160 57762 555212
rect 57716 555008 57744 555160
rect 57698 554956 57704 555008
rect 57756 554956 57762 555008
rect 58618 554752 58624 554804
rect 58676 554752 58682 554804
rect 124122 554752 124128 554804
rect 124180 554792 124186 554804
rect 262950 554792 262956 554804
rect 124180 554764 262956 554792
rect 124180 554752 124186 554764
rect 262950 554752 262956 554764
rect 263008 554752 263014 554804
rect 275922 554752 275928 554804
rect 275980 554792 275986 554804
rect 492858 554792 492864 554804
rect 275980 554764 492864 554792
rect 275980 554752 275986 554764
rect 492858 554752 492864 554764
rect 492916 554752 492922 554804
rect 58636 554600 58664 554752
rect 73154 554684 73160 554736
rect 73212 554724 73218 554736
rect 350074 554724 350080 554736
rect 73212 554696 350080 554724
rect 73212 554684 73218 554696
rect 350074 554684 350080 554696
rect 350132 554684 350138 554736
rect 88978 554616 88984 554668
rect 89036 554656 89042 554668
rect 310606 554656 310612 554668
rect 89036 554628 310612 554656
rect 89036 554616 89042 554628
rect 310606 554616 310612 554628
rect 310664 554616 310670 554668
rect 58618 554548 58624 554600
rect 58676 554548 58682 554600
rect 107562 554548 107568 554600
rect 107620 554588 107626 554600
rect 297450 554588 297456 554600
rect 107620 554560 297456 554588
rect 107620 554548 107626 554560
rect 297450 554548 297456 554560
rect 297508 554548 297514 554600
rect 136082 554004 136088 554056
rect 136140 554044 136146 554056
rect 320818 554044 320824 554056
rect 136140 554016 320824 554044
rect 136140 554004 136146 554016
rect 320818 554004 320824 554016
rect 320876 554004 320882 554056
rect 115842 553460 115848 553512
rect 115900 553500 115906 553512
rect 247310 553500 247316 553512
rect 115900 553472 247316 553500
rect 115900 553460 115906 553472
rect 247310 553460 247316 553472
rect 247368 553460 247374 553512
rect 299290 553460 299296 553512
rect 299348 553500 299354 553512
rect 489086 553500 489092 553512
rect 299348 553472 489092 553500
rect 299348 553460 299354 553472
rect 489086 553460 489092 553472
rect 489144 553460 489150 553512
rect 108298 553392 108304 553444
rect 108356 553432 108362 553444
rect 258258 553432 258264 553444
rect 108356 553404 258264 553432
rect 108356 553392 108362 553404
rect 258258 553392 258264 553404
rect 258316 553392 258322 553444
rect 293954 553392 293960 553444
rect 294012 553432 294018 553444
rect 493042 553432 493048 553444
rect 294012 553404 493048 553432
rect 294012 553392 294018 553404
rect 493042 553392 493048 553404
rect 493100 553392 493106 553444
rect 81434 553324 81440 553376
rect 81492 553364 81498 553376
rect 347038 553364 347044 553376
rect 81492 553336 347044 553364
rect 81492 553324 81498 553336
rect 347038 553324 347044 553336
rect 347096 553324 347102 553376
rect 57790 553256 57796 553308
rect 57848 553296 57854 553308
rect 286410 553296 286416 553308
rect 57848 553268 286416 553296
rect 57848 553256 57854 553268
rect 286410 553256 286416 553268
rect 286468 553256 286474 553308
rect 299290 553256 299296 553308
rect 299348 553296 299354 553308
rect 303522 553296 303528 553308
rect 299348 553268 303528 553296
rect 299348 553256 299354 553268
rect 303522 553256 303528 553268
rect 303580 553256 303586 553308
rect 98638 553188 98644 553240
rect 98696 553228 98702 553240
rect 305546 553228 305552 553240
rect 98696 553200 305552 553228
rect 98696 553188 98702 553200
rect 305546 553188 305552 553200
rect 305604 553188 305610 553240
rect 179414 553120 179420 553172
rect 179472 553160 179478 553172
rect 297726 553160 297732 553172
rect 179472 553132 297732 553160
rect 179472 553120 179478 553132
rect 297726 553120 297732 553132
rect 297784 553120 297790 553172
rect 47578 552644 47584 552696
rect 47636 552684 47642 552696
rect 60550 552684 60556 552696
rect 47636 552656 60556 552684
rect 47636 552644 47642 552656
rect 60550 552644 60556 552656
rect 60608 552684 60614 552696
rect 151078 552684 151084 552696
rect 60608 552656 151084 552684
rect 60608 552644 60614 552656
rect 151078 552644 151084 552656
rect 151136 552644 151142 552696
rect 304258 552644 304264 552696
rect 304316 552684 304322 552696
rect 332594 552684 332600 552696
rect 304316 552656 332600 552684
rect 304316 552644 304322 552656
rect 332594 552644 332600 552656
rect 332652 552644 332658 552696
rect 173802 552372 173808 552424
rect 173860 552412 173866 552424
rect 509326 552412 509332 552424
rect 173860 552384 509332 552412
rect 173860 552372 173866 552384
rect 509326 552372 509332 552384
rect 509384 552372 509390 552424
rect 295334 552304 295340 552356
rect 295392 552344 295398 552356
rect 358354 552344 358360 552356
rect 295392 552316 358360 552344
rect 295392 552304 295398 552316
rect 358354 552304 358360 552316
rect 358412 552304 358418 552356
rect 291746 552236 291752 552288
rect 291804 552276 291810 552288
rect 439682 552276 439688 552288
rect 291804 552248 439688 552276
rect 291804 552236 291810 552248
rect 439682 552236 439688 552248
rect 439740 552236 439746 552288
rect 278682 552168 278688 552220
rect 278740 552208 278746 552220
rect 491294 552208 491300 552220
rect 278740 552180 491300 552208
rect 278740 552168 278746 552180
rect 491294 552168 491300 552180
rect 491352 552168 491358 552220
rect 175826 552100 175832 552152
rect 175884 552140 175890 552152
rect 502518 552140 502524 552152
rect 175884 552112 502524 552140
rect 175884 552100 175890 552112
rect 502518 552100 502524 552112
rect 502576 552100 502582 552152
rect 58710 552032 58716 552084
rect 58768 552072 58774 552084
rect 169754 552072 169760 552084
rect 58768 552044 169760 552072
rect 58768 552032 58774 552044
rect 169754 552032 169760 552044
rect 169812 552032 169818 552084
rect 52454 551964 52460 552016
rect 52512 552004 52518 552016
rect 356146 552004 356152 552016
rect 52512 551976 356152 552004
rect 52512 551964 52518 551976
rect 356146 551964 356152 551976
rect 356204 551964 356210 552016
rect 59262 551896 59268 551948
rect 59320 551936 59326 551948
rect 348050 551936 348056 551948
rect 59320 551908 348056 551936
rect 59320 551896 59326 551908
rect 348050 551896 348056 551908
rect 348108 551896 348114 551948
rect 99374 551828 99380 551880
rect 99432 551868 99438 551880
rect 379882 551868 379888 551880
rect 99432 551840 379888 551868
rect 99432 551828 99438 551840
rect 379882 551828 379888 551840
rect 379940 551828 379946 551880
rect 81434 551760 81440 551812
rect 81492 551800 81498 551812
rect 328822 551800 328828 551812
rect 81492 551772 328828 551800
rect 81492 551760 81498 551772
rect 328822 551760 328828 551772
rect 328880 551760 328886 551812
rect 124858 551352 124864 551404
rect 124916 551392 124922 551404
rect 134702 551392 134708 551404
rect 124916 551364 134708 551392
rect 124916 551352 124922 551364
rect 134702 551352 134708 551364
rect 134760 551352 134766 551404
rect 60090 551284 60096 551336
rect 60148 551324 60154 551336
rect 359182 551324 359188 551336
rect 60148 551296 359188 551324
rect 60148 551284 60154 551296
rect 359182 551284 359188 551296
rect 359240 551284 359246 551336
rect 269114 550740 269120 550792
rect 269172 550780 269178 550792
rect 469398 550780 469404 550792
rect 269172 550752 469404 550780
rect 269172 550740 269178 550752
rect 469398 550740 469404 550752
rect 469456 550740 469462 550792
rect 241422 550672 241428 550724
rect 241480 550712 241486 550724
rect 492950 550712 492956 550724
rect 241480 550684 492956 550712
rect 241480 550672 241486 550684
rect 492950 550672 492956 550684
rect 493008 550672 493014 550724
rect 178034 550604 178040 550656
rect 178092 550644 178098 550656
rect 497458 550644 497464 550656
rect 178092 550616 497464 550644
rect 178092 550604 178098 550616
rect 497458 550604 497464 550616
rect 497516 550604 497522 550656
rect 85482 550536 85488 550588
rect 85540 550576 85546 550588
rect 365254 550576 365260 550588
rect 85540 550548 365260 550576
rect 85540 550536 85546 550548
rect 365254 550536 365260 550548
rect 365312 550536 365318 550588
rect 100754 550468 100760 550520
rect 100812 550508 100818 550520
rect 353110 550508 353116 550520
rect 100812 550480 353116 550508
rect 100812 550468 100818 550480
rect 353110 550468 353116 550480
rect 353168 550468 353174 550520
rect 179414 550400 179420 550452
rect 179472 550440 179478 550452
rect 380894 550440 380900 550452
rect 179472 550412 380900 550440
rect 179472 550400 179478 550412
rect 380894 550400 380900 550412
rect 380952 550400 380958 550452
rect 169754 550332 169760 550384
rect 169812 550372 169818 550384
rect 326798 550372 326804 550384
rect 169812 550344 326804 550372
rect 169812 550332 169818 550344
rect 326798 550332 326804 550344
rect 326856 550332 326862 550384
rect 233142 550264 233148 550316
rect 233200 550304 233206 550316
rect 283834 550304 283840 550316
rect 233200 550276 283840 550304
rect 233200 550264 233206 550276
rect 283834 550264 283840 550276
rect 283892 550264 283898 550316
rect 273898 550060 273904 550112
rect 273956 550100 273962 550112
rect 352098 550100 352104 550112
rect 273956 550072 352104 550100
rect 273956 550060 273962 550072
rect 352098 550060 352104 550072
rect 352156 550060 352162 550112
rect 283742 549992 283748 550044
rect 283800 550032 283806 550044
rect 364610 550032 364616 550044
rect 283800 550004 364616 550032
rect 283800 549992 283806 550004
rect 364610 549992 364616 550004
rect 364668 549992 364674 550044
rect 134610 549924 134616 549976
rect 134668 549964 134674 549976
rect 328638 549964 328644 549976
rect 134668 549936 328644 549964
rect 134668 549924 134674 549936
rect 328638 549924 328644 549936
rect 328696 549924 328702 549976
rect 177298 549856 177304 549908
rect 177356 549896 177362 549908
rect 491662 549896 491668 549908
rect 177356 549868 491668 549896
rect 177356 549856 177362 549868
rect 491662 549856 491668 549868
rect 491720 549856 491726 549908
rect 86862 549488 86868 549500
rect 84166 549460 86868 549488
rect 71038 549244 71044 549296
rect 71096 549284 71102 549296
rect 75822 549284 75828 549296
rect 71096 549256 75828 549284
rect 71096 549244 71102 549256
rect 75822 549244 75828 549256
rect 75880 549244 75886 549296
rect 81802 549244 81808 549296
rect 81860 549284 81866 549296
rect 84166 549284 84194 549460
rect 86862 549448 86868 549460
rect 86920 549448 86926 549500
rect 81860 549256 84194 549284
rect 81860 549244 81866 549256
rect 224954 549244 224960 549296
rect 225012 549284 225018 549296
rect 260788 549284 260794 549296
rect 225012 549256 260794 549284
rect 225012 549244 225018 549256
rect 260788 549244 260794 549256
rect 260846 549244 260852 549296
rect 260926 549244 260932 549296
rect 260984 549284 260990 549296
rect 487614 549284 487620 549296
rect 260984 549256 487620 549284
rect 260984 549244 260990 549256
rect 487614 549244 487620 549256
rect 487672 549244 487678 549296
rect 86862 549176 86868 549228
rect 86920 549216 86926 549228
rect 342990 549216 342996 549228
rect 86920 549188 342996 549216
rect 86920 549176 86926 549188
rect 342990 549176 342996 549188
rect 343048 549176 343054 549228
rect 75822 549108 75828 549160
rect 75880 549148 75886 549160
rect 260834 549148 260840 549160
rect 75880 549120 260840 549148
rect 75880 549108 75886 549120
rect 260834 549108 260840 549120
rect 260892 549108 260898 549160
rect 265636 549120 270494 549148
rect 126882 549040 126888 549092
rect 126940 549080 126946 549092
rect 265636 549080 265664 549120
rect 126940 549052 265664 549080
rect 270466 549080 270494 549120
rect 280062 549108 280068 549160
rect 280120 549148 280126 549160
rect 313642 549148 313648 549160
rect 280120 549120 313648 549148
rect 280120 549108 280126 549120
rect 313642 549108 313648 549120
rect 313700 549108 313706 549160
rect 322750 549080 322756 549092
rect 270466 549052 322756 549080
rect 126940 549040 126946 549052
rect 322750 549040 322756 549052
rect 322808 549040 322814 549092
rect 59262 548972 59268 549024
rect 59320 549012 59326 549024
rect 159358 549012 159364 549024
rect 59320 548984 159364 549012
rect 59320 548972 59326 548984
rect 159358 548972 159364 548984
rect 159416 548972 159422 549024
rect 260926 548972 260932 549024
rect 260984 549012 260990 549024
rect 279694 549012 279700 549024
rect 260984 548984 279700 549012
rect 260984 548972 260990 548984
rect 279694 548972 279700 548984
rect 279752 548972 279758 549024
rect 162302 548632 162308 548684
rect 162360 548672 162366 548684
rect 363046 548672 363052 548684
rect 162360 548644 363052 548672
rect 162360 548632 162366 548644
rect 363046 548632 363052 548644
rect 363104 548632 363110 548684
rect 432598 548632 432604 548684
rect 432656 548672 432662 548684
rect 443638 548672 443644 548684
rect 432656 548644 443644 548672
rect 432656 548632 432662 548644
rect 443638 548632 443644 548644
rect 443696 548632 443702 548684
rect 202782 548564 202788 548616
rect 202840 548604 202846 548616
rect 502334 548604 502340 548616
rect 202840 548576 502340 548604
rect 202840 548564 202846 548576
rect 502334 548564 502340 548576
rect 502392 548564 502398 548616
rect 177114 548496 177120 548548
rect 177172 548536 177178 548548
rect 493134 548536 493140 548548
rect 177172 548508 493140 548536
rect 177172 548496 177178 548508
rect 493134 548496 493140 548508
rect 493192 548496 493198 548548
rect 58710 548292 58716 548344
rect 58768 548332 58774 548344
rect 59262 548332 59268 548344
rect 58768 548304 59268 548332
rect 58768 548292 58774 548304
rect 59262 548292 59268 548304
rect 59320 548292 59326 548344
rect 278682 547884 278688 547936
rect 278740 547924 278746 547936
rect 514846 547924 514852 547936
rect 278740 547896 514852 547924
rect 278740 547884 278746 547896
rect 514846 547884 514852 547896
rect 514904 547884 514910 547936
rect 78582 547816 78588 547868
rect 78640 547856 78646 547868
rect 375650 547856 375656 547868
rect 78640 547828 375656 547856
rect 78640 547816 78646 547828
rect 375650 547816 375656 547828
rect 375708 547816 375714 547868
rect 89714 547748 89720 547800
rect 89772 547788 89778 547800
rect 346026 547788 346032 547800
rect 89772 547760 346032 547788
rect 89772 547748 89778 547760
rect 346026 547748 346032 547760
rect 346084 547748 346090 547800
rect 126882 547680 126888 547732
rect 126940 547720 126946 547732
rect 320726 547720 320732 547732
rect 126940 547692 320732 547720
rect 126940 547680 126946 547692
rect 320726 547680 320732 547692
rect 320784 547680 320790 547732
rect 216674 547612 216680 547664
rect 216732 547652 216738 547664
rect 306558 547652 306564 547664
rect 216732 547624 306564 547652
rect 216732 547612 216738 547624
rect 306558 547612 306564 547624
rect 306616 547612 306622 547664
rect 135990 547272 135996 547324
rect 136048 547312 136054 547324
rect 356790 547312 356796 547324
rect 136048 547284 356796 547312
rect 136048 547272 136054 547284
rect 356790 547272 356796 547284
rect 356848 547272 356854 547324
rect 226058 547204 226064 547256
rect 226116 547244 226122 547256
rect 486142 547244 486148 547256
rect 226116 547216 486148 547244
rect 226116 547204 226122 547216
rect 486142 547204 486148 547216
rect 486200 547204 486206 547256
rect 188614 547136 188620 547188
rect 188672 547176 188678 547188
rect 495434 547176 495440 547188
rect 188672 547148 495440 547176
rect 188672 547136 188678 547148
rect 495434 547136 495440 547148
rect 495492 547136 495498 547188
rect 230382 546524 230388 546576
rect 230440 546564 230446 546576
rect 305178 546564 305184 546576
rect 230440 546536 305184 546564
rect 230440 546524 230446 546536
rect 305178 546524 305184 546536
rect 305236 546524 305242 546576
rect 173802 546456 173808 546508
rect 173860 546496 173866 546508
rect 456886 546496 456892 546508
rect 173860 546468 456892 546496
rect 173860 546456 173866 546468
rect 456886 546456 456892 546468
rect 456944 546456 456950 546508
rect 60182 546388 60188 546440
rect 60240 546428 60246 546440
rect 372338 546428 372344 546440
rect 60240 546400 372344 546428
rect 60240 546388 60246 546400
rect 372338 546388 372344 546400
rect 372396 546388 372402 546440
rect 189626 546320 189632 546372
rect 189684 546360 189690 546372
rect 485774 546360 485780 546372
rect 189684 546332 485780 546360
rect 189684 546320 189690 546332
rect 485774 546320 485780 546332
rect 485832 546320 485838 546372
rect 79318 546252 79324 546304
rect 79376 546292 79382 546304
rect 362218 546292 362224 546304
rect 79376 546264 362224 546292
rect 79376 546252 79382 546264
rect 362218 546252 362224 546264
rect 362276 546252 362282 546304
rect 121454 546184 121460 546236
rect 121512 546224 121518 546236
rect 323762 546224 323768 546236
rect 121512 546196 323768 546224
rect 121512 546184 121518 546196
rect 323762 546184 323768 546196
rect 323820 546184 323826 546236
rect 89714 546116 89720 546168
rect 89772 546156 89778 546168
rect 284938 546156 284944 546168
rect 89772 546128 284944 546156
rect 89772 546116 89778 546128
rect 284938 546116 284944 546128
rect 284996 546116 285002 546168
rect 223482 546048 223488 546100
rect 223540 546088 223546 546100
rect 382642 546088 382648 546100
rect 223540 546060 382648 546088
rect 223540 546048 223546 546060
rect 382642 546048 382648 546060
rect 382700 546048 382706 546100
rect 207842 545708 207848 545760
rect 207900 545748 207906 545760
rect 503990 545748 503996 545760
rect 207900 545720 503996 545748
rect 207900 545708 207906 545720
rect 503990 545708 503996 545720
rect 504048 545708 504054 545760
rect 75822 545164 75828 545216
rect 75880 545204 75886 545216
rect 81802 545204 81808 545216
rect 75880 545176 81808 545204
rect 75880 545164 75886 545176
rect 81802 545164 81808 545176
rect 81860 545164 81866 545216
rect 92474 545028 92480 545080
rect 92532 545068 92538 545080
rect 381170 545068 381176 545080
rect 92532 545040 381176 545068
rect 92532 545028 92538 545040
rect 381170 545028 381176 545040
rect 381228 545028 381234 545080
rect 127618 544960 127624 545012
rect 127676 545000 127682 545012
rect 371326 545000 371332 545012
rect 127676 544972 371332 545000
rect 127676 544960 127682 544972
rect 371326 544960 371332 544972
rect 371384 544960 371390 545012
rect 153102 544892 153108 544944
rect 153160 544932 153166 544944
rect 308582 544932 308588 544944
rect 153160 544904 308588 544932
rect 153160 544892 153166 544904
rect 308582 544892 308588 544904
rect 308640 544892 308646 544944
rect 172422 544824 172428 544876
rect 172480 544864 172486 544876
rect 302510 544864 302516 544876
rect 172480 544836 302516 544864
rect 172480 544824 172486 544836
rect 302510 544824 302516 544836
rect 302568 544824 302574 544876
rect 215938 544416 215944 544468
rect 215996 544456 216002 544468
rect 494238 544456 494244 544468
rect 215996 544428 494244 544456
rect 215996 544416 216002 544428
rect 494238 544416 494244 544428
rect 494296 544416 494302 544468
rect 199746 544348 199752 544400
rect 199804 544388 199810 544400
rect 480530 544388 480536 544400
rect 199804 544360 480536 544388
rect 199804 544348 199810 544360
rect 480530 544348 480536 544360
rect 480588 544348 480594 544400
rect 293954 543804 293960 543856
rect 294012 543844 294018 543856
rect 348970 543844 348976 543856
rect 294012 543816 348976 543844
rect 294012 543804 294018 543816
rect 348970 543804 348976 543816
rect 349028 543804 349034 543856
rect 75822 543776 75828 543788
rect 74506 543748 75828 543776
rect 72418 543668 72424 543720
rect 72476 543708 72482 543720
rect 74506 543708 74534 543748
rect 75822 543736 75828 543748
rect 75880 543736 75886 543788
rect 175274 543736 175280 543788
rect 175332 543776 175338 543788
rect 436554 543776 436560 543788
rect 175332 543748 436560 543776
rect 175332 543736 175338 543748
rect 436554 543736 436560 543748
rect 436612 543736 436618 543788
rect 72476 543680 74534 543708
rect 72476 543668 72482 543680
rect 95142 543668 95148 543720
rect 95200 543708 95206 543720
rect 345014 543708 345020 543720
rect 95200 543680 345020 543708
rect 95200 543668 95206 543680
rect 345014 543668 345020 543680
rect 345072 543668 345078 543720
rect 125502 543600 125508 543652
rect 125560 543640 125566 543652
rect 318702 543640 318708 543652
rect 125560 543612 318708 543640
rect 125560 543600 125566 543612
rect 318702 543600 318708 543612
rect 318760 543600 318766 543652
rect 175274 543532 175280 543584
rect 175332 543572 175338 543584
rect 307570 543572 307576 543584
rect 175332 543544 307576 543572
rect 175332 543532 175338 543544
rect 307570 543532 307576 543544
rect 307628 543532 307634 543584
rect 283742 543124 283748 543176
rect 283800 543164 283806 543176
rect 357158 543164 357164 543176
rect 283800 543136 357164 543164
rect 283800 543124 283806 543136
rect 357158 543124 357164 543136
rect 357216 543124 357222 543176
rect 138750 543056 138756 543108
rect 138808 543096 138814 543108
rect 369210 543096 369216 543108
rect 138808 543068 369216 543096
rect 138808 543056 138814 543068
rect 369210 543056 369216 543068
rect 369268 543056 369274 543108
rect 177390 542988 177396 543040
rect 177448 543028 177454 543040
rect 494422 543028 494428 543040
rect 177448 543000 494428 543028
rect 177448 542988 177454 543000
rect 494422 542988 494428 543000
rect 494480 542988 494486 543040
rect 230382 542444 230388 542496
rect 230440 542484 230446 542496
rect 496998 542484 497004 542496
rect 230440 542456 497004 542484
rect 230440 542444 230446 542456
rect 496998 542444 497004 542456
rect 497056 542444 497062 542496
rect 172514 542376 172520 542428
rect 172572 542416 172578 542428
rect 466270 542416 466276 542428
rect 172572 542388 466276 542416
rect 172572 542376 172578 542388
rect 466270 542376 466276 542388
rect 466328 542376 466334 542428
rect 111794 542308 111800 542360
rect 111852 542348 111858 542360
rect 364242 542348 364248 542360
rect 111852 542320 364248 542348
rect 111852 542308 111858 542320
rect 364242 542308 364248 542320
rect 364300 542308 364306 542360
rect 224218 542240 224224 542292
rect 224276 542280 224282 542292
rect 386782 542280 386788 542292
rect 224276 542252 386788 542280
rect 224276 542240 224282 542252
rect 386782 542240 386788 542252
rect 386840 542240 386846 542292
rect 172514 542172 172520 542224
rect 172572 542212 172578 542224
rect 314654 542212 314660 542224
rect 172572 542184 314660 542212
rect 172572 542172 172578 542184
rect 314654 542172 314660 542184
rect 314712 542172 314718 542224
rect 135898 541832 135904 541884
rect 135956 541872 135962 541884
rect 355226 541872 355232 541884
rect 135956 541844 355232 541872
rect 135956 541832 135962 541844
rect 355226 541832 355232 541844
rect 355284 541832 355290 541884
rect 196710 541764 196716 541816
rect 196768 541804 196774 541816
rect 480622 541804 480628 541816
rect 196768 541776 480628 541804
rect 196768 541764 196774 541776
rect 480622 541764 480628 541776
rect 480680 541764 480686 541816
rect 187602 541696 187608 541748
rect 187660 541736 187666 541748
rect 496906 541736 496912 541748
rect 187660 541708 496912 541736
rect 187660 541696 187666 541708
rect 496906 541696 496912 541708
rect 496964 541696 496970 541748
rect 182542 541628 182548 541680
rect 182600 541668 182606 541680
rect 495526 541668 495532 541680
rect 182600 541640 495532 541668
rect 182600 541628 182606 541640
rect 495526 541628 495532 541640
rect 495584 541628 495590 541680
rect 233142 540948 233148 541000
rect 233200 540988 233206 541000
rect 494330 540988 494336 541000
rect 233200 540960 494336 540988
rect 233200 540948 233206 540960
rect 494330 540948 494336 540960
rect 494388 540948 494394 541000
rect 91094 540880 91100 540932
rect 91152 540920 91158 540932
rect 352006 540920 352012 540932
rect 91152 540892 352012 540920
rect 91152 540880 91158 540892
rect 352006 540880 352012 540892
rect 352064 540880 352070 540932
rect 121454 540812 121460 540864
rect 121512 540852 121518 540864
rect 349062 540852 349068 540864
rect 121512 540824 349068 540852
rect 121512 540812 121518 540824
rect 349062 540812 349068 540824
rect 349120 540812 349126 540864
rect 75822 540744 75828 540796
rect 75880 540784 75886 540796
rect 276842 540784 276848 540796
rect 75880 540756 276848 540784
rect 75880 540744 75886 540756
rect 276842 540744 276848 540756
rect 276900 540744 276906 540796
rect 272518 540676 272524 540728
rect 272576 540716 272582 540728
rect 317690 540716 317696 540728
rect 272576 540688 317696 540716
rect 272576 540676 272582 540688
rect 317690 540676 317696 540688
rect 317748 540676 317754 540728
rect 443638 540472 443644 540524
rect 443696 540512 443702 540524
rect 453298 540512 453304 540524
rect 443696 540484 453304 540512
rect 443696 540472 443702 540484
rect 453298 540472 453304 540484
rect 453356 540472 453362 540524
rect 208854 540404 208860 540456
rect 208912 540444 208918 540456
rect 487798 540444 487804 540456
rect 208912 540416 487804 540444
rect 208912 540404 208918 540416
rect 487798 540404 487804 540416
rect 487856 540404 487862 540456
rect 169018 540336 169024 540388
rect 169076 540376 169082 540388
rect 470962 540376 470968 540388
rect 169076 540348 470968 540376
rect 169076 540336 169082 540348
rect 470962 540336 470968 540348
rect 471020 540336 471026 540388
rect 177482 540268 177488 540320
rect 177540 540308 177546 540320
rect 493226 540308 493232 540320
rect 177540 540280 493232 540308
rect 177540 540268 177546 540280
rect 493226 540268 493232 540280
rect 493284 540268 493290 540320
rect 183554 540200 183560 540252
rect 183612 540240 183618 540252
rect 503898 540240 503904 540252
rect 183612 540212 503904 540240
rect 183612 540200 183618 540212
rect 503898 540200 503904 540212
rect 503956 540200 503962 540252
rect 86862 539520 86868 539572
rect 86920 539560 86926 539572
rect 373350 539560 373356 539572
rect 86920 539532 373356 539560
rect 86920 539520 86926 539532
rect 373350 539520 373356 539532
rect 373408 539520 373414 539572
rect 118694 539452 118700 539504
rect 118752 539492 118758 539504
rect 332870 539492 332876 539504
rect 118752 539464 332876 539492
rect 118752 539452 118758 539464
rect 332870 539452 332876 539464
rect 332928 539452 332934 539504
rect 131114 539384 131120 539436
rect 131172 539424 131178 539436
rect 316678 539424 316684 539436
rect 131172 539396 316684 539424
rect 131172 539384 131178 539396
rect 316678 539384 316684 539396
rect 316736 539384 316742 539436
rect 298738 539316 298744 539368
rect 298796 539356 298802 539368
rect 304258 539356 304264 539368
rect 298796 539328 304264 539356
rect 298796 539316 298802 539328
rect 304258 539316 304264 539328
rect 304316 539316 304322 539368
rect 138658 538976 138664 539028
rect 138716 539016 138722 539028
rect 372430 539016 372436 539028
rect 138716 538988 372436 539016
rect 138716 538976 138722 538988
rect 372430 538976 372436 538988
rect 372488 538976 372494 539028
rect 209866 538908 209872 538960
rect 209924 538948 209930 538960
rect 486050 538948 486056 538960
rect 209924 538920 486056 538948
rect 209924 538908 209930 538920
rect 486050 538908 486056 538920
rect 486108 538908 486114 538960
rect 194686 538840 194692 538892
rect 194744 538880 194750 538892
rect 480714 538880 480720 538892
rect 194744 538852 480720 538880
rect 194744 538840 194750 538852
rect 480714 538840 480720 538852
rect 480772 538840 480778 538892
rect 256694 538296 256700 538348
rect 256752 538336 256758 538348
rect 491478 538336 491484 538348
rect 256752 538308 491484 538336
rect 256752 538296 256758 538308
rect 491478 538296 491484 538308
rect 491536 538296 491542 538348
rect 171962 538228 171968 538280
rect 172020 538268 172026 538280
rect 447502 538268 447508 538280
rect 172020 538240 447508 538268
rect 172020 538228 172026 538240
rect 447502 538228 447508 538240
rect 447560 538228 447566 538280
rect 60826 538160 60832 538212
rect 60884 538200 60890 538212
rect 381078 538200 381084 538212
rect 60884 538172 381084 538200
rect 60884 538160 60890 538172
rect 381078 538160 381084 538172
rect 381136 538160 381142 538212
rect 82814 538092 82820 538144
rect 82872 538132 82878 538144
rect 370314 538132 370320 538144
rect 82872 538104 370320 538132
rect 82872 538092 82878 538104
rect 370314 538092 370320 538104
rect 370372 538092 370378 538144
rect 124122 538024 124128 538076
rect 124180 538064 124186 538076
rect 367278 538064 367284 538076
rect 124180 538036 367284 538064
rect 124180 538024 124186 538036
rect 367278 538024 367284 538036
rect 367336 538024 367342 538076
rect 171778 537956 171784 538008
rect 171836 537996 171842 538008
rect 331858 537996 331864 538008
rect 171836 537968 331864 537996
rect 171836 537956 171842 537968
rect 331858 537956 331864 537968
rect 331916 537956 331922 538008
rect 291838 537888 291844 537940
rect 291896 537928 291902 537940
rect 381630 537928 381636 537940
rect 291896 537900 381636 537928
rect 291896 537888 291902 537900
rect 381630 537888 381636 537900
rect 381688 537888 381694 537940
rect 252462 537820 252468 537872
rect 252520 537860 252526 537872
rect 315666 537860 315672 537872
rect 252520 537832 315672 537860
rect 252520 537820 252526 537832
rect 315666 537820 315672 537832
rect 315724 537820 315730 537872
rect 203794 537548 203800 537600
rect 203852 537588 203858 537600
rect 480990 537588 480996 537600
rect 203852 537560 480996 537588
rect 203852 537548 203858 537560
rect 480990 537548 480996 537560
rect 481048 537548 481054 537600
rect 195790 537480 195796 537532
rect 195848 537520 195854 537532
rect 480806 537520 480812 537532
rect 195848 537492 480812 537520
rect 195848 537480 195854 537492
rect 480806 537480 480812 537492
rect 480864 537480 480870 537532
rect 171042 536800 171048 536852
rect 171100 536840 171106 536852
rect 508130 536840 508136 536852
rect 171100 536812 508136 536840
rect 171100 536800 171106 536812
rect 508130 536800 508136 536812
rect 508188 536800 508194 536852
rect 97902 536732 97908 536784
rect 97960 536772 97966 536784
rect 344002 536772 344008 536784
rect 97960 536744 344008 536772
rect 97960 536732 97966 536744
rect 344002 536732 344008 536744
rect 344060 536732 344066 536784
rect 128354 536664 128360 536716
rect 128412 536704 128418 536716
rect 341978 536704 341984 536716
rect 128412 536676 341984 536704
rect 128412 536664 128418 536676
rect 341978 536664 341984 536676
rect 342036 536664 342042 536716
rect 178034 536596 178040 536648
rect 178092 536636 178098 536648
rect 330846 536636 330852 536648
rect 178092 536608 330852 536636
rect 178092 536596 178098 536608
rect 330846 536596 330852 536608
rect 330904 536596 330910 536648
rect 292574 536528 292580 536580
rect 292632 536568 292638 536580
rect 311618 536568 311624 536580
rect 292632 536540 311624 536568
rect 292632 536528 292638 536540
rect 311618 536528 311624 536540
rect 311676 536528 311682 536580
rect 179598 536052 179604 536104
rect 179656 536092 179662 536104
rect 506750 536092 506756 536104
rect 179656 536064 506756 536092
rect 179656 536052 179662 536064
rect 506750 536052 506756 536064
rect 506808 536052 506814 536104
rect 218054 535576 218060 535628
rect 218112 535616 218118 535628
rect 487890 535616 487896 535628
rect 218112 535588 487896 535616
rect 218112 535576 218118 535588
rect 487890 535576 487896 535588
rect 487948 535576 487954 535628
rect 173986 535508 173992 535560
rect 174044 535548 174050 535560
rect 463142 535548 463148 535560
rect 174044 535520 463148 535548
rect 174044 535508 174050 535520
rect 463142 535508 463148 535520
rect 463200 535508 463206 535560
rect 205634 535440 205640 535492
rect 205692 535480 205698 535492
rect 501138 535480 501144 535492
rect 205692 535452 501144 535480
rect 205692 535440 205698 535452
rect 501138 535440 501144 535452
rect 501196 535440 501202 535492
rect 97902 535372 97908 535424
rect 97960 535412 97966 535424
rect 358170 535412 358176 535424
rect 97960 535384 358176 535412
rect 97960 535372 97966 535384
rect 358170 535372 358176 535384
rect 358228 535372 358234 535424
rect 155862 535304 155868 535356
rect 155920 535344 155926 535356
rect 321738 535344 321744 535356
rect 155920 535316 321744 535344
rect 155920 535304 155926 535316
rect 321738 535304 321744 535316
rect 321796 535304 321802 535356
rect 179230 534760 179236 534812
rect 179288 534800 179294 534812
rect 461486 534800 461492 534812
rect 179288 534772 461492 534800
rect 179288 534760 179294 534772
rect 461486 534760 461492 534772
rect 461544 534760 461550 534812
rect 175182 534692 175188 534744
rect 175240 534732 175246 534744
rect 464706 534732 464712 534744
rect 175240 534704 464712 534732
rect 175240 534692 175246 534704
rect 464706 534692 464712 534704
rect 464764 534692 464770 534744
rect 243538 534284 243544 534336
rect 243596 534324 243602 534336
rect 487982 534324 487988 534336
rect 243596 534296 487988 534324
rect 243596 534284 243602 534296
rect 487982 534284 487988 534296
rect 488040 534284 488046 534336
rect 164142 534216 164148 534268
rect 164200 534256 164206 534268
rect 427078 534256 427084 534268
rect 164200 534228 427084 534256
rect 164200 534216 164206 534228
rect 427078 534216 427084 534228
rect 427136 534216 427142 534268
rect 212442 534148 212448 534200
rect 212500 534188 212506 534200
rect 480898 534188 480904 534200
rect 212500 534160 480904 534188
rect 212500 534148 212506 534160
rect 480898 534148 480904 534160
rect 480956 534148 480962 534200
rect 70486 534080 70492 534132
rect 70544 534120 70550 534132
rect 72418 534120 72424 534132
rect 70544 534092 72424 534120
rect 70544 534080 70550 534092
rect 72418 534080 72424 534092
rect 72476 534080 72482 534132
rect 194502 534080 194508 534132
rect 194560 534120 194566 534132
rect 500954 534120 500960 534132
rect 194560 534092 500960 534120
rect 194560 534080 194566 534092
rect 500954 534080 500960 534092
rect 501012 534080 501018 534132
rect 60734 534012 60740 534064
rect 60792 534052 60798 534064
rect 369302 534052 369308 534064
rect 60792 534024 369308 534052
rect 60792 534012 60798 534024
rect 369302 534012 369308 534024
rect 369360 534012 369366 534064
rect 70394 533944 70400 533996
rect 70452 533984 70458 533996
rect 354122 533984 354128 533996
rect 70452 533956 354128 533984
rect 70452 533944 70458 533956
rect 354122 533944 354128 533956
rect 354180 533944 354186 533996
rect 59170 533876 59176 533928
rect 59228 533916 59234 533928
rect 280890 533916 280896 533928
rect 59228 533888 280896 533916
rect 59228 533876 59234 533888
rect 280890 533876 280896 533888
rect 280948 533876 280954 533928
rect 166994 533808 167000 533860
rect 167052 533848 167058 533860
rect 338942 533848 338948 533860
rect 167052 533820 338948 533848
rect 167052 533808 167058 533820
rect 338942 533808 338948 533820
rect 339000 533808 339006 533860
rect 175826 533740 175832 533792
rect 175884 533780 175890 533792
rect 327810 533780 327816 533792
rect 175884 533752 327816 533780
rect 175884 533740 175890 533752
rect 327810 533740 327816 533752
rect 327868 533740 327874 533792
rect 177574 533400 177580 533452
rect 177632 533400 177638 533452
rect 177592 533372 177620 533400
rect 491754 533372 491760 533384
rect 177592 533344 491760 533372
rect 491754 533332 491760 533344
rect 491812 533332 491818 533384
rect 67910 532788 67916 532840
rect 67968 532828 67974 532840
rect 71038 532828 71044 532840
rect 67968 532800 71044 532828
rect 67968 532788 67974 532800
rect 71038 532788 71044 532800
rect 71096 532788 71102 532840
rect 244366 532788 244372 532840
rect 244424 532828 244430 532840
rect 502426 532828 502432 532840
rect 244424 532800 502432 532828
rect 244424 532788 244430 532800
rect 502426 532788 502432 532800
rect 502484 532788 502490 532840
rect 191742 532720 191748 532772
rect 191800 532760 191806 532772
rect 493502 532760 493508 532772
rect 191800 532732 493508 532760
rect 191800 532720 191806 532732
rect 493502 532720 493508 532732
rect 493560 532720 493566 532772
rect 96522 532652 96528 532704
rect 96580 532692 96586 532704
rect 368290 532692 368296 532704
rect 96580 532664 368296 532692
rect 96580 532652 96586 532664
rect 368290 532652 368296 532664
rect 368348 532652 368354 532704
rect 117222 532584 117228 532636
rect 117280 532624 117286 532636
rect 340966 532624 340972 532636
rect 117280 532596 340972 532624
rect 117280 532584 117286 532596
rect 340966 532584 340972 532596
rect 341024 532584 341030 532636
rect 131114 532516 131120 532568
rect 131172 532556 131178 532568
rect 329834 532556 329840 532568
rect 131172 532528 329840 532556
rect 131172 532516 131178 532528
rect 329834 532516 329840 532528
rect 329892 532516 329898 532568
rect 178034 532448 178040 532500
rect 178092 532488 178098 532500
rect 285030 532488 285036 532500
rect 178092 532460 285036 532488
rect 178092 532448 178098 532460
rect 285030 532448 285036 532460
rect 285088 532448 285094 532500
rect 290458 532176 290464 532228
rect 290516 532216 290522 532228
rect 330202 532216 330208 532228
rect 290516 532188 330208 532216
rect 290516 532176 290522 532188
rect 330202 532176 330208 532188
rect 330260 532176 330266 532228
rect 178862 532108 178868 532160
rect 178920 532148 178926 532160
rect 403710 532148 403716 532160
rect 178920 532120 403716 532148
rect 178920 532108 178926 532120
rect 403710 532108 403716 532120
rect 403768 532108 403774 532160
rect 178678 532040 178684 532092
rect 178736 532080 178742 532092
rect 450630 532080 450636 532092
rect 178736 532052 450636 532080
rect 178736 532040 178742 532052
rect 450630 532040 450636 532052
rect 450688 532040 450694 532092
rect 174630 531972 174636 532024
rect 174688 532012 174694 532024
rect 455322 532012 455328 532024
rect 174688 531984 455328 532012
rect 174688 531972 174694 531984
rect 455322 531972 455328 531984
rect 455380 531972 455386 532024
rect 213822 531292 213828 531344
rect 213880 531332 213886 531344
rect 494146 531332 494152 531344
rect 213880 531304 494152 531332
rect 213880 531292 213886 531304
rect 494146 531292 494152 531304
rect 494204 531292 494210 531344
rect 59906 531224 59912 531276
rect 59964 531264 59970 531276
rect 366266 531264 366272 531276
rect 59964 531236 366272 531264
rect 59964 531224 59970 531236
rect 366266 531224 366272 531236
rect 366324 531224 366330 531276
rect 67542 531156 67548 531208
rect 67600 531196 67606 531208
rect 355134 531196 355140 531208
rect 67600 531168 355140 531196
rect 67600 531156 67606 531168
rect 355134 531156 355140 531168
rect 355192 531156 355198 531208
rect 111794 531088 111800 531140
rect 111852 531128 111858 531140
rect 335906 531128 335912 531140
rect 111852 531100 335912 531128
rect 111852 531088 111858 531100
rect 335906 531088 335912 531100
rect 335964 531088 335970 531140
rect 59170 531020 59176 531072
rect 59228 531060 59234 531072
rect 278130 531060 278136 531072
rect 59228 531032 278136 531060
rect 59228 531020 59234 531032
rect 278130 531020 278136 531032
rect 278188 531020 278194 531072
rect 211062 530952 211068 531004
rect 211120 530992 211126 531004
rect 337930 530992 337936 531004
rect 211120 530964 337936 530992
rect 211120 530952 211126 530964
rect 337930 530952 337936 530964
rect 337988 530952 337994 531004
rect 64782 530544 64788 530596
rect 64840 530584 64846 530596
rect 67910 530584 67916 530596
rect 64840 530556 67916 530584
rect 64840 530544 64846 530556
rect 67910 530544 67916 530556
rect 67968 530544 67974 530596
rect 113174 530544 113180 530596
rect 113232 530584 113238 530596
rect 124858 530584 124864 530596
rect 113232 530556 124864 530584
rect 113232 530544 113238 530556
rect 124858 530544 124864 530556
rect 124916 530544 124922 530596
rect 177666 530544 177672 530596
rect 177724 530584 177730 530596
rect 489270 530584 489276 530596
rect 177724 530556 489276 530584
rect 177724 530544 177730 530556
rect 489270 530544 489276 530556
rect 489328 530544 489334 530596
rect 295334 530068 295340 530120
rect 295392 530108 295398 530120
rect 497182 530108 497188 530120
rect 295392 530080 497188 530108
rect 295392 530068 295398 530080
rect 497182 530068 497188 530080
rect 497240 530068 497246 530120
rect 289722 530000 289728 530052
rect 289780 530040 289786 530052
rect 497090 530040 497096 530052
rect 289780 530012 497096 530040
rect 289780 530000 289786 530012
rect 497090 530000 497096 530012
rect 497148 530000 497154 530052
rect 251082 529932 251088 529984
rect 251140 529972 251146 529984
rect 479610 529972 479616 529984
rect 251140 529944 479616 529972
rect 251140 529932 251146 529944
rect 479610 529932 479616 529944
rect 479668 529932 479674 529984
rect 59446 529864 59452 529916
rect 59504 529904 59510 529916
rect 378226 529904 378232 529916
rect 59504 529876 378232 529904
rect 59504 529864 59510 529876
rect 378226 529864 378232 529876
rect 378284 529864 378290 529916
rect 59170 529796 59176 529848
rect 59228 529836 59234 529848
rect 363230 529836 363236 529848
rect 59228 529808 363236 529836
rect 59228 529796 59234 529808
rect 363230 529796 363236 529808
rect 363288 529796 363294 529848
rect 68646 529728 68652 529780
rect 68704 529768 68710 529780
rect 70302 529768 70308 529780
rect 68704 529740 70308 529768
rect 68704 529728 68710 529740
rect 70302 529728 70308 529740
rect 70360 529728 70366 529780
rect 127618 529728 127624 529780
rect 127676 529768 127682 529780
rect 375374 529768 375380 529780
rect 127676 529740 375380 529768
rect 127676 529728 127682 529740
rect 375374 529728 375380 529740
rect 375432 529728 375438 529780
rect 135162 529660 135168 529712
rect 135220 529700 135226 529712
rect 378318 529700 378324 529712
rect 135220 529672 378324 529700
rect 135220 529660 135226 529672
rect 378318 529660 378324 529672
rect 378376 529660 378382 529712
rect 166258 529592 166264 529644
rect 166316 529632 166322 529644
rect 374546 529632 374552 529644
rect 166316 529604 374552 529632
rect 166316 529592 166322 529604
rect 374546 529592 374552 529604
rect 374604 529592 374610 529644
rect 181530 529184 181536 529236
rect 181588 529224 181594 529236
rect 501046 529224 501052 529236
rect 181588 529196 501052 529224
rect 181588 529184 181594 529196
rect 501046 529184 501052 529196
rect 501104 529184 501110 529236
rect 289722 528640 289728 528692
rect 289780 528680 289786 528692
rect 499850 528680 499856 528692
rect 289780 528652 499856 528680
rect 289780 528640 289786 528652
rect 499850 528640 499856 528652
rect 499908 528640 499914 528692
rect 177482 528572 177488 528624
rect 177540 528612 177546 528624
rect 493318 528612 493324 528624
rect 177540 528584 493324 528612
rect 177540 528572 177546 528584
rect 493318 528572 493324 528584
rect 493376 528572 493382 528624
rect 175826 528504 175832 528556
rect 175884 528544 175890 528556
rect 378410 528544 378416 528556
rect 175884 528516 378416 528544
rect 175884 528504 175890 528516
rect 378410 528504 378416 528516
rect 378468 528504 378474 528556
rect 175182 528436 175188 528488
rect 175240 528476 175246 528488
rect 374730 528476 374736 528488
rect 175240 528448 374736 528476
rect 175240 528436 175246 528448
rect 374730 528436 374736 528448
rect 374788 528436 374794 528488
rect 220630 528368 220636 528420
rect 220688 528408 220694 528420
rect 378594 528408 378600 528420
rect 220688 528380 378600 528408
rect 220688 528368 220694 528380
rect 378594 528368 378600 528380
rect 378652 528368 378658 528420
rect 279970 528300 279976 528352
rect 280028 528340 280034 528352
rect 375834 528340 375840 528352
rect 280028 528312 375840 528340
rect 280028 528300 280034 528312
rect 375834 528300 375840 528312
rect 375892 528300 375898 528352
rect 92474 527892 92480 527944
rect 92532 527932 92538 527944
rect 113174 527932 113180 527944
rect 92532 527904 113180 527932
rect 92532 527892 92538 527904
rect 113174 527892 113180 527904
rect 113232 527892 113238 527944
rect 60366 527824 60372 527876
rect 60424 527864 60430 527876
rect 155218 527864 155224 527876
rect 60424 527836 155224 527864
rect 60424 527824 60430 527836
rect 155218 527824 155224 527836
rect 155276 527824 155282 527876
rect 186590 527824 186596 527876
rect 186648 527864 186654 527876
rect 498286 527864 498292 527876
rect 186648 527836 498292 527864
rect 186648 527824 186654 527836
rect 498286 527824 498292 527836
rect 498344 527824 498350 527876
rect 286318 527212 286324 527264
rect 286376 527252 286382 527264
rect 497274 527252 497280 527264
rect 286376 527224 497280 527252
rect 286376 527212 286382 527224
rect 497274 527212 497280 527224
rect 497332 527212 497338 527264
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 60366 527184 60372 527196
rect 3476 527156 60372 527184
rect 3476 527144 3482 527156
rect 60366 527144 60372 527156
rect 60424 527144 60430 527196
rect 62206 527144 62212 527196
rect 62264 527184 62270 527196
rect 64782 527184 64788 527196
rect 62264 527156 64788 527184
rect 62264 527144 62270 527156
rect 64782 527144 64788 527156
rect 64840 527144 64846 527196
rect 66162 527144 66168 527196
rect 66220 527184 66226 527196
rect 68646 527184 68652 527196
rect 66220 527156 68652 527184
rect 66220 527144 66226 527156
rect 68646 527144 68652 527156
rect 68704 527144 68710 527196
rect 169754 527144 169760 527196
rect 169812 527184 169818 527196
rect 472526 527184 472532 527196
rect 169812 527156 472532 527184
rect 169812 527144 169818 527156
rect 472526 527144 472532 527156
rect 472584 527144 472590 527196
rect 108298 527076 108304 527128
rect 108356 527116 108362 527128
rect 372154 527116 372160 527128
rect 108356 527088 372160 527116
rect 108356 527076 108362 527088
rect 372154 527076 372160 527088
rect 372212 527076 372218 527128
rect 107562 527008 107568 527060
rect 107620 527048 107626 527060
rect 333882 527048 333888 527060
rect 107620 527020 333888 527048
rect 107620 527008 107626 527020
rect 333882 527008 333888 527020
rect 333940 527008 333946 527060
rect 109034 526940 109040 526992
rect 109092 526980 109098 526992
rect 312630 526980 312636 526992
rect 109092 526952 312636 526980
rect 109092 526940 109098 526952
rect 312630 526940 312636 526952
rect 312688 526940 312694 526992
rect 109126 526872 109132 526924
rect 109184 526912 109190 526924
rect 283650 526912 283656 526924
rect 109184 526884 283656 526912
rect 109184 526872 109190 526884
rect 283650 526872 283656 526884
rect 283708 526872 283714 526924
rect 111058 526464 111064 526516
rect 111116 526504 111122 526516
rect 211338 526504 211344 526516
rect 111116 526476 211344 526504
rect 111116 526464 111122 526476
rect 211338 526464 211344 526476
rect 211396 526464 211402 526516
rect 255406 526464 255412 526516
rect 255464 526504 255470 526516
rect 283742 526504 283748 526516
rect 255464 526476 283748 526504
rect 255464 526464 255470 526476
rect 283742 526464 283748 526476
rect 283800 526464 283806 526516
rect 175918 526396 175924 526448
rect 175976 526436 175982 526448
rect 433426 526436 433432 526448
rect 175976 526408 433432 526436
rect 175976 526396 175982 526408
rect 433426 526396 433432 526408
rect 433484 526396 433490 526448
rect 453298 526396 453304 526448
rect 453356 526436 453362 526448
rect 463602 526436 463608 526448
rect 453356 526408 463608 526436
rect 453356 526396 453362 526408
rect 463602 526396 463608 526408
rect 463660 526396 463666 526448
rect 66162 525960 66168 525972
rect 64846 525932 66168 525960
rect 62850 525716 62856 525768
rect 62908 525756 62914 525768
rect 64846 525756 64874 525932
rect 66162 525920 66168 525932
rect 66220 525920 66226 525972
rect 300762 525920 300768 525972
rect 300820 525960 300826 525972
rect 499666 525960 499672 525972
rect 300820 525932 499672 525960
rect 300820 525920 300826 525932
rect 499666 525920 499672 525932
rect 499724 525920 499730 525972
rect 289722 525852 289728 525904
rect 289780 525892 289786 525904
rect 498470 525892 498476 525904
rect 289780 525864 498476 525892
rect 289780 525852 289786 525864
rect 498470 525852 498476 525864
rect 498528 525852 498534 525904
rect 172422 525784 172428 525836
rect 172480 525824 172486 525836
rect 505186 525824 505192 525836
rect 172480 525796 505192 525824
rect 172480 525784 172486 525796
rect 505186 525784 505192 525796
rect 505244 525784 505250 525836
rect 62908 525728 64874 525756
rect 62908 525716 62914 525728
rect 100754 525716 100760 525768
rect 100812 525756 100818 525768
rect 379514 525756 379520 525768
rect 100812 525728 379520 525756
rect 100812 525716 100818 525728
rect 379514 525716 379520 525728
rect 379572 525716 379578 525768
rect 120074 525648 120080 525700
rect 120132 525688 120138 525700
rect 351086 525688 351092 525700
rect 120132 525660 351092 525688
rect 120132 525648 120138 525660
rect 351086 525648 351092 525660
rect 351144 525648 351150 525700
rect 175918 525580 175924 525632
rect 175976 525620 175982 525632
rect 386690 525620 386696 525632
rect 175976 525592 386696 525620
rect 175976 525580 175982 525592
rect 386690 525580 386696 525592
rect 386748 525580 386754 525632
rect 133782 525512 133788 525564
rect 133840 525552 133846 525564
rect 325786 525552 325792 525564
rect 133840 525524 325792 525552
rect 133840 525512 133846 525524
rect 325786 525512 325792 525524
rect 325844 525512 325850 525564
rect 102134 525444 102140 525496
rect 102192 525484 102198 525496
rect 274082 525484 274088 525496
rect 102192 525456 274088 525484
rect 102192 525444 102198 525456
rect 274082 525444 274088 525456
rect 274140 525444 274146 525496
rect 299382 525444 299388 525496
rect 299440 525484 299446 525496
rect 372062 525484 372068 525496
rect 299440 525456 372068 525484
rect 299440 525444 299446 525456
rect 372062 525444 372068 525456
rect 372120 525444 372126 525496
rect 118694 525376 118700 525428
rect 118752 525416 118758 525428
rect 274174 525416 274180 525428
rect 118752 525388 274180 525416
rect 118752 525376 118758 525388
rect 274174 525376 274180 525388
rect 274232 525376 274238 525428
rect 255314 525036 255320 525088
rect 255372 525076 255378 525088
rect 298738 525076 298744 525088
rect 255372 525048 298744 525076
rect 255372 525036 255378 525048
rect 298738 525036 298744 525048
rect 298796 525036 298802 525088
rect 465810 525036 465816 525088
rect 465868 525076 465874 525088
rect 513374 525076 513380 525088
rect 465868 525048 513380 525076
rect 465868 525036 465874 525048
rect 513374 525036 513380 525048
rect 513432 525036 513438 525088
rect 180242 524492 180248 524544
rect 180300 524532 180306 524544
rect 508222 524532 508228 524544
rect 180300 524504 508228 524532
rect 180300 524492 180306 524504
rect 508222 524492 508228 524504
rect 508280 524492 508286 524544
rect 55766 524424 55772 524476
rect 55824 524464 55830 524476
rect 58618 524464 58624 524476
rect 55824 524436 58624 524464
rect 55824 524424 55830 524436
rect 58618 524424 58624 524436
rect 58676 524424 58682 524476
rect 175182 524424 175188 524476
rect 175240 524464 175246 524476
rect 506842 524464 506848 524476
rect 175240 524436 506848 524464
rect 175240 524424 175246 524436
rect 506842 524424 506848 524436
rect 506900 524424 506906 524476
rect 59170 524356 59176 524408
rect 59228 524396 59234 524408
rect 380986 524396 380992 524408
rect 59228 524368 380992 524396
rect 59228 524356 59234 524368
rect 380986 524356 380992 524368
rect 381044 524356 381050 524408
rect 63494 524288 63500 524340
rect 63552 524328 63558 524340
rect 378134 524328 378140 524340
rect 63552 524300 378140 524328
rect 63552 524288 63558 524300
rect 378134 524288 378140 524300
rect 378192 524288 378198 524340
rect 66162 524220 66168 524272
rect 66220 524260 66226 524272
rect 375466 524260 375472 524272
rect 66220 524232 375472 524260
rect 66220 524220 66226 524232
rect 375466 524220 375472 524232
rect 375524 524220 375530 524272
rect 69658 524152 69664 524204
rect 69716 524192 69722 524204
rect 375742 524192 375748 524204
rect 69716 524164 375748 524192
rect 69716 524152 69722 524164
rect 375742 524152 375748 524164
rect 375800 524152 375806 524204
rect 169754 524084 169760 524136
rect 169812 524124 169818 524136
rect 383930 524124 383936 524136
rect 169812 524096 383936 524124
rect 169812 524084 169818 524096
rect 383930 524084 383936 524096
rect 383988 524084 383994 524136
rect 178034 524016 178040 524068
rect 178092 524056 178098 524068
rect 382366 524056 382372 524068
rect 178092 524028 382372 524056
rect 178092 524016 178098 524028
rect 382366 524016 382372 524028
rect 382424 524016 382430 524068
rect 274634 523948 274640 524000
rect 274692 523988 274698 524000
rect 297358 523988 297364 524000
rect 274692 523960 297364 523988
rect 274692 523948 274698 523960
rect 297358 523948 297364 523960
rect 297416 523948 297422 524000
rect 299382 523744 299388 523796
rect 299440 523784 299446 523796
rect 481634 523784 481640 523796
rect 299440 523756 481640 523784
rect 299440 523744 299446 523756
rect 481634 523744 481640 523756
rect 481692 523744 481698 523796
rect 86862 522996 86868 523048
rect 86920 523036 86926 523048
rect 92474 523036 92480 523048
rect 86920 523008 92480 523036
rect 86920 522996 86926 523008
rect 92474 522996 92480 523008
rect 92532 522996 92538 523048
rect 292574 522996 292580 523048
rect 292632 523036 292638 523048
rect 312998 523036 313004 523048
rect 292632 523008 313004 523036
rect 292632 522996 292638 523008
rect 312998 522996 313004 523008
rect 313056 522996 313062 523048
rect 56502 522928 56508 522980
rect 56560 522968 56566 522980
rect 386598 522968 386604 522980
rect 56560 522940 386604 522968
rect 56560 522928 56566 522940
rect 386598 522928 386604 522940
rect 386656 522928 386662 522980
rect 463602 522928 463608 522980
rect 463660 522968 463666 522980
rect 467834 522968 467840 522980
rect 463660 522940 467840 522968
rect 463660 522928 463666 522940
rect 467834 522928 467840 522940
rect 467892 522928 467898 522980
rect 63494 522860 63500 522912
rect 63552 522900 63558 522912
rect 385402 522900 385408 522912
rect 63552 522872 385408 522900
rect 63552 522860 63558 522872
rect 385402 522860 385408 522872
rect 385460 522860 385466 522912
rect 59906 522792 59912 522844
rect 59964 522832 59970 522844
rect 375558 522832 375564 522844
rect 59964 522804 375564 522832
rect 59964 522792 59970 522804
rect 375558 522792 375564 522804
rect 375616 522792 375622 522844
rect 62114 522724 62120 522776
rect 62172 522764 62178 522776
rect 378502 522764 378508 522776
rect 62172 522736 378508 522764
rect 62172 522724 62178 522736
rect 378502 522724 378508 522736
rect 378560 522724 378566 522776
rect 80054 522656 80060 522708
rect 80112 522696 80118 522708
rect 371970 522696 371976 522708
rect 80112 522668 371976 522696
rect 80112 522656 80118 522668
rect 371970 522656 371976 522668
rect 372028 522656 372034 522708
rect 114462 522588 114468 522640
rect 114520 522628 114526 522640
rect 382550 522628 382556 522640
rect 114520 522600 382556 522628
rect 114520 522588 114526 522600
rect 382550 522588 382556 522600
rect 382608 522588 382614 522640
rect 477402 522588 477408 522640
rect 477460 522628 477466 522640
rect 503714 522628 503720 522640
rect 477460 522600 503720 522628
rect 477460 522588 477466 522600
rect 503714 522588 503720 522600
rect 503772 522588 503778 522640
rect 474274 522520 474280 522572
rect 474332 522560 474338 522572
rect 504174 522560 504180 522572
rect 474332 522532 504180 522560
rect 474332 522520 474338 522532
rect 504174 522520 504180 522532
rect 504232 522520 504238 522572
rect 475930 522452 475936 522504
rect 475988 522492 475994 522504
rect 506566 522492 506572 522504
rect 475988 522464 506572 522492
rect 475988 522452 475994 522464
rect 506566 522452 506572 522464
rect 506624 522452 506630 522504
rect 465718 522384 465724 522436
rect 465776 522424 465782 522436
rect 497550 522424 497556 522436
rect 465776 522396 497556 522424
rect 465776 522384 465782 522396
rect 497550 522384 497556 522396
rect 497608 522384 497614 522436
rect 464430 522316 464436 522368
rect 464488 522356 464494 522368
rect 502610 522356 502616 522368
rect 464488 522328 502616 522356
rect 464488 522316 464494 522328
rect 502610 522316 502616 522328
rect 502668 522316 502674 522368
rect 468754 522248 468760 522300
rect 468812 522288 468818 522300
rect 510614 522288 510620 522300
rect 468812 522260 510620 522288
rect 468812 522248 468818 522260
rect 510614 522248 510620 522260
rect 510672 522248 510678 522300
rect 471882 521704 471888 521756
rect 471940 521744 471946 521756
rect 490558 521744 490564 521756
rect 471940 521716 490564 521744
rect 471940 521704 471946 521716
rect 490558 521704 490564 521716
rect 490616 521704 490622 521756
rect 293954 521636 293960 521688
rect 294012 521676 294018 521688
rect 494514 521676 494520 521688
rect 294012 521648 494520 521676
rect 294012 521636 294018 521648
rect 494514 521636 494520 521648
rect 494572 521636 494578 521688
rect 60734 521568 60740 521620
rect 60792 521608 60798 521620
rect 62206 521608 62212 521620
rect 60792 521580 62212 521608
rect 60792 521568 60798 521580
rect 62206 521568 62212 521580
rect 62264 521568 62270 521620
rect 99374 521568 99380 521620
rect 99432 521608 99438 521620
rect 385126 521608 385132 521620
rect 99432 521580 385132 521608
rect 99432 521568 99438 521580
rect 385126 521568 385132 521580
rect 385184 521568 385190 521620
rect 60826 521500 60832 521552
rect 60884 521540 60890 521552
rect 62850 521540 62856 521552
rect 60884 521512 62856 521540
rect 60884 521500 60890 521512
rect 62850 521500 62856 521512
rect 62908 521500 62914 521552
rect 110414 521500 110420 521552
rect 110472 521540 110478 521552
rect 383654 521540 383660 521552
rect 110472 521512 383660 521540
rect 110472 521500 110478 521512
rect 383654 521500 383660 521512
rect 383712 521500 383718 521552
rect 114462 521432 114468 521484
rect 114520 521472 114526 521484
rect 385310 521472 385316 521484
rect 114520 521444 385316 521472
rect 114520 521432 114526 521444
rect 385310 521432 385316 521444
rect 385368 521432 385374 521484
rect 115750 521364 115756 521416
rect 115808 521404 115814 521416
rect 382458 521404 382464 521416
rect 115808 521376 382464 521404
rect 115808 521364 115814 521376
rect 382458 521364 382464 521376
rect 382516 521364 382522 521416
rect 117222 521296 117228 521348
rect 117280 521336 117286 521348
rect 301498 521336 301504 521348
rect 117280 521308 301504 521336
rect 117280 521296 117286 521308
rect 301498 521296 301504 521308
rect 301556 521296 301562 521348
rect 253290 521228 253296 521280
rect 253348 521268 253354 521280
rect 256602 521268 256608 521280
rect 253348 521240 256608 521268
rect 253348 521228 253354 521240
rect 256602 521228 256608 521240
rect 256660 521228 256666 521280
rect 471330 521228 471336 521280
rect 471388 521268 471394 521280
rect 504266 521268 504272 521280
rect 471388 521240 504272 521268
rect 471388 521228 471394 521240
rect 504266 521228 504272 521240
rect 504324 521228 504330 521280
rect 254578 521160 254584 521212
rect 254636 521200 254642 521212
rect 276934 521200 276940 521212
rect 254636 521172 276940 521200
rect 254636 521160 254642 521172
rect 276934 521160 276940 521172
rect 276992 521160 276998 521212
rect 468478 521160 468484 521212
rect 468536 521200 468542 521212
rect 505370 521200 505376 521212
rect 468536 521172 505376 521200
rect 468536 521160 468542 521172
rect 505370 521160 505376 521172
rect 505428 521160 505434 521212
rect 61930 521092 61936 521144
rect 61988 521132 61994 521144
rect 86862 521132 86868 521144
rect 61988 521104 86868 521132
rect 61988 521092 61994 521104
rect 86862 521092 86868 521104
rect 86920 521092 86926 521144
rect 216122 521092 216128 521144
rect 216180 521132 216186 521144
rect 281534 521132 281540 521144
rect 216180 521104 281540 521132
rect 216180 521092 216186 521104
rect 281534 521092 281540 521104
rect 281592 521092 281598 521144
rect 295978 521092 295984 521144
rect 296036 521132 296042 521144
rect 367554 521132 367560 521144
rect 296036 521104 367560 521132
rect 296036 521092 296042 521104
rect 367554 521092 367560 521104
rect 367612 521092 367618 521144
rect 468662 521092 468668 521144
rect 468720 521132 468726 521144
rect 512178 521132 512184 521144
rect 468720 521104 512184 521132
rect 468720 521092 468726 521104
rect 512178 521092 512184 521104
rect 512236 521092 512242 521144
rect 62022 521024 62028 521076
rect 62080 521064 62086 521076
rect 255406 521064 255412 521076
rect 62080 521036 255412 521064
rect 62080 521024 62086 521036
rect 255406 521024 255412 521036
rect 255464 521024 255470 521076
rect 289078 521024 289084 521076
rect 289136 521064 289142 521076
rect 366082 521064 366088 521076
rect 289136 521036 366088 521064
rect 289136 521024 289142 521036
rect 366082 521024 366088 521036
rect 366140 521024 366146 521076
rect 461762 521024 461768 521076
rect 461820 521064 461826 521076
rect 505278 521064 505284 521076
rect 461820 521036 505284 521064
rect 461820 521024 461826 521036
rect 505278 521024 505284 521036
rect 505336 521024 505342 521076
rect 58802 520956 58808 521008
rect 58860 520996 58866 521008
rect 255314 520996 255320 521008
rect 58860 520968 255320 520996
rect 58860 520956 58866 520968
rect 255314 520956 255320 520968
rect 255372 520956 255378 521008
rect 264238 520956 264244 521008
rect 264296 520996 264302 521008
rect 370774 520996 370780 521008
rect 264296 520968 370780 520996
rect 264296 520956 264302 520968
rect 370774 520956 370780 520968
rect 370832 520956 370838 521008
rect 373902 520956 373908 521008
rect 373960 520996 373966 521008
rect 381538 520996 381544 521008
rect 373960 520968 381544 520996
rect 373960 520956 373966 520968
rect 381538 520956 381544 520968
rect 381596 520956 381602 521008
rect 427078 520956 427084 521008
rect 427136 520996 427142 521008
rect 475470 520996 475476 521008
rect 427136 520968 475476 520996
rect 427136 520956 427142 520968
rect 475470 520956 475476 520968
rect 475528 520956 475534 521008
rect 68278 520888 68284 520940
rect 68336 520928 68342 520940
rect 294138 520928 294144 520940
rect 68336 520900 294144 520928
rect 68336 520888 68342 520900
rect 294138 520888 294144 520900
rect 294196 520888 294202 520940
rect 360838 520888 360844 520940
rect 360896 520928 360902 520940
rect 473998 520928 474004 520940
rect 360896 520900 474004 520928
rect 360896 520888 360902 520900
rect 473998 520888 474004 520900
rect 474056 520888 474062 520940
rect 258442 520276 258448 520328
rect 258500 520316 258506 520328
rect 431678 520316 431684 520328
rect 258500 520288 431684 520316
rect 258500 520276 258506 520288
rect 431678 520276 431684 520288
rect 431736 520276 431742 520328
rect 55122 520208 55128 520260
rect 55180 520248 55186 520260
rect 137830 520248 137836 520260
rect 55180 520220 137836 520248
rect 55180 520208 55186 520220
rect 137830 520208 137836 520220
rect 137888 520208 137894 520260
rect 475378 520208 475384 520260
rect 475436 520248 475442 520260
rect 479702 520248 479708 520260
rect 475436 520220 479708 520248
rect 475436 520208 475442 520220
rect 479702 520208 479708 520220
rect 479760 520208 479766 520260
rect 45922 520140 45928 520192
rect 45980 520180 45986 520192
rect 289170 520180 289176 520192
rect 45980 520152 289176 520180
rect 45980 520140 45986 520152
rect 289170 520140 289176 520152
rect 289228 520140 289234 520192
rect 291010 520140 291016 520192
rect 291068 520180 291074 520192
rect 383746 520180 383752 520192
rect 291068 520152 383752 520180
rect 291068 520140 291074 520152
rect 383746 520140 383752 520152
rect 383804 520140 383810 520192
rect 44174 520072 44180 520124
rect 44232 520112 44238 520124
rect 44232 520084 277394 520112
rect 44232 520072 44238 520084
rect 50154 520004 50160 520056
rect 50212 520044 50218 520056
rect 275370 520044 275376 520056
rect 50212 520016 275376 520044
rect 50212 520004 50218 520016
rect 275370 520004 275376 520016
rect 275428 520004 275434 520056
rect 277366 520044 277394 520084
rect 282914 520072 282920 520124
rect 282972 520112 282978 520124
rect 371878 520112 371884 520124
rect 282972 520084 371884 520112
rect 282972 520072 282978 520084
rect 371878 520072 371884 520084
rect 371936 520072 371942 520124
rect 283558 520044 283564 520056
rect 277366 520016 283564 520044
rect 283558 520004 283564 520016
rect 283616 520004 283622 520056
rect 467834 520004 467840 520056
rect 467892 520044 467898 520056
rect 480162 520044 480168 520056
rect 467892 520016 480168 520044
rect 467892 520004 467898 520016
rect 480162 520004 480168 520016
rect 480220 520004 480226 520056
rect 57698 519936 57704 519988
rect 57756 519976 57762 519988
rect 271138 519976 271144 519988
rect 57756 519948 271144 519976
rect 57756 519936 57762 519948
rect 271138 519936 271144 519948
rect 271196 519936 271202 519988
rect 476022 519936 476028 519988
rect 476080 519976 476086 519988
rect 494882 519976 494888 519988
rect 476080 519948 494888 519976
rect 476080 519936 476086 519948
rect 494882 519936 494888 519948
rect 494940 519936 494946 519988
rect 270402 519868 270408 519920
rect 270460 519908 270466 519920
rect 385034 519908 385040 519920
rect 270460 519880 385040 519908
rect 270460 519868 270466 519880
rect 385034 519868 385040 519880
rect 385092 519868 385098 519920
rect 471238 519868 471244 519920
rect 471296 519908 471302 519920
rect 494698 519908 494704 519920
rect 471296 519880 494704 519908
rect 471296 519868 471302 519880
rect 494698 519868 494704 519880
rect 494756 519868 494762 519920
rect 164142 519800 164148 519852
rect 164200 519840 164206 519852
rect 273990 519840 273996 519852
rect 164200 519812 273996 519840
rect 164200 519800 164206 519812
rect 273990 519800 273996 519812
rect 274048 519800 274054 519852
rect 471422 519800 471428 519852
rect 471480 519840 471486 519852
rect 495894 519840 495900 519852
rect 471480 519812 495900 519840
rect 471480 519800 471486 519812
rect 495894 519800 495900 519812
rect 495952 519800 495958 519852
rect 467282 519732 467288 519784
rect 467340 519772 467346 519784
rect 498654 519772 498660 519784
rect 467340 519744 498660 519772
rect 467340 519732 467346 519744
rect 498654 519732 498660 519744
rect 498712 519732 498718 519784
rect 56134 519664 56140 519716
rect 56192 519704 56198 519716
rect 138014 519704 138020 519716
rect 56192 519676 138020 519704
rect 56192 519664 56198 519676
rect 138014 519664 138020 519676
rect 138072 519664 138078 519716
rect 467190 519664 467196 519716
rect 467248 519704 467254 519716
rect 500034 519704 500040 519716
rect 467248 519676 500040 519704
rect 467248 519664 467254 519676
rect 500034 519664 500040 519676
rect 500092 519664 500098 519716
rect 58434 519596 58440 519648
rect 58492 519636 58498 519648
rect 154114 519636 154120 519648
rect 58492 519608 154120 519636
rect 58492 519596 58498 519608
rect 154114 519596 154120 519608
rect 154172 519596 154178 519648
rect 467098 519596 467104 519648
rect 467156 519636 467162 519648
rect 500126 519636 500132 519648
rect 467156 519608 500132 519636
rect 467156 519596 467162 519608
rect 500126 519596 500132 519608
rect 500184 519596 500190 519648
rect 56502 519528 56508 519580
rect 56560 519568 56566 519580
rect 162118 519568 162124 519580
rect 56560 519540 162124 519568
rect 56560 519528 56566 519540
rect 162118 519528 162124 519540
rect 162176 519528 162182 519580
rect 468570 519528 468576 519580
rect 468628 519568 468634 519580
rect 509234 519568 509240 519580
rect 468628 519540 509240 519568
rect 468628 519528 468634 519540
rect 509234 519528 509240 519540
rect 509292 519528 509298 519580
rect 177942 519460 177948 519512
rect 178000 519500 178006 519512
rect 483014 519500 483020 519512
rect 178000 519472 483020 519500
rect 178000 519460 178006 519472
rect 483014 519460 483020 519472
rect 483072 519460 483078 519512
rect 55122 518984 55128 519036
rect 55180 519024 55186 519036
rect 58710 519024 58716 519036
rect 55180 518996 58716 519024
rect 55180 518984 55186 518996
rect 58710 518984 58716 518996
rect 58768 518984 58774 519036
rect 37918 518916 37924 518968
rect 37976 518956 37982 518968
rect 56502 518956 56508 518968
rect 37976 518928 56508 518956
rect 37976 518916 37982 518928
rect 56502 518916 56508 518928
rect 56560 518916 56566 518968
rect 291838 518916 291844 518968
rect 291896 518956 291902 518968
rect 494054 518956 494060 518968
rect 291896 518928 494060 518956
rect 291896 518916 291902 518928
rect 494054 518916 494060 518928
rect 494112 518916 494118 518968
rect 58894 518848 58900 518900
rect 58952 518888 58958 518900
rect 389174 518888 389180 518900
rect 58952 518860 389180 518888
rect 58952 518848 58958 518860
rect 389174 518848 389180 518860
rect 389232 518848 389238 518900
rect 58986 518780 58992 518832
rect 59044 518820 59050 518832
rect 386414 518820 386420 518832
rect 59044 518792 386420 518820
rect 59044 518780 59050 518792
rect 386414 518780 386420 518792
rect 386472 518780 386478 518832
rect 269022 518712 269028 518764
rect 269080 518752 269086 518764
rect 385218 518752 385224 518764
rect 269080 518724 385224 518752
rect 269080 518712 269086 518724
rect 385218 518712 385224 518724
rect 385276 518712 385282 518764
rect 481634 518576 481640 518628
rect 481692 518616 481698 518628
rect 482094 518616 482100 518628
rect 481692 518588 482100 518616
rect 481692 518576 481698 518588
rect 482094 518576 482100 518588
rect 482152 518576 482158 518628
rect 478782 518508 478788 518560
rect 478840 518548 478846 518560
rect 491386 518548 491392 518560
rect 478840 518520 491392 518548
rect 478840 518508 478846 518520
rect 491386 518508 491392 518520
rect 491444 518508 491450 518560
rect 477402 518440 477408 518492
rect 477460 518480 477466 518492
rect 490650 518480 490656 518492
rect 477460 518452 490656 518480
rect 477460 518440 477466 518452
rect 490650 518440 490656 518452
rect 490708 518440 490714 518492
rect 477310 518372 477316 518424
rect 477368 518412 477374 518424
rect 492674 518412 492680 518424
rect 477368 518384 492680 518412
rect 477368 518372 477374 518384
rect 492674 518372 492680 518384
rect 492732 518372 492738 518424
rect 480070 518304 480076 518356
rect 480128 518344 480134 518356
rect 482094 518344 482100 518356
rect 480128 518316 482100 518344
rect 480128 518304 480134 518316
rect 482094 518304 482100 518316
rect 482152 518304 482158 518356
rect 59538 518236 59544 518288
rect 59596 518276 59602 518288
rect 171134 518276 171140 518288
rect 59596 518248 171140 518276
rect 59596 518236 59602 518248
rect 171134 518236 171140 518248
rect 171192 518236 171198 518288
rect 476758 518236 476764 518288
rect 476816 518276 476822 518288
rect 493410 518276 493416 518288
rect 476816 518248 493416 518276
rect 476816 518236 476822 518248
rect 493410 518236 493416 518248
rect 493468 518236 493474 518288
rect 56778 518168 56784 518220
rect 56836 518208 56842 518220
rect 62022 518208 62028 518220
rect 56836 518180 62028 518208
rect 56836 518168 56842 518180
rect 62022 518168 62028 518180
rect 62080 518168 62086 518220
rect 374638 518208 374644 518220
rect 64846 518180 374644 518208
rect 60918 518100 60924 518152
rect 60976 518140 60982 518152
rect 61930 518140 61936 518152
rect 60976 518112 61936 518140
rect 60976 518100 60982 518112
rect 61930 518100 61936 518112
rect 61988 518100 61994 518152
rect 64846 518072 64874 518180
rect 374638 518168 374644 518180
rect 374696 518168 374702 518220
rect 474090 518168 474096 518220
rect 474148 518208 474154 518220
rect 491846 518208 491852 518220
rect 474148 518180 491852 518208
rect 474148 518168 474154 518180
rect 491846 518168 491852 518180
rect 491904 518168 491910 518220
rect 476114 518100 476120 518152
rect 476172 518140 476178 518152
rect 494790 518140 494796 518152
rect 476172 518112 494796 518140
rect 476172 518100 476178 518112
rect 494790 518100 494796 518112
rect 494848 518100 494854 518152
rect 59004 518044 64874 518072
rect 59004 517880 59032 518044
rect 478782 518032 478788 518084
rect 478840 518072 478846 518084
rect 483106 518072 483112 518084
rect 478840 518044 483112 518072
rect 478840 518032 478846 518044
rect 483106 518032 483112 518044
rect 483164 518032 483170 518084
rect 478966 517964 478972 518016
rect 479024 518004 479030 518016
rect 480070 518004 480076 518016
rect 479024 517976 480076 518004
rect 479024 517964 479030 517976
rect 480070 517964 480076 517976
rect 480128 517964 480134 518016
rect 58986 517828 58992 517880
rect 59044 517828 59050 517880
rect 60918 517664 60924 517676
rect 57440 517636 60924 517664
rect 57440 517064 57468 517636
rect 60918 517624 60924 517636
rect 60976 517624 60982 517676
rect 57698 517556 57704 517608
rect 57756 517596 57762 517608
rect 60826 517596 60832 517608
rect 57756 517568 60832 517596
rect 57756 517556 57762 517568
rect 60826 517556 60832 517568
rect 60884 517556 60890 517608
rect 60366 517488 60372 517540
rect 60424 517528 60430 517540
rect 60734 517528 60740 517540
rect 60424 517500 60740 517528
rect 60424 517488 60430 517500
rect 60734 517488 60740 517500
rect 60792 517488 60798 517540
rect 57422 517012 57428 517064
rect 57480 517012 57486 517064
rect 56502 516128 56508 516180
rect 56560 516168 56566 516180
rect 57238 516168 57244 516180
rect 56560 516140 57244 516168
rect 56560 516128 56566 516140
rect 57238 516128 57244 516140
rect 57296 516128 57302 516180
rect 56962 511980 56968 512032
rect 57020 512020 57026 512032
rect 58434 512020 58440 512032
rect 57020 511992 58440 512020
rect 57020 511980 57026 511992
rect 58434 511980 58440 511992
rect 58492 511980 58498 512032
rect 481634 510552 481640 510604
rect 481692 510592 481698 510604
rect 483106 510592 483112 510604
rect 481692 510564 483112 510592
rect 481692 510552 481698 510564
rect 483106 510552 483112 510564
rect 483164 510552 483170 510604
rect 482094 510484 482100 510536
rect 482152 510524 482158 510536
rect 482554 510524 482560 510536
rect 482152 510496 482560 510524
rect 482152 510484 482158 510496
rect 482554 510484 482560 510496
rect 482612 510484 482618 510536
rect 482830 506404 482836 506456
rect 482888 506444 482894 506456
rect 491386 506444 491392 506456
rect 482888 506416 491392 506444
rect 482888 506404 482894 506416
rect 491386 506404 491392 506416
rect 491444 506404 491450 506456
rect 482922 506336 482928 506388
rect 482980 506376 482986 506388
rect 490650 506376 490656 506388
rect 482980 506348 490656 506376
rect 482980 506336 482986 506348
rect 490650 506336 490656 506348
rect 490708 506336 490714 506388
rect 57698 500896 57704 500948
rect 57756 500936 57762 500948
rect 58802 500936 58808 500948
rect 57756 500908 58808 500936
rect 57756 500896 57762 500908
rect 58802 500896 58808 500908
rect 58860 500896 58866 500948
rect 482830 500896 482836 500948
rect 482888 500936 482894 500948
rect 494054 500936 494060 500948
rect 482888 500908 494060 500936
rect 482888 500896 482894 500908
rect 494054 500896 494060 500908
rect 494112 500896 494118 500948
rect 482922 500828 482928 500880
rect 482980 500868 482986 500880
rect 492674 500868 492680 500880
rect 482980 500840 492680 500868
rect 482980 500828 482986 500840
rect 492674 500828 492680 500840
rect 492732 500828 492738 500880
rect 56870 499672 56876 499724
rect 56928 499712 56934 499724
rect 57146 499712 57152 499724
rect 56928 499684 57152 499712
rect 56928 499672 56934 499684
rect 57146 499672 57152 499684
rect 57204 499672 57210 499724
rect 57054 490560 57060 490612
rect 57112 490600 57118 490612
rect 57330 490600 57336 490612
rect 57112 490572 57336 490600
rect 57112 490560 57118 490572
rect 57330 490560 57336 490572
rect 57388 490560 57394 490612
rect 482094 480156 482100 480208
rect 482152 480196 482158 480208
rect 494790 480196 494796 480208
rect 482152 480168 494796 480196
rect 482152 480156 482158 480168
rect 494790 480156 494796 480168
rect 494848 480156 494854 480208
rect 482094 478796 482100 478848
rect 482152 478836 482158 478848
rect 497550 478836 497556 478848
rect 482152 478808 497556 478836
rect 482152 478796 482158 478808
rect 497550 478796 497556 478808
rect 497608 478796 497614 478848
rect 479242 477980 479248 478032
rect 479300 478020 479306 478032
rect 479518 478020 479524 478032
rect 479300 477992 479524 478020
rect 479300 477980 479306 477992
rect 479518 477980 479524 477992
rect 479576 477980 479582 478032
rect 3418 476008 3424 476060
rect 3476 476048 3482 476060
rect 37918 476048 37924 476060
rect 3476 476020 37924 476048
rect 3476 476008 3482 476020
rect 37918 476008 37924 476020
rect 37976 476008 37982 476060
rect 482094 474648 482100 474700
rect 482152 474688 482158 474700
rect 485866 474688 485872 474700
rect 482152 474660 485872 474688
rect 482152 474648 482158 474660
rect 485866 474648 485872 474660
rect 485924 474648 485930 474700
rect 482094 473288 482100 473340
rect 482152 473328 482158 473340
rect 488810 473328 488816 473340
rect 482152 473300 488816 473328
rect 482152 473288 482158 473300
rect 488810 473288 488816 473300
rect 488868 473288 488874 473340
rect 482094 471928 482100 471980
rect 482152 471968 482158 471980
rect 498654 471968 498660 471980
rect 482152 471940 498660 471968
rect 482152 471928 482158 471940
rect 498654 471928 498660 471940
rect 498712 471928 498718 471980
rect 482002 471860 482008 471912
rect 482060 471900 482066 471912
rect 487430 471900 487436 471912
rect 482060 471872 487436 471900
rect 482060 471860 482066 471872
rect 487430 471860 487436 471872
rect 487488 471860 487494 471912
rect 482094 470500 482100 470552
rect 482152 470540 482158 470552
rect 500126 470540 500132 470552
rect 482152 470512 500132 470540
rect 482152 470500 482158 470512
rect 500126 470500 500132 470512
rect 500184 470500 500190 470552
rect 482002 470432 482008 470484
rect 482060 470472 482066 470484
rect 486694 470472 486700 470484
rect 482060 470444 486700 470472
rect 482060 470432 482066 470444
rect 486694 470432 486700 470444
rect 486752 470432 486758 470484
rect 482094 469140 482100 469192
rect 482152 469180 482158 469192
rect 500034 469180 500040 469192
rect 482152 469152 500040 469180
rect 482152 469140 482158 469152
rect 500034 469140 500040 469152
rect 500092 469140 500098 469192
rect 482002 469072 482008 469124
rect 482060 469112 482066 469124
rect 494698 469112 494704 469124
rect 482060 469084 494704 469112
rect 482060 469072 482066 469084
rect 494698 469072 494704 469084
rect 494756 469072 494762 469124
rect 482094 467780 482100 467832
rect 482152 467820 482158 467832
rect 487246 467820 487252 467832
rect 482152 467792 487252 467820
rect 482152 467780 482158 467792
rect 487246 467780 487252 467792
rect 487304 467780 487310 467832
rect 482002 467712 482008 467764
rect 482060 467752 482066 467764
rect 487338 467752 487344 467764
rect 482060 467724 487344 467752
rect 482060 467712 482066 467724
rect 487338 467712 487344 467724
rect 487396 467712 487402 467764
rect 482002 464992 482008 465044
rect 482060 465032 482066 465044
rect 505370 465032 505376 465044
rect 482060 465004 505376 465032
rect 482060 464992 482066 465004
rect 505370 464992 505376 465004
rect 505428 464992 505434 465044
rect 482094 464924 482100 464976
rect 482152 464964 482158 464976
rect 504266 464964 504272 464976
rect 482152 464936 504272 464964
rect 482152 464924 482158 464936
rect 504266 464924 504272 464936
rect 504324 464924 504330 464976
rect 482094 464788 482100 464840
rect 482152 464828 482158 464840
rect 489362 464828 489368 464840
rect 482152 464800 489368 464828
rect 482152 464788 482158 464800
rect 489362 464788 489368 464800
rect 489420 464788 489426 464840
rect 482094 463632 482100 463684
rect 482152 463672 482158 463684
rect 490190 463672 490196 463684
rect 482152 463644 490196 463672
rect 482152 463632 482158 463644
rect 490190 463632 490196 463644
rect 490248 463632 490254 463684
rect 482094 463292 482100 463344
rect 482152 463332 482158 463344
rect 488074 463332 488080 463344
rect 482152 463304 488080 463332
rect 482152 463292 482158 463304
rect 488074 463292 488080 463304
rect 488132 463292 488138 463344
rect 482002 462272 482008 462324
rect 482060 462312 482066 462324
rect 505278 462312 505284 462324
rect 482060 462284 505284 462312
rect 482060 462272 482066 462284
rect 505278 462272 505284 462284
rect 505336 462272 505342 462324
rect 481910 462204 481916 462256
rect 481968 462244 481974 462256
rect 502610 462244 502616 462256
rect 481968 462216 502616 462244
rect 481968 462204 481974 462216
rect 502610 462204 502616 462216
rect 502668 462204 502674 462256
rect 482094 462136 482100 462188
rect 482152 462176 482158 462188
rect 490098 462176 490104 462188
rect 482152 462148 490104 462176
rect 482152 462136 482158 462148
rect 490098 462136 490104 462148
rect 490156 462136 490162 462188
rect 482094 460776 482100 460828
rect 482152 460816 482158 460828
rect 488626 460816 488632 460828
rect 482152 460788 488632 460816
rect 482152 460776 482158 460788
rect 488626 460776 488632 460788
rect 488684 460776 488690 460828
rect 482002 459484 482008 459536
rect 482060 459524 482066 459536
rect 504174 459524 504180 459536
rect 482060 459496 504180 459524
rect 482060 459484 482066 459496
rect 504174 459484 504180 459496
rect 504232 459484 504238 459536
rect 482094 459416 482100 459468
rect 482152 459456 482158 459468
rect 495894 459456 495900 459468
rect 482152 459428 495900 459456
rect 482152 459416 482158 459428
rect 495894 459416 495900 459428
rect 495952 459416 495958 459468
rect 482002 458124 482008 458176
rect 482060 458164 482066 458176
rect 491846 458164 491852 458176
rect 482060 458136 491852 458164
rect 482060 458124 482066 458136
rect 491846 458124 491852 458136
rect 491904 458124 491910 458176
rect 482094 458056 482100 458108
rect 482152 458096 482158 458108
rect 490006 458096 490012 458108
rect 482152 458068 490012 458096
rect 482152 458056 482158 458068
rect 490006 458056 490012 458068
rect 490064 458056 490070 458108
rect 482094 456696 482100 456748
rect 482152 456736 482158 456748
rect 509418 456736 509424 456748
rect 482152 456708 509424 456736
rect 482152 456696 482158 456708
rect 509418 456696 509424 456708
rect 509476 456696 509482 456748
rect 482002 455336 482008 455388
rect 482060 455376 482066 455388
rect 493410 455376 493416 455388
rect 482060 455348 493416 455376
rect 482060 455336 482066 455348
rect 493410 455336 493416 455348
rect 493468 455336 493474 455388
rect 482094 455268 482100 455320
rect 482152 455308 482158 455320
rect 489914 455308 489920 455320
rect 482152 455280 489920 455308
rect 482152 455268 482158 455280
rect 489914 455268 489920 455280
rect 489972 455268 489978 455320
rect 482094 453976 482100 454028
rect 482152 454016 482158 454028
rect 491662 454016 491668 454028
rect 482152 453988 491668 454016
rect 482152 453976 482158 453988
rect 491662 453976 491668 453988
rect 491720 453976 491726 454028
rect 482094 452548 482100 452600
rect 482152 452588 482158 452600
rect 497458 452588 497464 452600
rect 482152 452560 497464 452588
rect 482152 452548 482158 452560
rect 497458 452548 497464 452560
rect 497516 452548 497522 452600
rect 482094 452412 482100 452464
rect 482152 452452 482158 452464
rect 489270 452452 489276 452464
rect 482152 452424 489276 452452
rect 482152 452412 482158 452424
rect 489270 452412 489276 452424
rect 489328 452412 489334 452464
rect 482186 449828 482192 449880
rect 482244 449868 482250 449880
rect 509326 449868 509332 449880
rect 482244 449840 509332 449868
rect 482244 449828 482250 449840
rect 509326 449828 509332 449840
rect 509384 449828 509390 449880
rect 482094 449760 482100 449812
rect 482152 449800 482158 449812
rect 494514 449800 494520 449812
rect 482152 449772 494520 449800
rect 482152 449760 482158 449772
rect 494514 449760 494520 449772
rect 494572 449760 494578 449812
rect 482186 449692 482192 449744
rect 482244 449732 482250 449744
rect 493226 449732 493232 449744
rect 482244 449704 493232 449732
rect 482244 449692 482250 449704
rect 493226 449692 493232 449704
rect 493284 449692 493290 449744
rect 482186 448468 482192 448520
rect 482244 448508 482250 448520
rect 494422 448508 494428 448520
rect 482244 448480 494428 448508
rect 482244 448468 482250 448480
rect 494422 448468 494428 448480
rect 494480 448468 494486 448520
rect 482094 448400 482100 448452
rect 482152 448440 482158 448452
rect 490558 448440 490564 448452
rect 482152 448412 490564 448440
rect 482152 448400 482158 448412
rect 490558 448400 490564 448412
rect 490616 448400 490622 448452
rect 482002 447040 482008 447092
rect 482060 447080 482066 447092
rect 508130 447080 508136 447092
rect 482060 447052 508136 447080
rect 482060 447040 482066 447052
rect 508130 447040 508136 447052
rect 508188 447040 508194 447092
rect 482094 446972 482100 447024
rect 482152 447012 482158 447024
rect 493042 447012 493048 447024
rect 482152 446984 493048 447012
rect 482152 446972 482158 446984
rect 493042 446972 493048 446984
rect 493100 446972 493106 447024
rect 482186 446904 482192 446956
rect 482244 446944 482250 446956
rect 491754 446944 491760 446956
rect 482244 446916 491760 446944
rect 482244 446904 482250 446916
rect 491754 446904 491760 446916
rect 491812 446904 491818 446956
rect 482094 445680 482100 445732
rect 482152 445720 482158 445732
rect 493318 445720 493324 445732
rect 482152 445692 493324 445720
rect 482152 445680 482158 445692
rect 493318 445680 493324 445692
rect 493376 445680 493382 445732
rect 482186 445612 482192 445664
rect 482244 445652 482250 445664
rect 493134 445652 493140 445664
rect 482244 445624 493140 445652
rect 482244 445612 482250 445624
rect 493134 445612 493140 445624
rect 493192 445612 493198 445664
rect 482186 444320 482192 444372
rect 482244 444360 482250 444372
rect 492766 444360 492772 444372
rect 482244 444332 492772 444360
rect 482244 444320 482250 444332
rect 492766 444320 492772 444332
rect 492824 444320 492830 444372
rect 482094 444252 482100 444304
rect 482152 444292 482158 444304
rect 492858 444292 492864 444304
rect 482152 444264 492864 444292
rect 482152 444252 482158 444264
rect 492858 444252 492864 444264
rect 492916 444252 492922 444304
rect 482186 442892 482192 442944
rect 482244 442932 482250 442944
rect 506842 442932 506848 442944
rect 482244 442904 506848 442932
rect 482244 442892 482250 442904
rect 506842 442892 506848 442904
rect 506900 442892 506906 442944
rect 482094 441532 482100 441584
rect 482152 441572 482158 441584
rect 508222 441572 508228 441584
rect 482152 441544 508228 441572
rect 482152 441532 482158 441544
rect 508222 441532 508228 441544
rect 508280 441532 508286 441584
rect 482186 441464 482192 441516
rect 482244 441504 482250 441516
rect 492950 441504 492956 441516
rect 482244 441476 492956 441504
rect 482244 441464 482250 441476
rect 492950 441464 492956 441476
rect 493008 441464 493014 441516
rect 482186 440172 482192 440224
rect 482244 440212 482250 440224
rect 505186 440212 505192 440224
rect 482244 440184 505192 440212
rect 482244 440172 482250 440184
rect 505186 440172 505192 440184
rect 505244 440172 505250 440224
rect 482094 438812 482100 438864
rect 482152 438852 482158 438864
rect 506750 438852 506756 438864
rect 482152 438824 506756 438852
rect 482152 438812 482158 438824
rect 506750 438812 506756 438824
rect 506808 438812 506814 438864
rect 482186 438744 482192 438796
rect 482244 438784 482250 438796
rect 502518 438784 502524 438796
rect 482244 438756 502524 438784
rect 482244 438744 482250 438756
rect 502518 438744 502524 438756
rect 502576 438744 502582 438796
rect 482186 428204 482192 428256
rect 482244 428244 482250 428256
rect 482830 428244 482836 428256
rect 482244 428216 482836 428244
rect 482244 428204 482250 428216
rect 482830 428204 482836 428216
rect 482888 428204 482894 428256
rect 482830 425008 482836 425060
rect 482888 425048 482894 425060
rect 491294 425048 491300 425060
rect 482888 425020 491300 425048
rect 482888 425008 482894 425020
rect 491294 425008 491300 425020
rect 491352 425008 491358 425060
rect 482830 423580 482836 423632
rect 482888 423620 482894 423632
rect 491478 423620 491484 423632
rect 482888 423592 491484 423620
rect 482888 423580 482894 423592
rect 491478 423580 491484 423592
rect 491536 423580 491542 423632
rect 482830 423308 482836 423360
rect 482888 423348 482894 423360
rect 486142 423348 486148 423360
rect 482888 423320 486148 423348
rect 482888 423308 482894 423320
rect 486142 423308 486148 423320
rect 486200 423308 486206 423360
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 26878 422328 26884 422340
rect 3476 422300 26884 422328
rect 3476 422288 3482 422300
rect 26878 422288 26884 422300
rect 26936 422288 26942 422340
rect 482830 418072 482836 418124
rect 482888 418112 482894 418124
rect 494238 418112 494244 418124
rect 482888 418084 494244 418112
rect 482888 418072 482894 418084
rect 494238 418072 494244 418084
rect 494296 418072 494302 418124
rect 482186 418004 482192 418056
rect 482244 418044 482250 418056
rect 494330 418044 494336 418056
rect 482244 418016 494336 418044
rect 482244 418004 482250 418016
rect 494330 418004 494336 418016
rect 494388 418004 494394 418056
rect 482830 416712 482836 416764
rect 482888 416752 482894 416764
rect 499850 416752 499856 416764
rect 482888 416724 499856 416752
rect 482888 416712 482894 416724
rect 499850 416712 499856 416724
rect 499908 416712 499914 416764
rect 482830 415352 482836 415404
rect 482888 415392 482894 415404
rect 497182 415392 497188 415404
rect 482888 415364 497188 415392
rect 482888 415352 482894 415364
rect 497182 415352 497188 415364
rect 497240 415352 497246 415404
rect 482186 415284 482192 415336
rect 482244 415324 482250 415336
rect 497274 415324 497280 415336
rect 482244 415296 497280 415324
rect 482244 415284 482250 415296
rect 497274 415284 497280 415296
rect 497332 415284 497338 415336
rect 482186 413924 482192 413976
rect 482244 413964 482250 413976
rect 498470 413964 498476 413976
rect 482244 413936 498476 413964
rect 482244 413924 482250 413936
rect 498470 413924 498476 413936
rect 498528 413924 498534 413976
rect 482830 413856 482836 413908
rect 482888 413896 482894 413908
rect 497090 413896 497096 413908
rect 482888 413868 497096 413896
rect 482888 413856 482894 413868
rect 497090 413856 497096 413868
rect 497148 413856 497154 413908
rect 482830 412496 482836 412548
rect 482888 412536 482894 412548
rect 487982 412536 487988 412548
rect 482888 412508 487988 412536
rect 482888 412496 482894 412508
rect 487982 412496 487988 412508
rect 488040 412496 488046 412548
rect 482830 411204 482836 411256
rect 482888 411244 482894 411256
rect 503990 411244 503996 411256
rect 482888 411216 503996 411244
rect 482888 411204 482894 411216
rect 503990 411204 503996 411216
rect 504048 411204 504054 411256
rect 482186 411136 482192 411188
rect 482244 411176 482250 411188
rect 486050 411176 486056 411188
rect 482244 411148 486056 411176
rect 482244 411136 482250 411148
rect 486050 411136 486056 411148
rect 486108 411136 486114 411188
rect 482186 410932 482192 410984
rect 482244 410972 482250 410984
rect 487798 410972 487804 410984
rect 482244 410944 487804 410972
rect 482244 410932 482250 410944
rect 487798 410932 487804 410944
rect 487856 410932 487862 410984
rect 482830 409776 482836 409828
rect 482888 409816 482894 409828
rect 487890 409816 487896 409828
rect 482888 409788 487896 409816
rect 482888 409776 482894 409788
rect 487890 409776 487896 409788
rect 487948 409776 487954 409828
rect 482830 408416 482836 408468
rect 482888 408456 482894 408468
rect 502334 408456 502340 408468
rect 482888 408428 502340 408456
rect 482888 408416 482894 408428
rect 502334 408416 502340 408428
rect 502392 408416 502398 408468
rect 482186 408348 482192 408400
rect 482244 408388 482250 408400
rect 487614 408388 487620 408400
rect 482244 408360 487620 408388
rect 482244 408348 482250 408360
rect 487614 408348 487620 408360
rect 487672 408348 487678 408400
rect 482830 407056 482836 407108
rect 482888 407096 482894 407108
rect 499666 407096 499672 407108
rect 482888 407068 499672 407096
rect 482888 407056 482894 407068
rect 499666 407056 499672 407068
rect 499724 407056 499730 407108
rect 482186 406988 482192 407040
rect 482244 407028 482250 407040
rect 496998 407028 497004 407040
rect 482244 407000 497004 407028
rect 482244 406988 482250 407000
rect 496998 406988 497004 407000
rect 497056 406988 497062 407040
rect 482830 405628 482836 405680
rect 482888 405668 482894 405680
rect 494146 405668 494152 405680
rect 482888 405640 494152 405668
rect 482888 405628 482894 405640
rect 494146 405628 494152 405640
rect 494204 405628 494210 405680
rect 482830 402908 482836 402960
rect 482888 402948 482894 402960
rect 501138 402948 501144 402960
rect 482888 402920 501144 402948
rect 482888 402908 482894 402920
rect 501138 402908 501144 402920
rect 501196 402908 501202 402960
rect 482830 401548 482836 401600
rect 482888 401588 482894 401600
rect 502426 401588 502432 401600
rect 482888 401560 502432 401588
rect 482888 401548 482894 401560
rect 502426 401548 502432 401560
rect 502484 401548 502490 401600
rect 482830 401276 482836 401328
rect 482888 401316 482894 401328
rect 489086 401316 489092 401328
rect 482888 401288 489092 401316
rect 482888 401276 482894 401288
rect 489086 401276 489092 401288
rect 489144 401276 489150 401328
rect 482186 400120 482192 400172
rect 482244 400160 482250 400172
rect 496906 400160 496912 400172
rect 482244 400132 496912 400160
rect 482244 400120 482250 400132
rect 496906 400120 496912 400132
rect 496964 400120 496970 400172
rect 482830 400052 482836 400104
rect 482888 400092 482894 400104
rect 495434 400092 495440 400104
rect 482888 400064 495440 400092
rect 482888 400052 482894 400064
rect 495434 400052 495440 400064
rect 495492 400052 495498 400104
rect 482002 398760 482008 398812
rect 482060 398800 482066 398812
rect 500954 398800 500960 398812
rect 482060 398772 500960 398800
rect 482060 398760 482066 398772
rect 500954 398760 500960 398772
rect 501012 398760 501018 398812
rect 482830 398692 482836 398744
rect 482888 398732 482894 398744
rect 498286 398732 498292 398744
rect 482888 398704 498292 398732
rect 482888 398692 482894 398704
rect 498286 398692 498292 398704
rect 498344 398692 498350 398744
rect 482186 398624 482192 398676
rect 482244 398664 482250 398676
rect 493502 398664 493508 398676
rect 482244 398636 493508 398664
rect 482244 398624 482250 398636
rect 493502 398624 493508 398636
rect 493560 398624 493566 398676
rect 482830 397400 482836 397452
rect 482888 397440 482894 397452
rect 503898 397440 503904 397452
rect 482888 397412 503904 397440
rect 482888 397400 482894 397412
rect 503898 397400 503904 397412
rect 503956 397400 503962 397452
rect 482186 397332 482192 397384
rect 482244 397372 482250 397384
rect 495526 397372 495532 397384
rect 482244 397344 495532 397372
rect 482244 397332 482250 397344
rect 495526 397332 495532 397344
rect 495584 397332 495590 397384
rect 482186 395972 482192 396024
rect 482244 396012 482250 396024
rect 514846 396012 514852 396024
rect 482244 395984 514852 396012
rect 482244 395972 482250 395984
rect 514846 395972 514852 395984
rect 514904 395972 514910 396024
rect 482830 395904 482836 395956
rect 482888 395944 482894 395956
rect 501046 395944 501052 395956
rect 482888 395916 501052 395944
rect 482888 395904 482894 395916
rect 501046 395904 501052 395916
rect 501104 395904 501110 395956
rect 482186 394612 482192 394664
rect 482244 394652 482250 394664
rect 514754 394652 514760 394664
rect 482244 394624 514760 394652
rect 482244 394612 482250 394624
rect 514754 394612 514760 394624
rect 514812 394612 514818 394664
rect 482830 394544 482836 394596
rect 482888 394584 482894 394596
rect 512086 394584 512092 394596
rect 482888 394556 512092 394584
rect 482888 394544 482894 394556
rect 512086 394544 512092 394556
rect 512144 394544 512150 394596
rect 482186 393252 482192 393304
rect 482244 393292 482250 393304
rect 482646 393292 482652 393304
rect 482244 393264 482652 393292
rect 482244 393252 482250 393264
rect 482646 393252 482652 393264
rect 482704 393252 482710 393304
rect 482830 393252 482836 393304
rect 482888 393292 482894 393304
rect 513374 393292 513380 393304
rect 482888 393264 513380 393292
rect 482888 393252 482894 393264
rect 513374 393252 513380 393264
rect 513432 393252 513438 393304
rect 482094 393184 482100 393236
rect 482152 393224 482158 393236
rect 509234 393224 509240 393236
rect 482152 393196 509240 393224
rect 482152 393184 482158 393196
rect 509234 393184 509240 393196
rect 509292 393184 509298 393236
rect 482922 393116 482928 393168
rect 482980 393156 482986 393168
rect 506658 393156 506664 393168
rect 482980 393128 506664 393156
rect 482980 393116 482986 393128
rect 506658 393116 506664 393128
rect 506716 393116 506722 393168
rect 482830 391892 482836 391944
rect 482888 391932 482894 391944
rect 511994 391932 512000 391944
rect 482888 391904 512000 391932
rect 482888 391892 482894 391904
rect 511994 391892 512000 391904
rect 512052 391892 512058 391944
rect 482922 391824 482928 391876
rect 482980 391864 482986 391876
rect 512178 391864 512184 391876
rect 482980 391836 512184 391864
rect 482980 391824 482986 391836
rect 512178 391824 512184 391836
rect 512236 391824 512242 391876
rect 482922 390464 482928 390516
rect 482980 390504 482986 390516
rect 510614 390504 510620 390516
rect 482980 390476 510620 390504
rect 482980 390464 482986 390476
rect 510614 390464 510620 390476
rect 510672 390464 510678 390516
rect 58802 389852 58808 389904
rect 58860 389892 58866 389904
rect 122098 389892 122104 389904
rect 58860 389864 122104 389892
rect 58860 389852 58866 389864
rect 122098 389852 122104 389864
rect 122156 389852 122162 389904
rect 60366 389784 60372 389836
rect 60424 389824 60430 389836
rect 265618 389824 265624 389836
rect 60424 389796 265624 389824
rect 60424 389784 60430 389796
rect 265618 389784 265624 389796
rect 265676 389784 265682 389836
rect 474642 389104 474648 389156
rect 474700 389144 474706 389156
rect 546494 389144 546500 389156
rect 474700 389116 546500 389144
rect 474700 389104 474706 389116
rect 546494 389104 546500 389116
rect 546552 389104 546558 389156
rect 26878 388424 26884 388476
rect 26936 388464 26942 388476
rect 95694 388464 95700 388476
rect 26936 388436 95700 388464
rect 26936 388424 26942 388436
rect 95694 388424 95700 388436
rect 95752 388424 95758 388476
rect 118694 387744 118700 387796
rect 118752 387784 118758 387796
rect 534718 387784 534724 387796
rect 118752 387756 534724 387784
rect 118752 387744 118758 387756
rect 534718 387744 534724 387756
rect 534776 387744 534782 387796
rect 57238 387676 57244 387728
rect 57296 387716 57302 387728
rect 150434 387716 150440 387728
rect 57296 387688 150440 387716
rect 57296 387676 57302 387688
rect 150434 387676 150440 387688
rect 150492 387676 150498 387728
rect 272518 387676 272524 387728
rect 272576 387716 272582 387728
rect 506474 387716 506480 387728
rect 272576 387688 506480 387716
rect 272576 387676 272582 387688
rect 506474 387676 506480 387688
rect 506532 387676 506538 387728
rect 58710 387608 58716 387660
rect 58768 387648 58774 387660
rect 143534 387648 143540 387660
rect 58768 387620 143540 387648
rect 58768 387608 58774 387620
rect 143534 387608 143540 387620
rect 143592 387648 143598 387660
rect 144362 387648 144368 387660
rect 143592 387620 144368 387648
rect 143592 387608 143598 387620
rect 144362 387608 144368 387620
rect 144420 387608 144426 387660
rect 274634 387608 274640 387660
rect 274692 387648 274698 387660
rect 505094 387648 505100 387660
rect 274692 387620 505100 387648
rect 274692 387608 274698 387620
rect 505094 387608 505100 387620
rect 505152 387608 505158 387660
rect 56134 387540 56140 387592
rect 56192 387580 56198 387592
rect 132494 387580 132500 387592
rect 56192 387552 132500 387580
rect 56192 387540 56198 387552
rect 132494 387540 132500 387552
rect 132552 387580 132558 387592
rect 137186 387580 137192 387592
rect 132552 387552 137192 387580
rect 132552 387540 132558 387552
rect 137186 387540 137192 387552
rect 137244 387540 137250 387592
rect 270402 387540 270408 387592
rect 270460 387580 270466 387592
rect 482646 387580 482652 387592
rect 270460 387552 482652 387580
rect 270460 387540 270466 387552
rect 482646 387540 482652 387552
rect 482704 387540 482710 387592
rect 498194 387540 498200 387592
rect 498252 387580 498258 387592
rect 498838 387580 498844 387592
rect 498252 387552 498844 387580
rect 498252 387540 498258 387552
rect 498838 387540 498844 387552
rect 498896 387540 498902 387592
rect 60550 387472 60556 387524
rect 60608 387512 60614 387524
rect 124122 387512 124128 387524
rect 60608 387484 124128 387512
rect 60608 387472 60614 387484
rect 124122 387472 124128 387484
rect 124180 387472 124186 387524
rect 106182 387336 106188 387388
rect 106240 387376 106246 387388
rect 147674 387376 147680 387388
rect 106240 387348 147680 387376
rect 106240 387336 106246 387348
rect 147674 387336 147680 387348
rect 147732 387336 147738 387388
rect 108298 387268 108304 387320
rect 108356 387308 108362 387320
rect 162302 387308 162308 387320
rect 108356 387280 162308 387308
rect 108356 387268 108362 387280
rect 162302 387268 162308 387280
rect 162360 387308 162366 387320
rect 162762 387308 162768 387320
rect 162360 387280 162768 387308
rect 162360 387268 162366 387280
rect 162762 387268 162768 387280
rect 162820 387268 162826 387320
rect 60274 387200 60280 387252
rect 60332 387240 60338 387252
rect 140774 387240 140780 387252
rect 60332 387212 140780 387240
rect 60332 387200 60338 387212
rect 140774 387200 140780 387212
rect 140832 387200 140838 387252
rect 62114 387132 62120 387184
rect 62172 387172 62178 387184
rect 154574 387172 154580 387184
rect 62172 387144 154580 387172
rect 62172 387132 62178 387144
rect 154574 387132 154580 387144
rect 154632 387172 154638 387184
rect 155126 387172 155132 387184
rect 154632 387144 155132 387172
rect 154632 387132 154638 387144
rect 155126 387132 155132 387144
rect 155184 387132 155190 387184
rect 277210 387132 277216 387184
rect 277268 387172 277274 387184
rect 445754 387172 445760 387184
rect 277268 387144 445760 387172
rect 277268 387132 277274 387144
rect 445754 387132 445760 387144
rect 445812 387132 445818 387184
rect 115842 387064 115848 387116
rect 115900 387104 115906 387116
rect 498194 387104 498200 387116
rect 115900 387076 498200 387104
rect 115900 387064 115906 387076
rect 498194 387064 498200 387076
rect 498252 387064 498258 387116
rect 458818 386860 458824 386912
rect 458876 386900 458882 386912
rect 460106 386900 460112 386912
rect 458876 386872 460112 386900
rect 458876 386860 458882 386872
rect 460106 386860 460112 386872
rect 460164 386860 460170 386912
rect 138658 386452 138664 386504
rect 138716 386492 138722 386504
rect 191006 386492 191012 386504
rect 138716 386464 191012 386492
rect 138716 386452 138722 386464
rect 191006 386452 191012 386464
rect 191064 386492 191070 386504
rect 191742 386492 191748 386504
rect 191064 386464 191748 386492
rect 191064 386452 191070 386464
rect 191742 386452 191748 386464
rect 191800 386452 191806 386504
rect 105538 386384 105544 386436
rect 105596 386424 105602 386436
rect 177298 386424 177304 386436
rect 105596 386396 177304 386424
rect 105596 386384 105602 386396
rect 177298 386384 177304 386396
rect 177356 386384 177362 386436
rect 471974 386316 471980 386368
rect 472032 386356 472038 386368
rect 479610 386356 479616 386368
rect 472032 386328 479616 386356
rect 472032 386316 472038 386328
rect 479610 386316 479616 386328
rect 479668 386316 479674 386368
rect 162762 384956 162768 385008
rect 162820 384996 162826 385008
rect 543826 384996 543832 385008
rect 162820 384968 543832 384996
rect 162820 384956 162826 384968
rect 543826 384956 543832 384968
rect 543884 384956 543890 385008
rect 191742 384888 191748 384940
rect 191800 384928 191806 384940
rect 547966 384928 547972 384940
rect 191800 384900 547972 384928
rect 191800 384888 191806 384900
rect 547966 384888 547972 384900
rect 548024 384888 548030 384940
rect 132494 384452 132500 384464
rect 122806 384424 132500 384452
rect 84102 384276 84108 384328
rect 84160 384316 84166 384328
rect 122806 384316 122834 384424
rect 132494 384412 132500 384424
rect 132552 384412 132558 384464
rect 84160 384288 122834 384316
rect 84160 384276 84166 384288
rect 177298 383596 177304 383648
rect 177356 383636 177362 383648
rect 547874 383636 547880 383648
rect 177356 383608 547880 383636
rect 177356 383596 177362 383608
rect 547874 383596 547880 383608
rect 547932 383596 547938 383648
rect 122098 382916 122104 382968
rect 122156 382956 122162 382968
rect 127618 382956 127624 382968
rect 122156 382928 127624 382956
rect 122156 382916 122162 382928
rect 127618 382916 127624 382928
rect 127676 382916 127682 382968
rect 449894 382916 449900 382968
rect 449952 382956 449958 382968
rect 471974 382956 471980 382968
rect 449952 382928 471980 382956
rect 449952 382916 449958 382928
rect 471974 382916 471980 382928
rect 472032 382916 472038 382968
rect 282822 380808 282828 380860
rect 282880 380848 282886 380860
rect 539962 380848 539968 380860
rect 282880 380820 539968 380848
rect 282880 380808 282886 380820
rect 539962 380808 539968 380820
rect 540020 380808 540026 380860
rect 127618 378088 127624 378140
rect 127676 378128 127682 378140
rect 133138 378128 133144 378140
rect 127676 378100 133144 378128
rect 127676 378088 127682 378100
rect 133138 378088 133144 378100
rect 133196 378088 133202 378140
rect 260742 378088 260748 378140
rect 260800 378128 260806 378140
rect 529382 378128 529388 378140
rect 260800 378100 529388 378128
rect 260800 378088 260806 378100
rect 529382 378088 529388 378100
rect 529440 378088 529446 378140
rect 282822 378020 282828 378072
rect 282880 378060 282886 378072
rect 539870 378060 539876 378072
rect 282880 378032 539876 378060
rect 282880 378020 282886 378032
rect 539870 378020 539876 378032
rect 539928 378020 539934 378072
rect 265618 377408 265624 377460
rect 265676 377448 265682 377460
rect 272518 377448 272524 377460
rect 265676 377420 272524 377448
rect 265676 377408 265682 377420
rect 272518 377408 272524 377420
rect 272576 377408 272582 377460
rect 438762 375980 438768 376032
rect 438820 376020 438826 376032
rect 449894 376020 449900 376032
rect 438820 375992 449900 376020
rect 438820 375980 438826 375992
rect 449894 375980 449900 375992
rect 449952 375980 449958 376032
rect 427906 373260 427912 373312
rect 427964 373300 427970 373312
rect 438762 373300 438768 373312
rect 427964 373272 438768 373300
rect 427964 373260 427970 373272
rect 438762 373260 438768 373272
rect 438820 373260 438826 373312
rect 426342 369928 426348 369980
rect 426400 369968 426406 369980
rect 427906 369968 427912 369980
rect 426400 369940 427912 369968
rect 426400 369928 426406 369940
rect 427906 369928 427912 369940
rect 427964 369928 427970 369980
rect 133138 368432 133144 368484
rect 133196 368472 133202 368484
rect 138014 368472 138020 368484
rect 133196 368444 138020 368472
rect 133196 368432 133202 368444
rect 138014 368432 138020 368444
rect 138072 368432 138078 368484
rect 420178 367752 420184 367804
rect 420236 367792 420242 367804
rect 426342 367792 426348 367804
rect 420236 367764 426348 367792
rect 420236 367752 420242 367764
rect 426342 367752 426348 367764
rect 426400 367752 426406 367804
rect 138014 365644 138020 365696
rect 138072 365684 138078 365696
rect 141418 365684 141424 365696
rect 138072 365656 141424 365684
rect 138072 365644 138078 365656
rect 141418 365644 141424 365656
rect 141476 365644 141482 365696
rect 417510 358708 417516 358760
rect 417568 358748 417574 358760
rect 420178 358748 420184 358760
rect 417568 358720 420184 358748
rect 417568 358708 417574 358720
rect 420178 358708 420184 358720
rect 420236 358708 420242 358760
rect 72602 355308 72608 355360
rect 72660 355348 72666 355360
rect 506566 355348 506572 355360
rect 72660 355320 506572 355348
rect 72660 355308 72666 355320
rect 506566 355308 506572 355320
rect 506624 355308 506630 355360
rect 141418 354696 141424 354748
rect 141476 354736 141482 354748
rect 144178 354736 144184 354748
rect 141476 354708 144184 354736
rect 141476 354696 141482 354708
rect 144178 354696 144184 354708
rect 144236 354696 144242 354748
rect 498838 353200 498844 353252
rect 498896 353240 498902 353252
rect 580166 353240 580172 353252
rect 498896 353212 580172 353240
rect 498896 353200 498902 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 272518 351160 272524 351212
rect 272576 351200 272582 351212
rect 287698 351200 287704 351212
rect 272576 351172 287704 351200
rect 272576 351160 272582 351172
rect 287698 351160 287704 351172
rect 287756 351160 287762 351212
rect 410518 347012 410524 347064
rect 410576 347052 410582 347064
rect 417510 347052 417516 347064
rect 410576 347024 417516 347052
rect 410576 347012 410582 347024
rect 417510 347012 417516 347024
rect 417568 347012 417574 347064
rect 56962 345652 56968 345704
rect 57020 345692 57026 345704
rect 288526 345692 288532 345704
rect 57020 345664 288532 345692
rect 57020 345652 57026 345664
rect 288526 345652 288532 345664
rect 288584 345652 288590 345704
rect 242802 344972 242808 345024
rect 242860 345012 242866 345024
rect 410518 345012 410524 345024
rect 242860 344984 410524 345012
rect 242860 344972 242866 344984
rect 410518 344972 410524 344984
rect 410576 344972 410582 345024
rect 76558 344292 76564 344344
rect 76616 344332 76622 344344
rect 494698 344332 494704 344344
rect 76616 344304 494704 344332
rect 76616 344292 76622 344304
rect 494698 344292 494704 344304
rect 494756 344292 494762 344344
rect 263594 343952 263600 344004
rect 263652 343992 263658 344004
rect 284294 343992 284300 344004
rect 263652 343964 284300 343992
rect 263652 343952 263658 343964
rect 284294 343952 284300 343964
rect 284352 343952 284358 344004
rect 256694 343884 256700 343936
rect 256752 343924 256758 343936
rect 280246 343924 280252 343936
rect 256752 343896 280252 343924
rect 256752 343884 256758 343896
rect 280246 343884 280252 343896
rect 280304 343884 280310 343936
rect 253198 343816 253204 343868
rect 253256 343856 253262 343868
rect 283190 343856 283196 343868
rect 253256 343828 283196 343856
rect 253256 343816 253262 343828
rect 283190 343816 283196 343828
rect 283248 343816 283254 343868
rect 255314 343748 255320 343800
rect 255372 343788 255378 343800
rect 287514 343788 287520 343800
rect 255372 343760 287520 343788
rect 255372 343748 255378 343760
rect 287514 343748 287520 343760
rect 287572 343748 287578 343800
rect 220170 343680 220176 343732
rect 220228 343720 220234 343732
rect 285950 343720 285956 343732
rect 220228 343692 285956 343720
rect 220228 343680 220234 343692
rect 285950 343680 285956 343692
rect 286008 343680 286014 343732
rect 144178 343612 144184 343664
rect 144236 343652 144242 343664
rect 147582 343652 147588 343664
rect 144236 343624 147588 343652
rect 144236 343612 144242 343624
rect 147582 343612 147588 343624
rect 147640 343612 147646 343664
rect 220078 343612 220084 343664
rect 220136 343652 220142 343664
rect 286042 343652 286048 343664
rect 220136 343624 286048 343652
rect 220136 343612 220142 343624
rect 286042 343612 286048 343624
rect 286100 343612 286106 343664
rect 251082 343068 251088 343120
rect 251140 343108 251146 343120
rect 284386 343108 284392 343120
rect 251140 343080 284392 343108
rect 251140 343068 251146 343080
rect 284386 343068 284392 343080
rect 284444 343068 284450 343120
rect 249702 343000 249708 343052
rect 249760 343040 249766 343052
rect 283282 343040 283288 343052
rect 249760 343012 283288 343040
rect 249760 343000 249766 343012
rect 283282 343000 283288 343012
rect 283340 343000 283346 343052
rect 245654 342932 245660 342984
rect 245712 342972 245718 342984
rect 283098 342972 283104 342984
rect 245712 342944 283104 342972
rect 245712 342932 245718 342944
rect 283098 342932 283104 342944
rect 283156 342932 283162 342984
rect 247034 342864 247040 342916
rect 247092 342904 247098 342916
rect 284478 342904 284484 342916
rect 247092 342876 284484 342904
rect 247092 342864 247098 342876
rect 284478 342864 284484 342876
rect 284536 342864 284542 342916
rect 243538 342796 243544 342848
rect 243596 342836 243602 342848
rect 285674 342836 285680 342848
rect 243596 342808 285680 342836
rect 243596 342796 243602 342808
rect 285674 342796 285680 342808
rect 285732 342796 285738 342848
rect 244274 342728 244280 342780
rect 244332 342768 244338 342780
rect 287606 342768 287612 342780
rect 244332 342740 287612 342768
rect 244332 342728 244338 342740
rect 287606 342728 287612 342740
rect 287664 342728 287670 342780
rect 240042 342660 240048 342712
rect 240100 342700 240106 342712
rect 283006 342700 283012 342712
rect 240100 342672 283012 342700
rect 240100 342660 240106 342672
rect 283006 342660 283012 342672
rect 283064 342660 283070 342712
rect 231210 342592 231216 342644
rect 231268 342632 231274 342644
rect 281534 342632 281540 342644
rect 231268 342604 281540 342632
rect 231268 342592 231274 342604
rect 281534 342592 281540 342604
rect 281592 342592 281598 342644
rect 231394 342524 231400 342576
rect 231452 342564 231458 342576
rect 284938 342564 284944 342576
rect 231452 342536 284944 342564
rect 231452 342524 231458 342536
rect 284938 342524 284944 342536
rect 284996 342524 285002 342576
rect 226334 342456 226340 342508
rect 226392 342496 226398 342508
rect 284846 342496 284852 342508
rect 226392 342468 284852 342496
rect 226392 342456 226398 342468
rect 284846 342456 284852 342468
rect 284904 342456 284910 342508
rect 223022 342388 223028 342440
rect 223080 342428 223086 342440
rect 283558 342428 283564 342440
rect 223080 342400 283564 342428
rect 223080 342388 223086 342400
rect 283558 342388 283564 342400
rect 283616 342388 283622 342440
rect 226610 342320 226616 342372
rect 226668 342360 226674 342372
rect 287422 342360 287428 342372
rect 226668 342332 287428 342360
rect 226668 342320 226674 342332
rect 287422 342320 287428 342332
rect 287480 342320 287486 342372
rect 220262 342252 220268 342304
rect 220320 342292 220326 342304
rect 285858 342292 285864 342304
rect 220320 342264 285864 342292
rect 220320 342252 220326 342264
rect 285858 342252 285864 342264
rect 285916 342252 285922 342304
rect 240042 341776 240048 341828
rect 240100 341816 240106 341828
rect 280614 341816 280620 341828
rect 240100 341788 280620 341816
rect 240100 341776 240106 341788
rect 280614 341776 280620 341788
rect 280672 341776 280678 341828
rect 237466 341708 237472 341760
rect 237524 341748 237530 341760
rect 280338 341748 280344 341760
rect 237524 341720 280344 341748
rect 237524 341708 237530 341720
rect 280338 341708 280344 341720
rect 280396 341708 280402 341760
rect 58618 341640 58624 341692
rect 58676 341680 58682 341692
rect 287054 341680 287060 341692
rect 58676 341652 287060 341680
rect 58676 341640 58682 341652
rect 287054 341640 287060 341652
rect 287112 341640 287118 341692
rect 236638 341572 236644 341624
rect 236696 341612 236702 341624
rect 490742 341612 490748 341624
rect 236696 341584 490748 341612
rect 236696 341572 236702 341584
rect 490742 341572 490748 341584
rect 490800 341572 490806 341624
rect 236914 341504 236920 341556
rect 236972 341544 236978 341556
rect 507302 341544 507308 341556
rect 236972 341516 507308 341544
rect 236972 341504 236978 341516
rect 507302 341504 507308 341516
rect 507360 341504 507366 341556
rect 237374 341436 237380 341488
rect 237432 341476 237438 341488
rect 280706 341476 280712 341488
rect 237432 341448 280712 341476
rect 237432 341436 237438 341448
rect 280706 341436 280712 341448
rect 280764 341436 280770 341488
rect 240778 341368 240784 341420
rect 240836 341408 240842 341420
rect 291838 341408 291844 341420
rect 240836 341380 291844 341408
rect 240836 341368 240842 341380
rect 291838 341368 291844 341380
rect 291896 341368 291902 341420
rect 227806 341300 227812 341352
rect 227864 341340 227870 341352
rect 284754 341340 284760 341352
rect 227864 341312 284760 341340
rect 227864 341300 227870 341312
rect 284754 341300 284760 341312
rect 284812 341300 284818 341352
rect 225690 341232 225696 341284
rect 225748 341272 225754 341284
rect 284570 341272 284576 341284
rect 225748 341244 284576 341272
rect 225748 341232 225754 341244
rect 284570 341232 284576 341244
rect 284628 341232 284634 341284
rect 223114 341164 223120 341216
rect 223172 341204 223178 341216
rect 283466 341204 283472 341216
rect 223172 341176 283472 341204
rect 223172 341164 223178 341176
rect 283466 341164 283472 341176
rect 283524 341164 283530 341216
rect 224954 341096 224960 341148
rect 225012 341136 225018 341148
rect 291378 341136 291384 341148
rect 225012 341108 291384 341136
rect 225012 341096 225018 341108
rect 291378 341096 291384 341108
rect 291436 341096 291442 341148
rect 225046 341028 225052 341080
rect 225104 341068 225110 341080
rect 291286 341068 291292 341080
rect 225104 341040 291292 341068
rect 225104 341028 225110 341040
rect 291286 341028 291292 341040
rect 291344 341028 291350 341080
rect 227714 340960 227720 341012
rect 227772 341000 227778 341012
rect 295334 341000 295340 341012
rect 227772 340972 295340 341000
rect 227772 340960 227778 340972
rect 295334 340960 295340 340972
rect 295392 340960 295398 341012
rect 225138 340892 225144 340944
rect 225196 340932 225202 340944
rect 292574 340932 292580 340944
rect 225196 340904 292580 340932
rect 225196 340892 225202 340904
rect 292574 340892 292580 340904
rect 292632 340892 292638 340944
rect 147582 340824 147588 340876
rect 147640 340864 147646 340876
rect 154482 340864 154488 340876
rect 147640 340836 154488 340864
rect 147640 340824 147646 340836
rect 154482 340824 154488 340836
rect 154540 340824 154546 340876
rect 239858 340348 239864 340400
rect 239916 340388 239922 340400
rect 280982 340388 280988 340400
rect 239916 340360 280988 340388
rect 239916 340348 239922 340360
rect 280982 340348 280988 340360
rect 281040 340348 281046 340400
rect 238386 340280 238392 340332
rect 238444 340320 238450 340332
rect 502978 340320 502984 340332
rect 238444 340292 502984 340320
rect 238444 340280 238450 340292
rect 502978 340280 502984 340292
rect 503036 340280 503042 340332
rect 237098 340212 237104 340264
rect 237156 340252 237162 340264
rect 580350 340252 580356 340264
rect 237156 340224 580356 340252
rect 237156 340212 237162 340224
rect 580350 340212 580356 340224
rect 580408 340212 580414 340264
rect 79318 340144 79324 340196
rect 79376 340184 79382 340196
rect 79778 340184 79784 340196
rect 79376 340156 79784 340184
rect 79376 340144 79382 340156
rect 79778 340144 79784 340156
rect 79836 340184 79842 340196
rect 503714 340184 503720 340196
rect 79836 340156 503720 340184
rect 79836 340144 79842 340156
rect 503714 340144 503720 340156
rect 503772 340144 503778 340196
rect 237466 340076 237472 340128
rect 237524 340116 237530 340128
rect 280430 340116 280436 340128
rect 237524 340088 280436 340116
rect 237524 340076 237530 340088
rect 280430 340076 280436 340088
rect 280488 340076 280494 340128
rect 237558 340008 237564 340060
rect 237616 340048 237622 340060
rect 280798 340048 280804 340060
rect 237616 340020 280804 340048
rect 237616 340008 237622 340020
rect 280798 340008 280804 340020
rect 280856 340008 280862 340060
rect 239950 339940 239956 339992
rect 240008 339980 240014 339992
rect 285030 339980 285036 339992
rect 240008 339952 285036 339980
rect 240008 339940 240014 339952
rect 285030 339940 285036 339952
rect 285088 339940 285094 339992
rect 240042 339872 240048 339924
rect 240100 339912 240106 339924
rect 285766 339912 285772 339924
rect 240100 339884 285772 339912
rect 240100 339872 240106 339884
rect 285766 339872 285772 339884
rect 285824 339872 285830 339924
rect 237374 339804 237380 339856
rect 237432 339844 237438 339856
rect 284662 339844 284668 339856
rect 237432 339816 284668 339844
rect 237432 339804 237438 339816
rect 284662 339804 284668 339816
rect 284720 339804 284726 339856
rect 228450 339736 228456 339788
rect 228508 339776 228514 339788
rect 281718 339776 281724 339788
rect 228508 339748 281724 339776
rect 228508 339736 228514 339748
rect 281718 339736 281724 339748
rect 281776 339736 281782 339788
rect 225874 339668 225880 339720
rect 225932 339708 225938 339720
rect 283374 339708 283380 339720
rect 225932 339680 283380 339708
rect 225932 339668 225938 339680
rect 283374 339668 283380 339680
rect 283432 339668 283438 339720
rect 223482 339600 223488 339652
rect 223540 339640 223546 339652
rect 283650 339640 283656 339652
rect 223540 339612 283656 339640
rect 223540 339600 223546 339612
rect 283650 339600 283656 339612
rect 283708 339600 283714 339652
rect 223390 339532 223396 339584
rect 223448 339572 223454 339584
rect 283742 339572 283748 339584
rect 223448 339544 283748 339572
rect 223448 339532 223454 339544
rect 283742 339532 283748 339544
rect 283800 339532 283806 339584
rect 235718 339464 235724 339516
rect 235776 339504 235782 339516
rect 580258 339504 580264 339516
rect 235776 339476 580264 339504
rect 235776 339464 235782 339476
rect 580258 339464 580264 339476
rect 580316 339464 580322 339516
rect 231302 339396 231308 339448
rect 231360 339436 231366 339448
rect 281626 339436 281632 339448
rect 231360 339408 281632 339436
rect 231360 339396 231366 339408
rect 281626 339396 281632 339408
rect 281684 339396 281690 339448
rect 239122 338512 239128 338564
rect 239180 338552 239186 338564
rect 239858 338552 239864 338564
rect 239180 338524 239864 338552
rect 239180 338512 239186 338524
rect 239858 338512 239864 338524
rect 239916 338512 239922 338564
rect 238018 337356 238024 337408
rect 238076 337396 238082 337408
rect 238386 337396 238392 337408
rect 238076 337368 238392 337396
rect 238076 337356 238082 337368
rect 238386 337356 238392 337368
rect 238444 337356 238450 337408
rect 154482 336676 154488 336728
rect 154540 336716 154546 336728
rect 158806 336716 158812 336728
rect 154540 336688 158812 336716
rect 154540 336676 154546 336688
rect 158806 336676 158812 336688
rect 158864 336676 158870 336728
rect 158806 332392 158812 332444
rect 158864 332432 158870 332444
rect 162118 332432 162124 332444
rect 158864 332404 162124 332432
rect 158864 332392 158870 332404
rect 162118 332392 162124 332404
rect 162176 332392 162182 332444
rect 162118 321580 162124 321632
rect 162176 321620 162182 321632
rect 166258 321620 166264 321632
rect 162176 321592 166264 321620
rect 162176 321580 162182 321592
rect 166258 321580 166264 321592
rect 166316 321580 166322 321632
rect 94038 312536 94044 312588
rect 94096 312576 94102 312588
rect 158714 312576 158720 312588
rect 94096 312548 158720 312576
rect 94096 312536 94102 312548
rect 158714 312536 158720 312548
rect 158772 312536 158778 312588
rect 92382 311108 92388 311160
rect 92440 311148 92446 311160
rect 154574 311148 154580 311160
rect 92440 311120 154580 311148
rect 92440 311108 92446 311120
rect 154574 311108 154580 311120
rect 154632 311108 154638 311160
rect 90726 309748 90732 309800
rect 90784 309788 90790 309800
rect 150434 309788 150440 309800
rect 90784 309760 150440 309788
rect 90784 309748 90790 309760
rect 150434 309748 150440 309760
rect 150492 309748 150498 309800
rect 87414 308388 87420 308440
rect 87472 308428 87478 308440
rect 143534 308428 143540 308440
rect 87472 308400 143540 308428
rect 87472 308388 87478 308400
rect 143534 308388 143540 308400
rect 143592 308388 143598 308440
rect 85758 307028 85764 307080
rect 85816 307068 85822 307080
rect 140774 307068 140780 307080
rect 85816 307040 140780 307068
rect 85816 307028 85822 307040
rect 140774 307028 140780 307040
rect 140832 307028 140838 307080
rect 82446 304240 82452 304292
rect 82504 304280 82510 304292
rect 132494 304280 132500 304292
rect 82504 304252 132500 304280
rect 82504 304240 82510 304252
rect 132494 304240 132500 304252
rect 132552 304240 132558 304292
rect 80790 302880 80796 302932
rect 80848 302920 80854 302932
rect 129734 302920 129740 302932
rect 80848 302892 129740 302920
rect 80848 302880 80854 302892
rect 129734 302880 129740 302892
rect 129792 302880 129798 302932
rect 75822 300092 75828 300144
rect 75880 300132 75886 300144
rect 119338 300132 119344 300144
rect 75880 300104 119344 300132
rect 75880 300092 75886 300104
rect 119338 300092 119344 300104
rect 119396 300092 119402 300144
rect 282178 299412 282184 299464
rect 282236 299452 282242 299464
rect 285030 299452 285036 299464
rect 282236 299424 285036 299452
rect 282236 299412 282242 299424
rect 285030 299412 285036 299424
rect 285088 299412 285094 299464
rect 74166 297372 74172 297424
rect 74224 297412 74230 297424
rect 115198 297412 115204 297424
rect 74224 297384 115204 297412
rect 74224 297372 74230 297384
rect 115198 297372 115204 297384
rect 115256 297372 115262 297424
rect 166258 292544 166264 292596
rect 166316 292584 166322 292596
rect 169018 292584 169024 292596
rect 166316 292556 169024 292584
rect 166316 292544 166322 292556
rect 169018 292544 169024 292556
rect 169076 292544 169082 292596
rect 496722 291796 496728 291848
rect 496780 291836 496786 291848
rect 503714 291836 503720 291848
rect 496780 291808 503720 291836
rect 496780 291796 496786 291808
rect 503714 291796 503720 291808
rect 503772 291796 503778 291848
rect 282178 289756 282184 289808
rect 282236 289796 282242 289808
rect 284938 289796 284944 289808
rect 282236 289768 284944 289796
rect 282236 289756 282242 289768
rect 284938 289756 284944 289768
rect 284996 289756 285002 289808
rect 282086 288328 282092 288380
rect 282144 288368 282150 288380
rect 284846 288368 284852 288380
rect 282144 288340 284852 288368
rect 282144 288328 282150 288340
rect 284846 288328 284852 288340
rect 284904 288328 284910 288380
rect 282730 288260 282736 288312
rect 282788 288300 282794 288312
rect 286042 288300 286048 288312
rect 282788 288272 286048 288300
rect 282788 288260 282794 288272
rect 286042 288260 286048 288272
rect 286100 288260 286106 288312
rect 282638 286696 282644 286748
rect 282696 286736 282702 286748
rect 285950 286736 285956 286748
rect 282696 286708 285956 286736
rect 282696 286696 282702 286708
rect 285950 286696 285956 286708
rect 286008 286696 286014 286748
rect 281534 285608 281540 285660
rect 281592 285648 281598 285660
rect 283742 285648 283748 285660
rect 281592 285620 283748 285648
rect 281592 285608 281598 285620
rect 283742 285608 283748 285620
rect 283800 285608 283806 285660
rect 282638 285540 282644 285592
rect 282696 285580 282702 285592
rect 285858 285580 285864 285592
rect 282696 285552 285864 285580
rect 282696 285540 282702 285552
rect 285858 285540 285864 285552
rect 285916 285540 285922 285592
rect 282086 284248 282092 284300
rect 282144 284288 282150 284300
rect 284754 284288 284760 284300
rect 282144 284260 284760 284288
rect 282144 284248 282150 284260
rect 284754 284248 284760 284260
rect 284812 284248 284818 284300
rect 77478 282140 77484 282192
rect 77536 282180 77542 282192
rect 122834 282180 122840 282192
rect 77536 282152 122840 282180
rect 77536 282140 77542 282152
rect 122834 282140 122840 282152
rect 122892 282140 122898 282192
rect 281994 281460 282000 281512
rect 282052 281500 282058 281512
rect 284570 281500 284576 281512
rect 282052 281472 284576 281500
rect 282052 281460 282058 281472
rect 284570 281460 284576 281472
rect 284628 281460 284634 281512
rect 281994 280100 282000 280152
rect 282052 280140 282058 280152
rect 284662 280140 284668 280152
rect 282052 280112 284668 280140
rect 282052 280100 282058 280112
rect 284662 280100 284668 280112
rect 284720 280100 284726 280152
rect 70854 279420 70860 279472
rect 70912 279460 70918 279472
rect 108298 279460 108304 279472
rect 70912 279432 108304 279460
rect 70912 279420 70918 279432
rect 108298 279420 108304 279432
rect 108356 279420 108362 279472
rect 169018 279420 169024 279472
rect 169076 279460 169082 279472
rect 182818 279460 182824 279472
rect 169076 279432 182824 279460
rect 169076 279420 169082 279432
rect 182818 279420 182824 279432
rect 182876 279420 182882 279472
rect 282822 277448 282828 277500
rect 282880 277488 282886 277500
rect 288618 277488 288624 277500
rect 282880 277460 288624 277488
rect 282880 277448 282886 277460
rect 288618 277448 288624 277460
rect 288676 277448 288682 277500
rect 282822 276088 282828 276140
rect 282880 276128 282886 276140
rect 288710 276128 288716 276140
rect 282880 276100 288716 276128
rect 282880 276088 282886 276100
rect 288710 276088 288716 276100
rect 288768 276088 288774 276140
rect 282730 276020 282736 276072
rect 282788 276060 282794 276072
rect 289906 276060 289912 276072
rect 282788 276032 289912 276060
rect 282788 276020 282794 276032
rect 289906 276020 289912 276032
rect 289964 276020 289970 276072
rect 493962 275272 493968 275324
rect 494020 275312 494026 275324
rect 506474 275312 506480 275324
rect 494020 275284 506480 275312
rect 494020 275272 494026 275284
rect 506474 275272 506480 275284
rect 506532 275272 506538 275324
rect 282822 274660 282828 274712
rect 282880 274700 282886 274712
rect 287146 274700 287152 274712
rect 282880 274672 287152 274700
rect 282880 274660 282886 274672
rect 287146 274660 287152 274672
rect 287204 274660 287210 274712
rect 282822 273300 282828 273352
rect 282880 273340 282886 273352
rect 287238 273340 287244 273352
rect 282880 273312 287244 273340
rect 282880 273300 282886 273312
rect 287238 273300 287244 273312
rect 287296 273300 287302 273352
rect 282730 273232 282736 273284
rect 282788 273272 282794 273284
rect 289998 273272 290004 273284
rect 282788 273244 290004 273272
rect 282788 273232 282794 273244
rect 289998 273232 290004 273244
rect 290056 273232 290062 273284
rect 282822 271872 282828 271924
rect 282880 271912 282886 271924
rect 287330 271912 287336 271924
rect 282880 271884 287336 271912
rect 282880 271872 282886 271884
rect 287330 271872 287336 271884
rect 287388 271872 287394 271924
rect 69198 271192 69204 271244
rect 69256 271232 69262 271244
rect 105630 271232 105636 271244
rect 69256 271204 105636 271232
rect 69256 271192 69262 271204
rect 105630 271192 105636 271204
rect 105688 271192 105694 271244
rect 89070 271124 89076 271176
rect 89128 271164 89134 271176
rect 147674 271164 147680 271176
rect 89128 271136 147680 271164
rect 89128 271124 89134 271136
rect 147674 271124 147680 271136
rect 147732 271124 147738 271176
rect 282822 270580 282828 270632
rect 282880 270620 282886 270632
rect 291562 270620 291568 270632
rect 282880 270592 291568 270620
rect 282880 270580 282886 270592
rect 291562 270580 291568 270592
rect 291620 270580 291626 270632
rect 282730 270512 282736 270564
rect 282788 270552 282794 270564
rect 291470 270552 291476 270564
rect 282788 270524 291476 270552
rect 282788 270512 282794 270524
rect 291470 270512 291476 270524
rect 291528 270512 291534 270564
rect 281902 270444 281908 270496
rect 281960 270484 281966 270496
rect 284478 270484 284484 270496
rect 281960 270456 284484 270484
rect 281960 270444 281966 270456
rect 284478 270444 284484 270456
rect 284536 270444 284542 270496
rect 281902 267656 281908 267708
rect 281960 267696 281966 267708
rect 284386 267696 284392 267708
rect 281960 267668 284392 267696
rect 281960 267656 281966 267668
rect 284386 267656 284392 267668
rect 284444 267656 284450 267708
rect 281810 266296 281816 266348
rect 281868 266336 281874 266348
rect 284294 266336 284300 266348
rect 281868 266308 284300 266336
rect 281868 266296 281874 266308
rect 284294 266296 284300 266308
rect 284352 266296 284358 266348
rect 54662 262964 54668 263016
rect 54720 263004 54726 263016
rect 72418 263004 72424 263016
rect 54720 262976 72424 263004
rect 54720 262964 54726 262976
rect 72418 262964 72424 262976
rect 72476 262964 72482 263016
rect 56318 262896 56324 262948
rect 56376 262936 56382 262948
rect 76558 262936 76564 262948
rect 56376 262908 76564 262936
rect 56376 262896 56382 262908
rect 76558 262896 76564 262908
rect 76616 262896 76622 262948
rect 57882 262828 57888 262880
rect 57940 262868 57946 262880
rect 79318 262868 79324 262880
rect 57940 262840 79324 262868
rect 57940 262828 57946 262840
rect 79318 262828 79324 262840
rect 79376 262828 79382 262880
rect 282822 262148 282828 262200
rect 282880 262188 282886 262200
rect 287606 262188 287612 262200
rect 282880 262160 287612 262188
rect 282880 262148 282886 262160
rect 287606 262148 287612 262160
rect 287664 262148 287670 262200
rect 39942 261468 39948 261520
rect 40000 261508 40006 261520
rect 233970 261508 233976 261520
rect 40000 261480 233976 261508
rect 40000 261468 40006 261480
rect 233970 261468 233976 261480
rect 234028 261468 234034 261520
rect 11698 260856 11704 260908
rect 11756 260896 11762 260908
rect 102134 260896 102140 260908
rect 11756 260868 102140 260896
rect 11756 260856 11762 260868
rect 102134 260856 102140 260868
rect 102192 260856 102198 260908
rect 282546 260788 282552 260840
rect 282604 260828 282610 260840
rect 285674 260828 285680 260840
rect 282604 260800 285680 260828
rect 282604 260788 282610 260800
rect 285674 260788 285680 260800
rect 285732 260788 285738 260840
rect 282546 257456 282552 257508
rect 282604 257496 282610 257508
rect 285766 257496 285772 257508
rect 282604 257468 285772 257496
rect 282604 257456 282610 257468
rect 285766 257456 285772 257468
rect 285824 257456 285830 257508
rect 282822 256640 282828 256692
rect 282880 256680 282886 256692
rect 287514 256680 287520 256692
rect 282880 256652 287520 256680
rect 282880 256640 282886 256652
rect 287514 256640 287520 256652
rect 287572 256640 287578 256692
rect 282822 253852 282828 253904
rect 282880 253892 282886 253904
rect 287422 253892 287428 253904
rect 282880 253864 287428 253892
rect 282880 253852 282886 253864
rect 287422 253852 287428 253864
rect 287480 253852 287486 253904
rect 182818 249704 182824 249756
rect 182876 249744 182882 249756
rect 189718 249744 189724 249756
rect 182876 249716 189724 249744
rect 182876 249704 182882 249716
rect 189718 249704 189724 249716
rect 189776 249704 189782 249756
rect 496722 245556 496728 245608
rect 496780 245596 496786 245608
rect 580166 245596 580172 245608
rect 496780 245568 580172 245596
rect 496780 245556 496786 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 282822 242904 282828 242956
rect 282880 242944 282886 242956
rect 288894 242944 288900 242956
rect 282880 242916 288900 242944
rect 282880 242904 282886 242916
rect 288894 242904 288900 242916
rect 288952 242904 288958 242956
rect 189718 235220 189724 235272
rect 189776 235260 189782 235272
rect 207658 235260 207664 235272
rect 189776 235232 207664 235260
rect 189776 235220 189782 235232
rect 207658 235220 207664 235232
rect 207716 235220 207722 235272
rect 282178 229100 282184 229152
rect 282236 229140 282242 229152
rect 284938 229140 284944 229152
rect 282236 229112 284944 229140
rect 282236 229100 282242 229112
rect 284938 229100 284944 229112
rect 284996 229100 285002 229152
rect 282270 227740 282276 227792
rect 282328 227780 282334 227792
rect 285122 227780 285128 227792
rect 282328 227752 285128 227780
rect 282328 227740 282334 227752
rect 285122 227740 285128 227752
rect 285180 227740 285186 227792
rect 282822 219444 282828 219496
rect 282880 219484 282886 219496
rect 290458 219484 290464 219496
rect 282880 219456 290464 219484
rect 282880 219444 282886 219456
rect 290458 219444 290464 219456
rect 290516 219444 290522 219496
rect 3418 215228 3424 215280
rect 3476 215268 3482 215280
rect 11698 215268 11704 215280
rect 3476 215240 11704 215268
rect 3476 215228 3482 215240
rect 11698 215228 11704 215240
rect 11756 215228 11762 215280
rect 111058 214548 111064 214600
rect 111116 214588 111122 214600
rect 158714 214588 158720 214600
rect 111116 214560 158720 214588
rect 111116 214548 111122 214560
rect 158714 214548 158720 214560
rect 158772 214548 158778 214600
rect 233878 213936 233884 213988
rect 233936 213976 233942 213988
rect 237374 213976 237380 213988
rect 233936 213948 237380 213976
rect 233936 213936 233942 213948
rect 237374 213936 237380 213948
rect 237432 213936 237438 213988
rect 207658 211760 207664 211812
rect 207716 211800 207722 211812
rect 218698 211800 218704 211812
rect 207716 211772 218704 211800
rect 207716 211760 207722 211772
rect 218698 211760 218704 211772
rect 218756 211760 218762 211812
rect 282822 211148 282828 211200
rect 282880 211188 282886 211200
rect 288986 211188 288992 211200
rect 282880 211160 288992 211188
rect 282880 211148 282886 211160
rect 288986 211148 288992 211160
rect 289044 211148 289050 211200
rect 494698 206932 494704 206984
rect 494756 206972 494762 206984
rect 580166 206972 580172 206984
rect 494756 206944 580172 206972
rect 494756 206932 494762 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 282822 204280 282828 204332
rect 282880 204320 282886 204332
rect 291746 204320 291752 204332
rect 282880 204292 291752 204320
rect 282880 204280 282886 204292
rect 291746 204280 291752 204292
rect 291804 204280 291810 204332
rect 233970 201424 233976 201476
rect 234028 201464 234034 201476
rect 237374 201464 237380 201476
rect 234028 201436 237380 201464
rect 234028 201424 234034 201436
rect 237374 201424 237380 201436
rect 237432 201424 237438 201476
rect 48222 200064 48228 200116
rect 48280 200104 48286 200116
rect 110414 200104 110420 200116
rect 48280 200076 110420 200104
rect 48280 200064 48286 200076
rect 110414 200064 110420 200076
rect 110472 200104 110478 200116
rect 111058 200104 111064 200116
rect 110472 200076 111064 200104
rect 110472 200064 110478 200076
rect 111058 200064 111064 200076
rect 111116 200064 111122 200116
rect 218698 199996 218704 200048
rect 218756 200036 218762 200048
rect 237374 200036 237380 200048
rect 218756 200008 237380 200036
rect 218756 199996 218762 200008
rect 237374 199996 237380 200008
rect 237432 199996 237438 200048
rect 104894 199928 104900 199980
rect 104952 199968 104958 199980
rect 231026 199968 231032 199980
rect 104952 199940 231032 199968
rect 104952 199928 104958 199940
rect 231026 199928 231032 199940
rect 231084 199928 231090 199980
rect 106274 199860 106280 199912
rect 106332 199900 106338 199912
rect 231302 199900 231308 199912
rect 106332 199872 231308 199900
rect 106332 199860 106338 199872
rect 231302 199860 231308 199872
rect 231360 199860 231366 199912
rect 95234 199792 95240 199844
rect 95292 199832 95298 199844
rect 220078 199832 220084 199844
rect 95292 199804 220084 199832
rect 95292 199792 95298 199804
rect 220078 199792 220084 199804
rect 220136 199792 220142 199844
rect 100662 199724 100668 199776
rect 100720 199764 100726 199776
rect 220170 199764 220176 199776
rect 100720 199736 220176 199764
rect 100720 199724 100726 199736
rect 220170 199724 220176 199736
rect 220228 199724 220234 199776
rect 103422 199656 103428 199708
rect 103480 199696 103486 199708
rect 220262 199696 220268 199708
rect 103480 199668 220268 199696
rect 103480 199656 103486 199668
rect 220262 199656 220268 199668
rect 220320 199656 220326 199708
rect 94498 199588 94504 199640
rect 94556 199628 94562 199640
rect 223022 199628 223028 199640
rect 94556 199600 223028 199628
rect 94556 199588 94562 199600
rect 223022 199588 223028 199600
rect 223080 199588 223086 199640
rect 107654 199520 107660 199572
rect 107712 199560 107718 199572
rect 228450 199560 228456 199572
rect 107712 199532 228456 199560
rect 107712 199520 107718 199532
rect 228450 199520 228456 199532
rect 228508 199520 228514 199572
rect 88334 198636 88340 198688
rect 88392 198676 88398 198688
rect 225874 198676 225880 198688
rect 88392 198648 225880 198676
rect 88392 198636 88398 198648
rect 225874 198636 225880 198648
rect 225932 198636 225938 198688
rect 86954 198568 86960 198620
rect 87012 198608 87018 198620
rect 223482 198608 223488 198620
rect 87012 198580 223488 198608
rect 87012 198568 87018 198580
rect 223482 198568 223488 198580
rect 223540 198568 223546 198620
rect 97994 198500 98000 198552
rect 98052 198540 98058 198552
rect 225690 198540 225696 198552
rect 98052 198512 225696 198540
rect 98052 198500 98058 198512
rect 225690 198500 225696 198512
rect 225748 198500 225754 198552
rect 96614 198432 96620 198484
rect 96672 198472 96678 198484
rect 223114 198472 223120 198484
rect 96672 198444 223120 198472
rect 96672 198432 96678 198444
rect 223114 198432 223120 198444
rect 223172 198432 223178 198484
rect 104158 198364 104164 198416
rect 104216 198404 104222 198416
rect 223390 198404 223396 198416
rect 104216 198376 223396 198404
rect 104216 198364 104222 198376
rect 223390 198364 223396 198376
rect 223448 198364 223454 198416
rect 85574 197684 85580 197736
rect 85632 197724 85638 197736
rect 238662 197724 238668 197736
rect 85632 197696 238668 197724
rect 85632 197684 85638 197696
rect 238662 197684 238668 197696
rect 238720 197684 238726 197736
rect 78582 197616 78588 197668
rect 78640 197656 78646 197668
rect 235442 197656 235448 197668
rect 78640 197628 235448 197656
rect 78640 197616 78646 197628
rect 235442 197616 235448 197628
rect 235500 197616 235506 197668
rect 79318 197548 79324 197600
rect 79376 197588 79382 197600
rect 238478 197588 238484 197600
rect 79376 197560 238484 197588
rect 79376 197548 79382 197560
rect 238478 197548 238484 197560
rect 238536 197548 238542 197600
rect 70394 197480 70400 197532
rect 70452 197520 70458 197532
rect 235350 197520 235356 197532
rect 70452 197492 235356 197520
rect 70452 197480 70458 197492
rect 235350 197480 235356 197492
rect 235408 197480 235414 197532
rect 73154 197412 73160 197464
rect 73212 197452 73218 197464
rect 238294 197452 238300 197464
rect 73212 197424 238300 197452
rect 73212 197412 73218 197424
rect 238294 197412 238300 197424
rect 238352 197412 238358 197464
rect 71774 197344 71780 197396
rect 71832 197384 71838 197396
rect 238202 197384 238208 197396
rect 71832 197356 238208 197384
rect 71832 197344 71838 197356
rect 238202 197344 238208 197356
rect 238260 197344 238266 197396
rect 287698 187688 287704 187740
rect 287756 187728 287762 187740
rect 291194 187728 291200 187740
rect 287756 187700 291200 187728
rect 287756 187688 287762 187700
rect 291194 187688 291200 187700
rect 291252 187688 291258 187740
rect 282454 178032 282460 178084
rect 282512 178072 282518 178084
rect 283742 178072 283748 178084
rect 282512 178044 283748 178072
rect 282512 178032 282518 178044
rect 283742 178032 283748 178044
rect 283800 178032 283806 178084
rect 282822 176672 282828 176724
rect 282880 176712 282886 176724
rect 289170 176712 289176 176724
rect 282880 176684 289176 176712
rect 282880 176672 282886 176684
rect 289170 176672 289176 176684
rect 289228 176672 289234 176724
rect 282822 172456 282828 172508
rect 282880 172496 282886 172508
rect 295334 172496 295340 172508
rect 282880 172468 295340 172496
rect 282880 172456 282886 172468
rect 295334 172456 295340 172468
rect 295392 172456 295398 172508
rect 282730 172388 282736 172440
rect 282788 172428 282794 172440
rect 291378 172428 291384 172440
rect 282788 172400 291384 172428
rect 282788 172388 282794 172400
rect 291378 172388 291384 172400
rect 291436 172388 291442 172440
rect 282822 171028 282828 171080
rect 282880 171068 282886 171080
rect 292574 171068 292580 171080
rect 282880 171040 292580 171068
rect 282880 171028 282886 171040
rect 292574 171028 292580 171040
rect 292632 171028 292638 171080
rect 282822 169668 282828 169720
rect 282880 169708 282886 169720
rect 291286 169708 291292 169720
rect 282880 169680 291292 169708
rect 282880 169668 282886 169680
rect 291286 169668 291292 169680
rect 291344 169668 291350 169720
rect 282822 169532 282828 169584
rect 282880 169572 282886 169584
rect 287054 169572 287060 169584
rect 282880 169544 287060 169572
rect 282880 169532 282886 169544
rect 287054 169532 287060 169544
rect 287112 169532 287118 169584
rect 282730 168308 282736 168360
rect 282788 168348 282794 168360
rect 291194 168348 291200 168360
rect 282788 168320 291200 168348
rect 282788 168308 282794 168320
rect 291194 168308 291200 168320
rect 291252 168308 291258 168360
rect 282822 168240 282828 168292
rect 282880 168280 282886 168292
rect 288526 168280 288532 168292
rect 282880 168252 288532 168280
rect 282880 168240 282886 168252
rect 288526 168240 288532 168252
rect 288584 168240 288590 168292
rect 493962 166948 493968 167000
rect 494020 166988 494026 167000
rect 580166 166988 580172 167000
rect 494020 166960 580172 166988
rect 494020 166948 494026 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 232682 141992 232688 142044
rect 232740 142032 232746 142044
rect 236822 142032 236828 142044
rect 232740 142004 236828 142032
rect 232740 141992 232746 142004
rect 236822 141992 236828 142004
rect 236880 141992 236886 142044
rect 238478 140632 238484 140684
rect 238536 140672 238542 140684
rect 580442 140672 580448 140684
rect 238536 140644 580448 140672
rect 238536 140632 238542 140644
rect 580442 140632 580448 140644
rect 580500 140632 580506 140684
rect 237742 140564 237748 140616
rect 237800 140604 237806 140616
rect 580350 140604 580356 140616
rect 237800 140576 580356 140604
rect 237800 140564 237806 140576
rect 580350 140564 580356 140576
rect 580408 140564 580414 140616
rect 238570 140496 238576 140548
rect 238628 140536 238634 140548
rect 580258 140536 580264 140548
rect 238628 140508 580264 140536
rect 238628 140496 238634 140508
rect 580258 140496 580264 140508
rect 580316 140496 580322 140548
rect 239674 140428 239680 140480
rect 239732 140468 239738 140480
rect 580534 140468 580540 140480
rect 239732 140440 580540 140468
rect 239732 140428 239738 140440
rect 580534 140428 580540 140440
rect 580592 140428 580598 140480
rect 239582 140360 239588 140412
rect 239640 140400 239646 140412
rect 458818 140400 458824 140412
rect 239640 140372 458824 140400
rect 239640 140360 239646 140372
rect 458818 140360 458824 140372
rect 458876 140360 458882 140412
rect 235350 140292 235356 140344
rect 235408 140332 235414 140344
rect 291562 140332 291568 140344
rect 235408 140304 291568 140332
rect 235408 140292 235414 140304
rect 291562 140292 291568 140304
rect 291620 140292 291626 140344
rect 235442 140224 235448 140276
rect 235500 140264 235506 140276
rect 291470 140264 291476 140276
rect 235500 140236 291476 140264
rect 235500 140224 235506 140236
rect 291470 140224 291476 140236
rect 291528 140224 291534 140276
rect 235902 140156 235908 140208
rect 235960 140196 235966 140208
rect 289170 140196 289176 140208
rect 235960 140168 289176 140196
rect 235960 140156 235966 140168
rect 289170 140156 289176 140168
rect 289228 140156 289234 140208
rect 238018 140088 238024 140140
rect 238076 140128 238082 140140
rect 287238 140128 287244 140140
rect 238076 140100 287244 140128
rect 238076 140088 238082 140100
rect 287238 140088 287244 140100
rect 287296 140088 287302 140140
rect 238110 140020 238116 140072
rect 238168 140060 238174 140072
rect 287330 140060 287336 140072
rect 238168 140032 287336 140060
rect 238168 140020 238174 140032
rect 287330 140020 287336 140032
rect 287388 140020 287394 140072
rect 266906 139952 266912 140004
rect 266964 139992 266970 140004
rect 283742 139992 283748 140004
rect 266964 139964 283748 139992
rect 266964 139952 266970 139964
rect 283742 139952 283748 139964
rect 283800 139952 283806 140004
rect 238202 139340 238208 139392
rect 238260 139380 238266 139392
rect 470870 139380 470876 139392
rect 238260 139352 470876 139380
rect 238260 139340 238266 139352
rect 470870 139340 470876 139352
rect 470928 139340 470934 139392
rect 240778 139272 240784 139324
rect 240836 139312 240842 139324
rect 467282 139312 467288 139324
rect 240836 139284 467288 139312
rect 240836 139272 240842 139284
rect 467282 139272 467288 139284
rect 467340 139272 467346 139324
rect 205634 139204 205640 139256
rect 205692 139244 205698 139256
rect 288986 139244 288992 139256
rect 205692 139216 288992 139244
rect 205692 139204 205698 139216
rect 288986 139204 288992 139216
rect 289044 139204 289050 139256
rect 215294 139136 215300 139188
rect 215352 139176 215358 139188
rect 290458 139176 290464 139188
rect 215352 139148 290464 139176
rect 215352 139136 215358 139148
rect 290458 139136 290464 139148
rect 290516 139136 290522 139188
rect 218054 139068 218060 139120
rect 218112 139108 218118 139120
rect 282178 139108 282184 139120
rect 218112 139080 282184 139108
rect 218112 139068 218118 139080
rect 282178 139068 282184 139080
rect 282236 139068 282242 139120
rect 235902 139000 235908 139052
rect 235960 139040 235966 139052
rect 288710 139040 288716 139052
rect 235960 139012 288716 139040
rect 235960 139000 235966 139012
rect 288710 139000 288716 139012
rect 288768 139000 288774 139052
rect 235626 138932 235632 138984
rect 235684 138972 235690 138984
rect 287146 138972 287152 138984
rect 235684 138944 287152 138972
rect 235684 138932 235690 138944
rect 287146 138932 287152 138944
rect 287204 138932 287210 138984
rect 233142 138864 233148 138916
rect 233200 138904 233206 138916
rect 283374 138904 283380 138916
rect 233200 138876 283380 138904
rect 233200 138864 233206 138876
rect 283374 138864 283380 138876
rect 283432 138864 283438 138916
rect 238754 138796 238760 138848
rect 238812 138836 238818 138848
rect 288894 138836 288900 138848
rect 238812 138808 288900 138836
rect 238812 138796 238818 138808
rect 288894 138796 288900 138808
rect 288952 138796 288958 138848
rect 235810 138728 235816 138780
rect 235868 138768 235874 138780
rect 285122 138768 285128 138780
rect 235868 138740 285128 138768
rect 235868 138728 235874 138740
rect 285122 138728 285128 138740
rect 285180 138728 285186 138780
rect 235902 138660 235908 138712
rect 235960 138700 235966 138712
rect 284938 138700 284944 138712
rect 235960 138672 284944 138700
rect 235960 138660 235966 138672
rect 284938 138660 284944 138672
rect 284996 138660 285002 138712
rect 235718 138592 235724 138644
rect 235776 138632 235782 138644
rect 282086 138632 282092 138644
rect 235776 138604 282092 138632
rect 235776 138592 235782 138604
rect 282086 138592 282092 138604
rect 282144 138592 282150 138644
rect 251174 138524 251180 138576
rect 251232 138564 251238 138576
rect 280338 138564 280344 138576
rect 251232 138536 280344 138564
rect 251232 138524 251238 138536
rect 280338 138524 280344 138536
rect 280396 138524 280402 138576
rect 237374 137912 237380 137964
rect 237432 137952 237438 137964
rect 249794 137952 249800 137964
rect 237432 137924 249800 137952
rect 237432 137912 237438 137924
rect 249794 137912 249800 137924
rect 249852 137912 249858 137964
rect 262122 137912 262128 137964
rect 262180 137952 262186 137964
rect 288618 137952 288624 137964
rect 262180 137924 288624 137952
rect 262180 137912 262186 137924
rect 288618 137912 288624 137924
rect 288676 137912 288682 137964
rect 66162 137844 66168 137896
rect 66220 137884 66226 137896
rect 245010 137884 245016 137896
rect 66220 137856 245016 137884
rect 66220 137844 66226 137856
rect 245010 137844 245016 137856
rect 245068 137844 245074 137896
rect 247034 137844 247040 137896
rect 247092 137884 247098 137896
rect 250990 137884 250996 137896
rect 247092 137856 250996 137884
rect 247092 137844 247098 137856
rect 250990 137844 250996 137856
rect 251048 137844 251054 137896
rect 115842 137776 115848 137828
rect 115900 137816 115906 137828
rect 246206 137816 246212 137828
rect 115900 137788 246212 137816
rect 115900 137776 115906 137788
rect 246206 137776 246212 137788
rect 246264 137776 246270 137828
rect 118694 137708 118700 137760
rect 118752 137748 118758 137760
rect 247402 137748 247408 137760
rect 118752 137720 247408 137748
rect 118752 137708 118758 137720
rect 247402 137708 247408 137720
rect 247460 137708 247466 137760
rect 233142 137640 233148 137692
rect 233200 137680 233206 137692
rect 248598 137680 248604 137692
rect 233200 137652 248604 137680
rect 233200 137640 233206 137652
rect 248598 137640 248604 137652
rect 248656 137640 248662 137692
rect 44174 137572 44180 137624
rect 44232 137612 44238 137624
rect 243814 137612 243820 137624
rect 44232 137584 243820 137612
rect 44232 137572 44238 137584
rect 243814 137572 243820 137584
rect 243872 137572 243878 137624
rect 271138 136620 271144 136672
rect 271196 136660 271202 136672
rect 272518 136660 272524 136672
rect 271196 136632 272524 136660
rect 271196 136620 271202 136632
rect 272518 136620 272524 136632
rect 272576 136620 272582 136672
rect 73062 87320 73068 87372
rect 73120 87360 73126 87372
rect 345658 87360 345664 87372
rect 73120 87332 345664 87360
rect 73120 87320 73126 87332
rect 345658 87320 345664 87332
rect 345716 87320 345722 87372
rect 74442 87252 74448 87304
rect 74500 87292 74506 87304
rect 86310 87292 86316 87304
rect 74500 87264 86316 87292
rect 74500 87252 74506 87264
rect 86310 87252 86316 87264
rect 86368 87252 86374 87304
rect 66990 87184 66996 87236
rect 67048 87224 67054 87236
rect 84930 87224 84936 87236
rect 67048 87196 84936 87224
rect 67048 87184 67054 87196
rect 84930 87184 84936 87196
rect 84988 87184 84994 87236
rect 70118 87116 70124 87168
rect 70176 87156 70182 87168
rect 98730 87156 98736 87168
rect 70176 87128 98736 87156
rect 70176 87116 70182 87128
rect 98730 87116 98736 87128
rect 98788 87116 98794 87168
rect 76466 87048 76472 87100
rect 76524 87088 76530 87100
rect 287698 87088 287704 87100
rect 76524 87060 287704 87088
rect 76524 87048 76530 87060
rect 287698 87048 287704 87060
rect 287756 87048 287762 87100
rect 82722 86980 82728 87032
rect 82780 87020 82786 87032
rect 90450 87020 90456 87032
rect 82780 86992 90456 87020
rect 82780 86980 82786 86992
rect 90450 86980 90456 86992
rect 90508 86980 90514 87032
rect 84930 83444 84936 83496
rect 84988 83484 84994 83496
rect 336274 83484 336280 83496
rect 84988 83456 336280 83484
rect 84988 83444 84994 83456
rect 336274 83444 336280 83456
rect 336332 83444 336338 83496
rect 84194 82764 84200 82816
rect 84252 82804 84258 82816
rect 295978 82804 295984 82816
rect 84252 82776 295984 82804
rect 84252 82764 84258 82776
rect 295978 82764 295984 82776
rect 296036 82764 296042 82816
rect 86310 69640 86316 69692
rect 86368 69680 86374 69692
rect 350442 69680 350448 69692
rect 86368 69652 350448 69680
rect 86368 69640 86374 69652
rect 350442 69640 350448 69652
rect 350500 69640 350506 69692
rect 88242 51688 88248 51740
rect 88300 51728 88306 51740
rect 110414 51728 110420 51740
rect 88300 51700 110420 51728
rect 88300 51688 88306 51700
rect 110414 51688 110420 51700
rect 110472 51688 110478 51740
rect 90450 50328 90456 50380
rect 90508 50368 90514 50380
rect 368198 50368 368204 50380
rect 90508 50340 368204 50368
rect 90508 50328 90514 50340
rect 368198 50328 368204 50340
rect 368256 50328 368262 50380
rect 566 40672 572 40724
rect 624 40712 630 40724
rect 86954 40712 86960 40724
rect 624 40684 86960 40712
rect 624 40672 630 40684
rect 86954 40672 86960 40684
rect 87012 40672 87018 40724
rect 98730 10276 98736 10328
rect 98788 10316 98794 10328
rect 339862 10316 339868 10328
rect 98788 10288 339868 10316
rect 98788 10276 98794 10288
rect 339862 10276 339868 10288
rect 339920 10276 339926 10328
rect 291838 6808 291844 6860
rect 291896 6848 291902 6860
rect 580166 6848 580172 6860
rect 291896 6820 580172 6848
rect 291896 6808 291902 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 287698 4768 287704 4820
rect 287756 4808 287762 4820
rect 354030 4808 354036 4820
rect 287756 4780 354036 4808
rect 287756 4768 287762 4780
rect 354030 4768 354036 4780
rect 354088 4768 354094 4820
rect 345658 4156 345664 4208
rect 345716 4196 345722 4208
rect 346946 4196 346952 4208
rect 345716 4168 346952 4196
rect 345716 4156 345722 4168
rect 346946 4156 346952 4168
rect 347004 4156 347010 4208
rect 241422 4088 241428 4140
rect 241480 4128 241486 4140
rect 282914 4128 282920 4140
rect 241480 4100 282920 4128
rect 241480 4088 241486 4100
rect 282914 4088 282920 4100
rect 282972 4088 282978 4140
rect 264974 4020 264980 4072
rect 265032 4060 265038 4072
rect 291746 4060 291752 4072
rect 265032 4032 291752 4060
rect 265032 4020 265038 4032
rect 291746 4020 291752 4032
rect 291804 4020 291810 4072
rect 295978 3408 295984 3460
rect 296036 3448 296042 3460
rect 371694 3448 371700 3460
rect 296036 3420 371700 3448
rect 296036 3408 296042 3420
rect 371694 3408 371700 3420
rect 371752 3408 371758 3460
rect 442258 3408 442264 3460
rect 442316 3448 442322 3460
rect 583386 3448 583392 3460
rect 442316 3420 583392 3448
rect 442316 3408 442322 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 438854 2796 438860 2848
rect 438912 2836 438918 2848
rect 580994 2836 581000 2848
rect 438912 2808 581000 2836
rect 438912 2796 438918 2808
rect 580994 2796 581000 2808
rect 581052 2796 581058 2848
<< via1 >>
rect 40500 700952 40552 701004
rect 59268 700952 59320 701004
rect 105452 700272 105504 700324
rect 137284 700272 137336 700324
rect 257344 700272 257396 700324
rect 267648 700272 267700 700324
rect 348792 700272 348844 700324
rect 365628 700272 365680 700324
rect 527180 700272 527232 700324
rect 546500 700272 546552 700324
rect 365628 695444 365680 695496
rect 371884 695444 371936 695496
rect 332508 694764 332560 694816
rect 338764 694764 338816 694816
rect 247684 687896 247736 687948
rect 257344 687896 257396 687948
rect 3424 683136 3476 683188
rect 55220 683136 55272 683188
rect 144184 683136 144236 683188
rect 338764 682388 338816 682440
rect 358728 682388 358780 682440
rect 358728 680280 358780 680332
rect 366364 680280 366416 680332
rect 244556 676132 244608 676184
rect 247684 676132 247736 676184
rect 507124 670692 507176 670744
rect 580172 670692 580224 670744
rect 232504 668584 232556 668636
rect 244556 668584 244608 668636
rect 371884 664436 371936 664488
rect 377404 664436 377456 664488
rect 366364 663008 366416 663060
rect 382280 663008 382332 663060
rect 382280 660288 382332 660340
rect 388444 660288 388496 660340
rect 137284 658180 137336 658232
rect 138020 658180 138072 658232
rect 170312 658180 170364 658232
rect 171140 658180 171192 658232
rect 172428 658180 172480 658232
rect 388444 658180 388496 658232
rect 393964 658180 394016 658232
rect 429844 657704 429896 657756
rect 478880 657704 478932 657756
rect 485596 657704 485648 657756
rect 494796 657704 494848 657756
rect 510068 657704 510120 657756
rect 298744 657636 298796 657688
rect 364984 657636 365036 657688
rect 512828 657636 512880 657688
rect 144184 657568 144236 657620
rect 521108 657568 521160 657620
rect 141424 657500 141476 657552
rect 519728 657500 519780 657552
rect 138020 657228 138072 657280
rect 518348 657228 518400 657280
rect 485688 657160 485740 657212
rect 507124 657160 507176 657212
rect 478880 657092 478932 657144
rect 480168 657092 480220 657144
rect 511448 657092 511500 657144
rect 172428 657024 172480 657076
rect 516968 657024 517020 657076
rect 528008 657024 528060 657076
rect 543832 657024 543884 657076
rect 162124 656956 162176 657008
rect 526628 656956 526680 657008
rect 533528 656956 533580 657008
rect 547880 656956 547932 657008
rect 487068 656888 487120 656940
rect 499028 656888 499080 656940
rect 539048 656888 539100 656940
rect 547972 656888 548024 656940
rect 505928 655664 505980 655716
rect 540336 655664 540388 655716
rect 155224 655596 155276 655648
rect 525248 655596 525300 655648
rect 148324 655528 148376 655580
rect 522488 655528 522540 655580
rect 151084 654440 151136 654492
rect 523500 654440 523552 654492
rect 159364 648592 159416 648644
rect 361948 648592 362000 648644
rect 393964 648524 394016 648576
rect 397368 648524 397420 648576
rect 204904 647436 204956 647488
rect 358084 647436 358136 647488
rect 202788 647368 202840 647420
rect 359372 647368 359424 647420
rect 233148 647300 233200 647352
rect 471244 647300 471296 647352
rect 208400 647232 208452 647284
rect 468484 647232 468536 647284
rect 222844 646484 222896 646536
rect 232504 646484 232556 646536
rect 212448 646008 212500 646060
rect 354220 646008 354272 646060
rect 186596 645940 186648 645992
rect 461768 645940 461820 645992
rect 194324 645872 194376 645924
rect 471336 645872 471388 645924
rect 215300 644920 215352 644972
rect 324596 644920 324648 644972
rect 231768 644852 231820 644904
rect 375472 644852 375524 644904
rect 106188 644784 106240 644836
rect 352932 644784 352984 644836
rect 227720 644716 227772 644768
rect 480352 644716 480404 644768
rect 102140 644648 102192 644700
rect 355508 644648 355560 644700
rect 397368 644648 397420 644700
rect 404360 644648 404412 644700
rect 191748 644580 191800 644632
rect 489368 644580 489420 644632
rect 189172 644512 189224 644564
rect 488080 644512 488132 644564
rect 187884 644444 187936 644496
rect 490104 644444 490156 644496
rect 377404 643696 377456 643748
rect 397460 643696 397512 643748
rect 176660 643560 176712 643612
rect 356796 643560 356848 643612
rect 233884 643492 233936 643544
rect 486700 643492 486752 643544
rect 207020 643424 207072 643476
rect 467196 643424 467248 643476
rect 88984 643356 89036 643408
rect 364524 643356 364576 643408
rect 86868 643288 86920 643340
rect 365812 643288 365864 643340
rect 80060 643220 80112 643272
rect 367100 643220 367152 643272
rect 204168 643152 204220 643204
rect 489920 643152 489972 643204
rect 179328 643084 179380 643136
rect 474004 643084 474056 643136
rect 223488 642200 223540 642252
rect 328460 642200 328512 642252
rect 92480 642132 92532 642184
rect 342628 642132 342680 642184
rect 85488 642064 85540 642116
rect 349068 642064 349120 642116
rect 179328 641996 179380 642048
rect 474096 641996 474148 642048
rect 177948 641928 178000 641980
rect 479432 641928 479484 641980
rect 177764 641860 177816 641912
rect 488540 641860 488592 641912
rect 177856 641792 177908 641844
rect 490012 641792 490064 641844
rect 249708 641724 249760 641776
rect 369676 641724 369728 641776
rect 218060 640840 218112 640892
rect 315580 640840 315632 640892
rect 214564 640772 214616 640824
rect 320732 640772 320784 640824
rect 91100 640704 91152 640756
rect 329748 640704 329800 640756
rect 230388 640636 230440 640688
rect 485872 640636 485924 640688
rect 216772 640568 216824 640620
rect 480444 640568 480496 640620
rect 211068 640500 211120 640552
rect 488816 640500 488868 640552
rect 185676 640432 185728 640484
rect 464436 640432 464488 640484
rect 190736 640364 190788 640416
rect 490196 640364 490248 640416
rect 56508 640296 56560 640348
rect 363236 640296 363288 640348
rect 404360 640296 404412 640348
rect 410524 640296 410576 640348
rect 397460 640228 397512 640280
rect 400864 640228 400916 640280
rect 220728 639548 220780 639600
rect 485780 639548 485832 639600
rect 122748 639412 122800 639464
rect 306564 639412 306616 639464
rect 95148 639344 95200 639396
rect 318156 639344 318208 639396
rect 251088 639276 251140 639328
rect 479340 639276 479392 639328
rect 82820 639208 82872 639260
rect 319444 639208 319496 639260
rect 81440 639140 81492 639192
rect 322020 639140 322072 639192
rect 125600 639072 125652 639124
rect 376852 639072 376904 639124
rect 234620 639004 234672 639056
rect 487252 639004 487304 639056
rect 58624 638936 58676 638988
rect 139032 638936 139084 638988
rect 213828 638936 213880 638988
rect 488632 638936 488684 638988
rect 129740 638392 129792 638444
rect 283748 638392 283800 638444
rect 123484 638324 123536 638376
rect 289084 638324 289136 638376
rect 278136 638256 278188 638308
rect 343916 638256 343968 638308
rect 211068 638188 211120 638240
rect 487160 638188 487212 638240
rect 280896 638120 280948 638172
rect 346492 638120 346544 638172
rect 283564 638052 283616 638104
rect 347780 638052 347832 638104
rect 110328 637984 110380 638036
rect 295984 637984 296036 638036
rect 108304 637916 108356 637968
rect 331036 637916 331088 637968
rect 247500 637848 247552 637900
rect 488540 637848 488592 637900
rect 224224 637780 224276 637832
rect 480260 637780 480312 637832
rect 230388 637712 230440 637764
rect 487436 637712 487488 637764
rect 115480 637644 115532 637696
rect 381544 637644 381596 637696
rect 109040 637576 109092 637628
rect 375564 637576 375616 637628
rect 73160 637032 73212 637084
rect 350356 637032 350408 637084
rect 241060 636964 241112 637016
rect 468576 636964 468628 637016
rect 273996 636896 274048 636948
rect 302700 636896 302752 636948
rect 101312 636828 101364 636880
rect 135996 636828 136048 636880
rect 249616 636828 249668 636880
rect 268384 636828 268436 636880
rect 279700 636828 279752 636880
rect 314292 636828 314344 636880
rect 124220 636760 124272 636812
rect 135904 636760 135956 636812
rect 238392 636760 238444 636812
rect 271236 636760 271288 636812
rect 275376 636760 275428 636812
rect 327172 636760 327224 636812
rect 99380 636692 99432 636744
rect 311716 636692 311768 636744
rect 114192 636624 114244 636676
rect 138664 636624 138716 636676
rect 243636 636624 243688 636676
rect 465816 636624 465868 636676
rect 111616 636556 111668 636608
rect 138756 636556 138808 636608
rect 239680 636556 239732 636608
rect 468668 636556 468720 636608
rect 106464 636488 106516 636540
rect 162308 636488 162360 636540
rect 237104 636488 237156 636540
rect 468760 636488 468812 636540
rect 78588 636420 78640 636472
rect 323308 636420 323360 636472
rect 75828 636352 75880 636404
rect 338764 636352 338816 636404
rect 131120 636284 131172 636336
rect 134708 636284 134760 636336
rect 129648 636216 129700 636268
rect 249708 636216 249760 636268
rect 369676 636216 369728 636268
rect 374552 636216 374604 636268
rect 79324 635672 79376 635724
rect 296720 635672 296772 635724
rect 53840 635604 53892 635656
rect 377036 635604 377088 635656
rect 170404 635536 170456 635588
rect 222844 635536 222896 635588
rect 271144 635536 271196 635588
rect 325884 635536 325936 635588
rect 39948 635468 40000 635520
rect 72976 635468 73028 635520
rect 112904 635468 112956 635520
rect 264244 635468 264296 635520
rect 276848 635468 276900 635520
rect 337476 635468 337528 635520
rect 119988 635400 120040 635452
rect 273904 635400 273956 635452
rect 274088 635400 274140 635452
rect 372252 635400 372304 635452
rect 121368 635332 121420 635384
rect 290464 635332 290516 635384
rect 97908 635264 97960 635316
rect 297548 635264 297600 635316
rect 252468 635196 252520 635248
rect 465724 635196 465776 635248
rect 289176 635128 289228 635180
rect 341340 635128 341392 635180
rect 244280 635060 244332 635112
rect 487344 635060 487396 635112
rect 226340 634992 226392 635044
rect 476764 634992 476816 635044
rect 71872 634924 71924 634976
rect 377220 634924 377272 634976
rect 70584 634856 70636 634908
rect 377128 634856 377180 634908
rect 246120 634788 246172 634840
rect 265624 634788 265676 634840
rect 286416 634584 286468 634636
rect 312636 634584 312688 634636
rect 284944 634516 284996 634568
rect 307668 634516 307720 634568
rect 274180 634448 274232 634500
rect 316500 634448 316552 634500
rect 129832 634380 129884 634432
rect 297180 634380 297232 634432
rect 139032 633360 139084 633412
rect 148324 633360 148376 633412
rect 3424 632680 3476 632732
rect 55588 632680 55640 632732
rect 374552 632680 374604 632732
rect 453304 632680 453356 632732
rect 410524 632000 410576 632052
rect 413284 632000 413336 632052
rect 377680 625540 377732 625592
rect 380992 625540 381044 625592
rect 377680 623772 377732 623824
rect 381084 623772 381136 623824
rect 164976 622412 165028 622464
rect 170404 622412 170456 622464
rect 377772 622412 377824 622464
rect 381176 622412 381228 622464
rect 377036 620984 377088 621036
rect 379520 620984 379572 621036
rect 400864 617516 400916 617568
rect 426348 617516 426400 617568
rect 540336 617516 540388 617568
rect 580172 617516 580224 617568
rect 283656 614116 283708 614168
rect 298008 614116 298060 614168
rect 453304 613368 453356 613420
rect 477500 613368 477552 613420
rect 413284 612756 413336 612808
rect 416044 612756 416096 612808
rect 477500 612756 477552 612808
rect 478788 612756 478840 612808
rect 487160 612756 487212 612808
rect 159548 612008 159600 612060
rect 164976 612008 165028 612060
rect 289360 611328 289412 611380
rect 298008 611328 298060 611380
rect 283840 609968 283892 610020
rect 298008 609968 298060 610020
rect 426348 609220 426400 609272
rect 442264 609220 442316 609272
rect 378048 605820 378100 605872
rect 385040 605820 385092 605872
rect 378048 604528 378100 604580
rect 386420 604528 386472 604580
rect 377956 604460 378008 604512
rect 389180 604460 389232 604512
rect 378048 603236 378100 603288
rect 385132 603236 385184 603288
rect 378048 603100 378100 603152
rect 386604 603100 386656 603152
rect 538588 600584 538640 600636
rect 539324 600584 539376 600636
rect 535736 600244 535788 600296
rect 542636 600244 542688 600296
rect 536840 600176 536892 600228
rect 542728 600176 542780 600228
rect 534724 600108 534776 600160
rect 540336 600108 540388 600160
rect 487068 599700 487120 599752
rect 498200 599700 498252 599752
rect 485596 599632 485648 599684
rect 505100 599632 505152 599684
rect 485688 599564 485740 599616
rect 506480 599564 506532 599616
rect 502984 598204 503036 598256
rect 539048 598204 539100 598256
rect 157064 597456 157116 597508
rect 159548 597456 159600 597508
rect 47952 594804 48004 594856
rect 56968 594804 57020 594856
rect 285312 594804 285364 594856
rect 298008 594804 298060 594856
rect 378048 594804 378100 594856
rect 385224 594804 385276 594856
rect 442264 594804 442316 594856
rect 448520 594804 448572 594856
rect 147404 594056 147456 594108
rect 157064 594056 157116 594108
rect 378048 592084 378100 592136
rect 383660 592084 383712 592136
rect 377956 592016 378008 592068
rect 386696 592016 386748 592068
rect 448520 591268 448572 591320
rect 454684 591268 454736 591320
rect 50620 590656 50672 590708
rect 56968 590656 57020 590708
rect 144276 590656 144328 590708
rect 147404 590656 147456 590708
rect 288164 590656 288216 590708
rect 298008 590656 298060 590708
rect 378048 590656 378100 590708
rect 385408 590656 385460 590708
rect 378048 589636 378100 589688
rect 385316 589636 385368 589688
rect 53380 589500 53432 589552
rect 56968 589500 57020 589552
rect 378048 587936 378100 587988
rect 382648 587936 382700 587988
rect 377036 587868 377088 587920
rect 379796 587868 379848 587920
rect 377864 587052 377916 587104
rect 381452 587052 381504 587104
rect 377864 586644 377916 586696
rect 381360 586644 381412 586696
rect 377220 585216 377272 585268
rect 379980 585216 380032 585268
rect 137560 585148 137612 585200
rect 144276 585148 144328 585200
rect 377036 585148 377088 585200
rect 379704 585148 379756 585200
rect 416044 584740 416096 584792
rect 423588 584740 423640 584792
rect 377772 583720 377824 583772
rect 381268 583720 381320 583772
rect 378048 582768 378100 582820
rect 382372 582768 382424 582820
rect 378048 582428 378100 582480
rect 383936 582428 383988 582480
rect 378048 581000 378100 581052
rect 383752 581000 383804 581052
rect 423588 580252 423640 580304
rect 432604 580252 432656 580304
rect 3424 579640 3476 579692
rect 47584 579640 47636 579692
rect 378048 579640 378100 579692
rect 382464 579640 382516 579692
rect 378048 578280 378100 578332
rect 382556 578280 382608 578332
rect 377036 578212 377088 578264
rect 379888 578212 379940 578264
rect 134708 575492 134760 575544
rect 137560 575492 137612 575544
rect 454684 574744 454736 574796
rect 475384 574744 475436 574796
rect 378048 574064 378100 574116
rect 386788 574064 386840 574116
rect 377588 572704 377640 572756
rect 380900 572704 380952 572756
rect 166632 569780 166684 569832
rect 172244 569780 172296 569832
rect 377956 568556 378008 568608
rect 381636 568556 381688 568608
rect 285036 567196 285088 567248
rect 296720 567196 296772 567248
rect 56968 563184 57020 563236
rect 57520 563184 57572 563236
rect 291936 560872 291988 560924
rect 298008 560872 298060 560924
rect 98736 560600 98788 560652
rect 160836 560600 160888 560652
rect 178592 560600 178644 560652
rect 288164 560600 288216 560652
rect 179420 560532 179472 560584
rect 285312 560532 285364 560584
rect 179236 560328 179288 560380
rect 179512 560328 179564 560380
rect 57336 560260 57388 560312
rect 58072 560260 58124 560312
rect 299756 560260 299808 560312
rect 309784 560260 309836 560312
rect 57612 560192 57664 560244
rect 376116 560192 376168 560244
rect 57336 560124 57388 560176
rect 297824 560124 297876 560176
rect 57520 560056 57572 560108
rect 297640 560056 297692 560108
rect 169392 559988 169444 560040
rect 173072 559988 173124 560040
rect 166816 559920 166868 559972
rect 173808 559920 173860 559972
rect 372068 559852 372120 559904
rect 379980 559852 380032 559904
rect 371884 559784 371936 559836
rect 379796 559784 379848 559836
rect 371976 559716 372028 559768
rect 381268 559716 381320 559768
rect 372160 559648 372212 559700
rect 381452 559648 381504 559700
rect 90916 559580 90968 559632
rect 139584 559580 139636 559632
rect 268384 559580 268436 559632
rect 514760 559580 514812 559632
rect 76012 559512 76064 559564
rect 135168 559512 135220 559564
rect 177212 559512 177264 559564
rect 487160 559512 487212 559564
rect 63776 558900 63828 558952
rect 68284 558900 68336 558952
rect 97816 558900 97868 558952
rect 254584 558900 254636 558952
rect 57612 558832 57664 558884
rect 381360 558832 381412 558884
rect 56508 558764 56560 558816
rect 361212 558764 361264 558816
rect 47952 558696 48004 558748
rect 98736 558696 98788 558748
rect 109132 558696 109184 558748
rect 289360 558696 289412 558748
rect 120080 558628 120132 558680
rect 163872 558628 163924 558680
rect 279792 558424 279844 558476
rect 506664 558424 506716 558476
rect 60464 558356 60516 558408
rect 297548 558356 297600 558408
rect 60556 558288 60608 558340
rect 298744 558288 298796 558340
rect 271236 558220 271288 558272
rect 512000 558220 512052 558272
rect 59636 558152 59688 558204
rect 360200 558152 360252 558204
rect 372620 558152 372672 558204
rect 377128 558152 377180 558204
rect 117964 557676 118016 557728
rect 216128 557676 216180 557728
rect 120172 557608 120224 557660
rect 253296 557608 253348 557660
rect 280160 557608 280212 557660
rect 492772 557608 492824 557660
rect 117780 557540 117832 557592
rect 259828 557540 259880 557592
rect 284208 557540 284260 557592
rect 509424 557540 509476 557592
rect 56508 557472 56560 557524
rect 379704 557472 379756 557524
rect 55864 557404 55916 557456
rect 377036 557404 377088 557456
rect 60096 557336 60148 557388
rect 376024 557336 376076 557388
rect 95148 557268 95200 557320
rect 297916 557268 297968 557320
rect 265624 556860 265676 556912
rect 512092 556860 512144 556912
rect 50620 556792 50672 556844
rect 92388 556792 92440 556844
rect 163780 556792 163832 556844
rect 175096 556792 175148 556844
rect 424048 556792 424100 556844
rect 86960 556180 87012 556232
rect 90916 556180 90968 556232
rect 178040 556180 178092 556232
rect 422484 556180 422536 556232
rect 100760 556112 100812 556164
rect 378692 556112 378744 556164
rect 121460 556044 121512 556096
rect 339960 556044 340012 556096
rect 332600 555568 332652 555620
rect 372620 555568 372672 555620
rect 137284 555500 137336 555552
rect 360844 555500 360896 555552
rect 57152 555432 57204 555484
rect 375932 555432 375984 555484
rect 57704 555160 57756 555212
rect 57704 554956 57756 555008
rect 58624 554752 58676 554804
rect 124128 554752 124180 554804
rect 262956 554752 263008 554804
rect 275928 554752 275980 554804
rect 492864 554752 492916 554804
rect 73160 554684 73212 554736
rect 350080 554684 350132 554736
rect 88984 554616 89036 554668
rect 310612 554616 310664 554668
rect 58624 554548 58676 554600
rect 107568 554548 107620 554600
rect 297456 554548 297508 554600
rect 136088 554004 136140 554056
rect 320824 554004 320876 554056
rect 115848 553460 115900 553512
rect 247316 553460 247368 553512
rect 299296 553460 299348 553512
rect 489092 553460 489144 553512
rect 108304 553392 108356 553444
rect 258264 553392 258316 553444
rect 293960 553392 294012 553444
rect 493048 553392 493100 553444
rect 81440 553324 81492 553376
rect 347044 553324 347096 553376
rect 57796 553256 57848 553308
rect 286416 553256 286468 553308
rect 299296 553256 299348 553308
rect 303528 553256 303580 553308
rect 98644 553188 98696 553240
rect 305552 553188 305604 553240
rect 179420 553120 179472 553172
rect 297732 553120 297784 553172
rect 47584 552644 47636 552696
rect 60556 552644 60608 552696
rect 151084 552644 151136 552696
rect 304264 552644 304316 552696
rect 332600 552644 332652 552696
rect 173808 552372 173860 552424
rect 509332 552372 509384 552424
rect 295340 552304 295392 552356
rect 358360 552304 358412 552356
rect 291752 552236 291804 552288
rect 439688 552236 439740 552288
rect 278688 552168 278740 552220
rect 491300 552168 491352 552220
rect 175832 552100 175884 552152
rect 502524 552100 502576 552152
rect 58716 552032 58768 552084
rect 169760 552032 169812 552084
rect 52460 551964 52512 552016
rect 356152 551964 356204 552016
rect 59268 551896 59320 551948
rect 348056 551896 348108 551948
rect 99380 551828 99432 551880
rect 379888 551828 379940 551880
rect 81440 551760 81492 551812
rect 328828 551760 328880 551812
rect 124864 551352 124916 551404
rect 134708 551352 134760 551404
rect 60096 551284 60148 551336
rect 359188 551284 359240 551336
rect 269120 550740 269172 550792
rect 469404 550740 469456 550792
rect 241428 550672 241480 550724
rect 492956 550672 493008 550724
rect 178040 550604 178092 550656
rect 497464 550604 497516 550656
rect 85488 550536 85540 550588
rect 365260 550536 365312 550588
rect 100760 550468 100812 550520
rect 353116 550468 353168 550520
rect 179420 550400 179472 550452
rect 380900 550400 380952 550452
rect 169760 550332 169812 550384
rect 326804 550332 326856 550384
rect 233148 550264 233200 550316
rect 283840 550264 283892 550316
rect 273904 550060 273956 550112
rect 352104 550060 352156 550112
rect 283748 549992 283800 550044
rect 364616 549992 364668 550044
rect 134616 549924 134668 549976
rect 328644 549924 328696 549976
rect 177304 549856 177356 549908
rect 491668 549856 491720 549908
rect 71044 549244 71096 549296
rect 75828 549244 75880 549296
rect 81808 549244 81860 549296
rect 86868 549448 86920 549500
rect 224960 549244 225012 549296
rect 260794 549244 260846 549296
rect 260932 549244 260984 549296
rect 487620 549244 487672 549296
rect 86868 549176 86920 549228
rect 342996 549176 343048 549228
rect 75828 549108 75880 549160
rect 260840 549108 260892 549160
rect 126888 549040 126940 549092
rect 280068 549108 280120 549160
rect 313648 549108 313700 549160
rect 322756 549040 322808 549092
rect 59268 548972 59320 549024
rect 159364 548972 159416 549024
rect 260932 548972 260984 549024
rect 279700 548972 279752 549024
rect 162308 548632 162360 548684
rect 363052 548632 363104 548684
rect 432604 548632 432656 548684
rect 443644 548632 443696 548684
rect 202788 548564 202840 548616
rect 502340 548564 502392 548616
rect 177120 548496 177172 548548
rect 493140 548496 493192 548548
rect 58716 548292 58768 548344
rect 59268 548292 59320 548344
rect 278688 547884 278740 547936
rect 514852 547884 514904 547936
rect 78588 547816 78640 547868
rect 375656 547816 375708 547868
rect 89720 547748 89772 547800
rect 346032 547748 346084 547800
rect 126888 547680 126940 547732
rect 320732 547680 320784 547732
rect 216680 547612 216732 547664
rect 306564 547612 306616 547664
rect 135996 547272 136048 547324
rect 356796 547272 356848 547324
rect 226064 547204 226116 547256
rect 486148 547204 486200 547256
rect 188620 547136 188672 547188
rect 495440 547136 495492 547188
rect 230388 546524 230440 546576
rect 305184 546524 305236 546576
rect 173808 546456 173860 546508
rect 456892 546456 456944 546508
rect 60188 546388 60240 546440
rect 372344 546388 372396 546440
rect 189632 546320 189684 546372
rect 485780 546320 485832 546372
rect 79324 546252 79376 546304
rect 362224 546252 362276 546304
rect 121460 546184 121512 546236
rect 323768 546184 323820 546236
rect 89720 546116 89772 546168
rect 284944 546116 284996 546168
rect 223488 546048 223540 546100
rect 382648 546048 382700 546100
rect 207848 545708 207900 545760
rect 503996 545708 504048 545760
rect 75828 545164 75880 545216
rect 81808 545164 81860 545216
rect 92480 545028 92532 545080
rect 381176 545028 381228 545080
rect 127624 544960 127676 545012
rect 371332 544960 371384 545012
rect 153108 544892 153160 544944
rect 308588 544892 308640 544944
rect 172428 544824 172480 544876
rect 302516 544824 302568 544876
rect 215944 544416 215996 544468
rect 494244 544416 494296 544468
rect 199752 544348 199804 544400
rect 480536 544348 480588 544400
rect 293960 543804 294012 543856
rect 348976 543804 349028 543856
rect 72424 543668 72476 543720
rect 75828 543736 75880 543788
rect 175280 543736 175332 543788
rect 436560 543736 436612 543788
rect 95148 543668 95200 543720
rect 345020 543668 345072 543720
rect 125508 543600 125560 543652
rect 318708 543600 318760 543652
rect 175280 543532 175332 543584
rect 307576 543532 307628 543584
rect 283748 543124 283800 543176
rect 357164 543124 357216 543176
rect 138756 543056 138808 543108
rect 369216 543056 369268 543108
rect 177396 542988 177448 543040
rect 494428 542988 494480 543040
rect 230388 542444 230440 542496
rect 497004 542444 497056 542496
rect 172520 542376 172572 542428
rect 466276 542376 466328 542428
rect 111800 542308 111852 542360
rect 364248 542308 364300 542360
rect 224224 542240 224276 542292
rect 386788 542240 386840 542292
rect 172520 542172 172572 542224
rect 314660 542172 314712 542224
rect 135904 541832 135956 541884
rect 355232 541832 355284 541884
rect 196716 541764 196768 541816
rect 480628 541764 480680 541816
rect 187608 541696 187660 541748
rect 496912 541696 496964 541748
rect 182548 541628 182600 541680
rect 495532 541628 495584 541680
rect 233148 540948 233200 541000
rect 494336 540948 494388 541000
rect 91100 540880 91152 540932
rect 352012 540880 352064 540932
rect 121460 540812 121512 540864
rect 349068 540812 349120 540864
rect 75828 540744 75880 540796
rect 276848 540744 276900 540796
rect 272524 540676 272576 540728
rect 317696 540676 317748 540728
rect 443644 540472 443696 540524
rect 453304 540472 453356 540524
rect 208860 540404 208912 540456
rect 487804 540404 487856 540456
rect 169024 540336 169076 540388
rect 470968 540336 471020 540388
rect 177488 540268 177540 540320
rect 493232 540268 493284 540320
rect 183560 540200 183612 540252
rect 503904 540200 503956 540252
rect 86868 539520 86920 539572
rect 373356 539520 373408 539572
rect 118700 539452 118752 539504
rect 332876 539452 332928 539504
rect 131120 539384 131172 539436
rect 316684 539384 316736 539436
rect 298744 539316 298796 539368
rect 304264 539316 304316 539368
rect 138664 538976 138716 539028
rect 372436 538976 372488 539028
rect 209872 538908 209924 538960
rect 486056 538908 486108 538960
rect 194692 538840 194744 538892
rect 480720 538840 480772 538892
rect 256700 538296 256752 538348
rect 491484 538296 491536 538348
rect 171968 538228 172020 538280
rect 447508 538228 447560 538280
rect 60832 538160 60884 538212
rect 381084 538160 381136 538212
rect 82820 538092 82872 538144
rect 370320 538092 370372 538144
rect 124128 538024 124180 538076
rect 367284 538024 367336 538076
rect 171784 537956 171836 538008
rect 331864 537956 331916 538008
rect 291844 537888 291896 537940
rect 381636 537888 381688 537940
rect 252468 537820 252520 537872
rect 315672 537820 315724 537872
rect 203800 537548 203852 537600
rect 480996 537548 481048 537600
rect 195796 537480 195848 537532
rect 480812 537480 480864 537532
rect 171048 536800 171100 536852
rect 508136 536800 508188 536852
rect 97908 536732 97960 536784
rect 344008 536732 344060 536784
rect 128360 536664 128412 536716
rect 341984 536664 342036 536716
rect 178040 536596 178092 536648
rect 330852 536596 330904 536648
rect 292580 536528 292632 536580
rect 311624 536528 311676 536580
rect 179604 536052 179656 536104
rect 506756 536052 506808 536104
rect 218060 535576 218112 535628
rect 487896 535576 487948 535628
rect 173992 535508 174044 535560
rect 463148 535508 463200 535560
rect 205640 535440 205692 535492
rect 501144 535440 501196 535492
rect 97908 535372 97960 535424
rect 358176 535372 358228 535424
rect 155868 535304 155920 535356
rect 321744 535304 321796 535356
rect 179236 534760 179288 534812
rect 461492 534760 461544 534812
rect 175188 534692 175240 534744
rect 464712 534692 464764 534744
rect 243544 534284 243596 534336
rect 487988 534284 488040 534336
rect 164148 534216 164200 534268
rect 427084 534216 427136 534268
rect 212448 534148 212500 534200
rect 480904 534148 480956 534200
rect 70492 534080 70544 534132
rect 72424 534080 72476 534132
rect 194508 534080 194560 534132
rect 500960 534080 501012 534132
rect 60740 534012 60792 534064
rect 369308 534012 369360 534064
rect 70400 533944 70452 533996
rect 354128 533944 354180 533996
rect 59176 533876 59228 533928
rect 280896 533876 280948 533928
rect 167000 533808 167052 533860
rect 338948 533808 339000 533860
rect 175832 533740 175884 533792
rect 327816 533740 327868 533792
rect 177580 533400 177632 533452
rect 491760 533332 491812 533384
rect 67916 532788 67968 532840
rect 71044 532788 71096 532840
rect 244372 532788 244424 532840
rect 502432 532788 502484 532840
rect 191748 532720 191800 532772
rect 493508 532720 493560 532772
rect 96528 532652 96580 532704
rect 368296 532652 368348 532704
rect 117228 532584 117280 532636
rect 340972 532584 341024 532636
rect 131120 532516 131172 532568
rect 329840 532516 329892 532568
rect 178040 532448 178092 532500
rect 285036 532448 285088 532500
rect 290464 532176 290516 532228
rect 330208 532176 330260 532228
rect 178868 532108 178920 532160
rect 403716 532108 403768 532160
rect 178684 532040 178736 532092
rect 450636 532040 450688 532092
rect 174636 531972 174688 532024
rect 455328 531972 455380 532024
rect 213828 531292 213880 531344
rect 494152 531292 494204 531344
rect 59912 531224 59964 531276
rect 366272 531224 366324 531276
rect 67548 531156 67600 531208
rect 355140 531156 355192 531208
rect 111800 531088 111852 531140
rect 335912 531088 335964 531140
rect 59176 531020 59228 531072
rect 278136 531020 278188 531072
rect 211068 530952 211120 531004
rect 337936 530952 337988 531004
rect 64788 530544 64840 530596
rect 67916 530544 67968 530596
rect 113180 530544 113232 530596
rect 124864 530544 124916 530596
rect 177672 530544 177724 530596
rect 489276 530544 489328 530596
rect 295340 530068 295392 530120
rect 497188 530068 497240 530120
rect 289728 530000 289780 530052
rect 497096 530000 497148 530052
rect 251088 529932 251140 529984
rect 479616 529932 479668 529984
rect 59452 529864 59504 529916
rect 378232 529864 378284 529916
rect 59176 529796 59228 529848
rect 363236 529796 363288 529848
rect 68652 529728 68704 529780
rect 70308 529728 70360 529780
rect 127624 529728 127676 529780
rect 375380 529728 375432 529780
rect 135168 529660 135220 529712
rect 378324 529660 378376 529712
rect 166264 529592 166316 529644
rect 374552 529592 374604 529644
rect 181536 529184 181588 529236
rect 501052 529184 501104 529236
rect 289728 528640 289780 528692
rect 499856 528640 499908 528692
rect 177488 528572 177540 528624
rect 493324 528572 493376 528624
rect 175832 528504 175884 528556
rect 378416 528504 378468 528556
rect 175188 528436 175240 528488
rect 374736 528436 374788 528488
rect 220636 528368 220688 528420
rect 378600 528368 378652 528420
rect 279976 528300 280028 528352
rect 375840 528300 375892 528352
rect 92480 527892 92532 527944
rect 113180 527892 113232 527944
rect 60372 527824 60424 527876
rect 155224 527824 155276 527876
rect 186596 527824 186648 527876
rect 498292 527824 498344 527876
rect 286324 527212 286376 527264
rect 497280 527212 497332 527264
rect 3424 527144 3476 527196
rect 60372 527144 60424 527196
rect 62212 527144 62264 527196
rect 64788 527144 64840 527196
rect 66168 527144 66220 527196
rect 68652 527144 68704 527196
rect 169760 527144 169812 527196
rect 472532 527144 472584 527196
rect 108304 527076 108356 527128
rect 372160 527076 372212 527128
rect 107568 527008 107620 527060
rect 333888 527008 333940 527060
rect 109040 526940 109092 526992
rect 312636 526940 312688 526992
rect 109132 526872 109184 526924
rect 283656 526872 283708 526924
rect 111064 526464 111116 526516
rect 211344 526464 211396 526516
rect 255412 526464 255464 526516
rect 283748 526464 283800 526516
rect 175924 526396 175976 526448
rect 433432 526396 433484 526448
rect 453304 526396 453356 526448
rect 463608 526396 463660 526448
rect 62856 525716 62908 525768
rect 66168 525920 66220 525972
rect 300768 525920 300820 525972
rect 499672 525920 499724 525972
rect 289728 525852 289780 525904
rect 498476 525852 498528 525904
rect 172428 525784 172480 525836
rect 505192 525784 505244 525836
rect 100760 525716 100812 525768
rect 379520 525716 379572 525768
rect 120080 525648 120132 525700
rect 351092 525648 351144 525700
rect 175924 525580 175976 525632
rect 386696 525580 386748 525632
rect 133788 525512 133840 525564
rect 325792 525512 325844 525564
rect 102140 525444 102192 525496
rect 274088 525444 274140 525496
rect 299388 525444 299440 525496
rect 372068 525444 372120 525496
rect 118700 525376 118752 525428
rect 274180 525376 274232 525428
rect 255320 525036 255372 525088
rect 298744 525036 298796 525088
rect 465816 525036 465868 525088
rect 513380 525036 513432 525088
rect 180248 524492 180300 524544
rect 508228 524492 508280 524544
rect 55772 524424 55824 524476
rect 58624 524424 58676 524476
rect 175188 524424 175240 524476
rect 506848 524424 506900 524476
rect 59176 524356 59228 524408
rect 380992 524356 381044 524408
rect 63500 524288 63552 524340
rect 378140 524288 378192 524340
rect 66168 524220 66220 524272
rect 375472 524220 375524 524272
rect 69664 524152 69716 524204
rect 375748 524152 375800 524204
rect 169760 524084 169812 524136
rect 383936 524084 383988 524136
rect 178040 524016 178092 524068
rect 382372 524016 382424 524068
rect 274640 523948 274692 524000
rect 297364 523948 297416 524000
rect 299388 523744 299440 523796
rect 481640 523744 481692 523796
rect 86868 522996 86920 523048
rect 92480 522996 92532 523048
rect 292580 522996 292632 523048
rect 313004 522996 313056 523048
rect 56508 522928 56560 522980
rect 386604 522928 386656 522980
rect 463608 522928 463660 522980
rect 467840 522928 467892 522980
rect 63500 522860 63552 522912
rect 385408 522860 385460 522912
rect 59912 522792 59964 522844
rect 375564 522792 375616 522844
rect 62120 522724 62172 522776
rect 378508 522724 378560 522776
rect 80060 522656 80112 522708
rect 371976 522656 372028 522708
rect 114468 522588 114520 522640
rect 382556 522588 382608 522640
rect 477408 522588 477460 522640
rect 503720 522588 503772 522640
rect 474280 522520 474332 522572
rect 504180 522520 504232 522572
rect 475936 522452 475988 522504
rect 506572 522452 506624 522504
rect 465724 522384 465776 522436
rect 497556 522384 497608 522436
rect 464436 522316 464488 522368
rect 502616 522316 502668 522368
rect 468760 522248 468812 522300
rect 510620 522248 510672 522300
rect 471888 521704 471940 521756
rect 490564 521704 490616 521756
rect 293960 521636 294012 521688
rect 494520 521636 494572 521688
rect 60740 521568 60792 521620
rect 62212 521568 62264 521620
rect 99380 521568 99432 521620
rect 385132 521568 385184 521620
rect 60832 521500 60884 521552
rect 62856 521500 62908 521552
rect 110420 521500 110472 521552
rect 383660 521500 383712 521552
rect 114468 521432 114520 521484
rect 385316 521432 385368 521484
rect 115756 521364 115808 521416
rect 382464 521364 382516 521416
rect 117228 521296 117280 521348
rect 301504 521296 301556 521348
rect 253296 521228 253348 521280
rect 256608 521228 256660 521280
rect 471336 521228 471388 521280
rect 504272 521228 504324 521280
rect 254584 521160 254636 521212
rect 276940 521160 276992 521212
rect 468484 521160 468536 521212
rect 505376 521160 505428 521212
rect 61936 521092 61988 521144
rect 86868 521092 86920 521144
rect 216128 521092 216180 521144
rect 281540 521092 281592 521144
rect 295984 521092 296036 521144
rect 367560 521092 367612 521144
rect 468668 521092 468720 521144
rect 512184 521092 512236 521144
rect 62028 521024 62080 521076
rect 255412 521024 255464 521076
rect 289084 521024 289136 521076
rect 366088 521024 366140 521076
rect 461768 521024 461820 521076
rect 505284 521024 505336 521076
rect 58808 520956 58860 521008
rect 255320 520956 255372 521008
rect 264244 520956 264296 521008
rect 370780 520956 370832 521008
rect 373908 520956 373960 521008
rect 381544 520956 381596 521008
rect 427084 520956 427136 521008
rect 475476 520956 475528 521008
rect 68284 520888 68336 520940
rect 294144 520888 294196 520940
rect 360844 520888 360896 520940
rect 474004 520888 474056 520940
rect 258448 520276 258500 520328
rect 431684 520276 431736 520328
rect 55128 520208 55180 520260
rect 137836 520208 137888 520260
rect 475384 520208 475436 520260
rect 479708 520208 479760 520260
rect 45928 520140 45980 520192
rect 289176 520140 289228 520192
rect 291016 520140 291068 520192
rect 383752 520140 383804 520192
rect 44180 520072 44232 520124
rect 50160 520004 50212 520056
rect 275376 520004 275428 520056
rect 282920 520072 282972 520124
rect 371884 520072 371936 520124
rect 283564 520004 283616 520056
rect 467840 520004 467892 520056
rect 480168 520004 480220 520056
rect 57704 519936 57756 519988
rect 271144 519936 271196 519988
rect 476028 519936 476080 519988
rect 494888 519936 494940 519988
rect 270408 519868 270460 519920
rect 385040 519868 385092 519920
rect 471244 519868 471296 519920
rect 494704 519868 494756 519920
rect 164148 519800 164200 519852
rect 273996 519800 274048 519852
rect 471428 519800 471480 519852
rect 495900 519800 495952 519852
rect 467288 519732 467340 519784
rect 498660 519732 498712 519784
rect 56140 519664 56192 519716
rect 138020 519664 138072 519716
rect 467196 519664 467248 519716
rect 500040 519664 500092 519716
rect 58440 519596 58492 519648
rect 154120 519596 154172 519648
rect 467104 519596 467156 519648
rect 500132 519596 500184 519648
rect 56508 519528 56560 519580
rect 162124 519528 162176 519580
rect 468576 519528 468628 519580
rect 509240 519528 509292 519580
rect 177948 519460 178000 519512
rect 483020 519460 483072 519512
rect 55128 518984 55180 519036
rect 58716 518984 58768 519036
rect 37924 518916 37976 518968
rect 56508 518916 56560 518968
rect 291844 518916 291896 518968
rect 494060 518916 494112 518968
rect 58900 518848 58952 518900
rect 389180 518848 389232 518900
rect 58992 518780 59044 518832
rect 386420 518780 386472 518832
rect 269028 518712 269080 518764
rect 385224 518712 385276 518764
rect 481640 518576 481692 518628
rect 482100 518576 482152 518628
rect 478788 518508 478840 518560
rect 491392 518508 491444 518560
rect 477408 518440 477460 518492
rect 490656 518440 490708 518492
rect 477316 518372 477368 518424
rect 492680 518372 492732 518424
rect 480076 518304 480128 518356
rect 482100 518304 482152 518356
rect 59544 518236 59596 518288
rect 171140 518236 171192 518288
rect 476764 518236 476816 518288
rect 493416 518236 493468 518288
rect 56784 518168 56836 518220
rect 62028 518168 62080 518220
rect 60924 518100 60976 518152
rect 61936 518100 61988 518152
rect 374644 518168 374696 518220
rect 474096 518168 474148 518220
rect 491852 518168 491904 518220
rect 476120 518100 476172 518152
rect 494796 518100 494848 518152
rect 478788 518032 478840 518084
rect 483112 518032 483164 518084
rect 478972 517964 479024 518016
rect 480076 517964 480128 518016
rect 58992 517828 59044 517880
rect 60924 517624 60976 517676
rect 57704 517556 57756 517608
rect 60832 517556 60884 517608
rect 60372 517488 60424 517540
rect 60740 517488 60792 517540
rect 57428 517012 57480 517064
rect 56508 516128 56560 516180
rect 57244 516128 57296 516180
rect 56968 511980 57020 512032
rect 58440 511980 58492 512032
rect 481640 510552 481692 510604
rect 483112 510552 483164 510604
rect 482100 510484 482152 510536
rect 482560 510484 482612 510536
rect 482836 506404 482888 506456
rect 491392 506404 491444 506456
rect 482928 506336 482980 506388
rect 490656 506336 490708 506388
rect 57704 500896 57756 500948
rect 58808 500896 58860 500948
rect 482836 500896 482888 500948
rect 494060 500896 494112 500948
rect 482928 500828 482980 500880
rect 492680 500828 492732 500880
rect 56876 499672 56928 499724
rect 57152 499672 57204 499724
rect 57060 490560 57112 490612
rect 57336 490560 57388 490612
rect 482100 480156 482152 480208
rect 494796 480156 494848 480208
rect 482100 478796 482152 478848
rect 497556 478796 497608 478848
rect 479248 477980 479300 478032
rect 479524 477980 479576 478032
rect 3424 476008 3476 476060
rect 37924 476008 37976 476060
rect 482100 474648 482152 474700
rect 485872 474648 485924 474700
rect 482100 473288 482152 473340
rect 488816 473288 488868 473340
rect 482100 471928 482152 471980
rect 498660 471928 498712 471980
rect 482008 471860 482060 471912
rect 487436 471860 487488 471912
rect 482100 470500 482152 470552
rect 500132 470500 500184 470552
rect 482008 470432 482060 470484
rect 486700 470432 486752 470484
rect 482100 469140 482152 469192
rect 500040 469140 500092 469192
rect 482008 469072 482060 469124
rect 494704 469072 494756 469124
rect 482100 467780 482152 467832
rect 487252 467780 487304 467832
rect 482008 467712 482060 467764
rect 487344 467712 487396 467764
rect 482008 464992 482060 465044
rect 505376 464992 505428 465044
rect 482100 464924 482152 464976
rect 504272 464924 504324 464976
rect 482100 464788 482152 464840
rect 489368 464788 489420 464840
rect 482100 463632 482152 463684
rect 490196 463632 490248 463684
rect 482100 463292 482152 463344
rect 488080 463292 488132 463344
rect 482008 462272 482060 462324
rect 505284 462272 505336 462324
rect 481916 462204 481968 462256
rect 502616 462204 502668 462256
rect 482100 462136 482152 462188
rect 490104 462136 490156 462188
rect 482100 460776 482152 460828
rect 488632 460776 488684 460828
rect 482008 459484 482060 459536
rect 504180 459484 504232 459536
rect 482100 459416 482152 459468
rect 495900 459416 495952 459468
rect 482008 458124 482060 458176
rect 491852 458124 491904 458176
rect 482100 458056 482152 458108
rect 490012 458056 490064 458108
rect 482100 456696 482152 456748
rect 509424 456696 509476 456748
rect 482008 455336 482060 455388
rect 493416 455336 493468 455388
rect 482100 455268 482152 455320
rect 489920 455268 489972 455320
rect 482100 453976 482152 454028
rect 491668 453976 491720 454028
rect 482100 452548 482152 452600
rect 497464 452548 497516 452600
rect 482100 452412 482152 452464
rect 489276 452412 489328 452464
rect 482192 449828 482244 449880
rect 509332 449828 509384 449880
rect 482100 449760 482152 449812
rect 494520 449760 494572 449812
rect 482192 449692 482244 449744
rect 493232 449692 493284 449744
rect 482192 448468 482244 448520
rect 494428 448468 494480 448520
rect 482100 448400 482152 448452
rect 490564 448400 490616 448452
rect 482008 447040 482060 447092
rect 508136 447040 508188 447092
rect 482100 446972 482152 447024
rect 493048 446972 493100 447024
rect 482192 446904 482244 446956
rect 491760 446904 491812 446956
rect 482100 445680 482152 445732
rect 493324 445680 493376 445732
rect 482192 445612 482244 445664
rect 493140 445612 493192 445664
rect 482192 444320 482244 444372
rect 492772 444320 492824 444372
rect 482100 444252 482152 444304
rect 492864 444252 492916 444304
rect 482192 442892 482244 442944
rect 506848 442892 506900 442944
rect 482100 441532 482152 441584
rect 508228 441532 508280 441584
rect 482192 441464 482244 441516
rect 492956 441464 493008 441516
rect 482192 440172 482244 440224
rect 505192 440172 505244 440224
rect 482100 438812 482152 438864
rect 506756 438812 506808 438864
rect 482192 438744 482244 438796
rect 502524 438744 502576 438796
rect 482192 428204 482244 428256
rect 482836 428204 482888 428256
rect 482836 425008 482888 425060
rect 491300 425008 491352 425060
rect 482836 423580 482888 423632
rect 491484 423580 491536 423632
rect 482836 423308 482888 423360
rect 486148 423308 486200 423360
rect 3424 422288 3476 422340
rect 26884 422288 26936 422340
rect 482836 418072 482888 418124
rect 494244 418072 494296 418124
rect 482192 418004 482244 418056
rect 494336 418004 494388 418056
rect 482836 416712 482888 416764
rect 499856 416712 499908 416764
rect 482836 415352 482888 415404
rect 497188 415352 497240 415404
rect 482192 415284 482244 415336
rect 497280 415284 497332 415336
rect 482192 413924 482244 413976
rect 498476 413924 498528 413976
rect 482836 413856 482888 413908
rect 497096 413856 497148 413908
rect 482836 412496 482888 412548
rect 487988 412496 488040 412548
rect 482836 411204 482888 411256
rect 503996 411204 504048 411256
rect 482192 411136 482244 411188
rect 486056 411136 486108 411188
rect 482192 410932 482244 410984
rect 487804 410932 487856 410984
rect 482836 409776 482888 409828
rect 487896 409776 487948 409828
rect 482836 408416 482888 408468
rect 502340 408416 502392 408468
rect 482192 408348 482244 408400
rect 487620 408348 487672 408400
rect 482836 407056 482888 407108
rect 499672 407056 499724 407108
rect 482192 406988 482244 407040
rect 497004 406988 497056 407040
rect 482836 405628 482888 405680
rect 494152 405628 494204 405680
rect 482836 402908 482888 402960
rect 501144 402908 501196 402960
rect 482836 401548 482888 401600
rect 502432 401548 502484 401600
rect 482836 401276 482888 401328
rect 489092 401276 489144 401328
rect 482192 400120 482244 400172
rect 496912 400120 496964 400172
rect 482836 400052 482888 400104
rect 495440 400052 495492 400104
rect 482008 398760 482060 398812
rect 500960 398760 501012 398812
rect 482836 398692 482888 398744
rect 498292 398692 498344 398744
rect 482192 398624 482244 398676
rect 493508 398624 493560 398676
rect 482836 397400 482888 397452
rect 503904 397400 503956 397452
rect 482192 397332 482244 397384
rect 495532 397332 495584 397384
rect 482192 395972 482244 396024
rect 514852 395972 514904 396024
rect 482836 395904 482888 395956
rect 501052 395904 501104 395956
rect 482192 394612 482244 394664
rect 514760 394612 514812 394664
rect 482836 394544 482888 394596
rect 512092 394544 512144 394596
rect 482192 393252 482244 393304
rect 482652 393252 482704 393304
rect 482836 393252 482888 393304
rect 513380 393252 513432 393304
rect 482100 393184 482152 393236
rect 509240 393184 509292 393236
rect 482928 393116 482980 393168
rect 506664 393116 506716 393168
rect 482836 391892 482888 391944
rect 512000 391892 512052 391944
rect 482928 391824 482980 391876
rect 512184 391824 512236 391876
rect 482928 390464 482980 390516
rect 510620 390464 510672 390516
rect 58808 389852 58860 389904
rect 122104 389852 122156 389904
rect 60372 389784 60424 389836
rect 265624 389784 265676 389836
rect 474648 389104 474700 389156
rect 546500 389104 546552 389156
rect 26884 388424 26936 388476
rect 95700 388424 95752 388476
rect 118700 387744 118752 387796
rect 534724 387744 534776 387796
rect 57244 387676 57296 387728
rect 150440 387676 150492 387728
rect 272524 387676 272576 387728
rect 506480 387676 506532 387728
rect 58716 387608 58768 387660
rect 143540 387608 143592 387660
rect 144368 387608 144420 387660
rect 274640 387608 274692 387660
rect 505100 387608 505152 387660
rect 56140 387540 56192 387592
rect 132500 387540 132552 387592
rect 137192 387540 137244 387592
rect 270408 387540 270460 387592
rect 482652 387540 482704 387592
rect 498200 387540 498252 387592
rect 498844 387540 498896 387592
rect 60556 387472 60608 387524
rect 124128 387472 124180 387524
rect 106188 387336 106240 387388
rect 147680 387336 147732 387388
rect 108304 387268 108356 387320
rect 162308 387268 162360 387320
rect 162768 387268 162820 387320
rect 60280 387200 60332 387252
rect 140780 387200 140832 387252
rect 62120 387132 62172 387184
rect 154580 387132 154632 387184
rect 155132 387132 155184 387184
rect 277216 387132 277268 387184
rect 445760 387132 445812 387184
rect 115848 387064 115900 387116
rect 498200 387064 498252 387116
rect 458824 386860 458876 386912
rect 460112 386860 460164 386912
rect 138664 386452 138716 386504
rect 191012 386452 191064 386504
rect 191748 386452 191800 386504
rect 105544 386384 105596 386436
rect 177304 386384 177356 386436
rect 471980 386316 472032 386368
rect 479616 386316 479668 386368
rect 162768 384956 162820 385008
rect 543832 384956 543884 385008
rect 191748 384888 191800 384940
rect 547972 384888 548024 384940
rect 84108 384276 84160 384328
rect 132500 384412 132552 384464
rect 177304 383596 177356 383648
rect 547880 383596 547932 383648
rect 122104 382916 122156 382968
rect 127624 382916 127676 382968
rect 449900 382916 449952 382968
rect 471980 382916 472032 382968
rect 282828 380808 282880 380860
rect 539968 380808 540020 380860
rect 127624 378088 127676 378140
rect 133144 378088 133196 378140
rect 260748 378088 260800 378140
rect 529388 378088 529440 378140
rect 282828 378020 282880 378072
rect 539876 378020 539928 378072
rect 265624 377408 265676 377460
rect 272524 377408 272576 377460
rect 438768 375980 438820 376032
rect 449900 375980 449952 376032
rect 427912 373260 427964 373312
rect 438768 373260 438820 373312
rect 426348 369928 426400 369980
rect 427912 369928 427964 369980
rect 133144 368432 133196 368484
rect 138020 368432 138072 368484
rect 420184 367752 420236 367804
rect 426348 367752 426400 367804
rect 138020 365644 138072 365696
rect 141424 365644 141476 365696
rect 417516 358708 417568 358760
rect 420184 358708 420236 358760
rect 72608 355308 72660 355360
rect 506572 355308 506624 355360
rect 141424 354696 141476 354748
rect 144184 354696 144236 354748
rect 498844 353200 498896 353252
rect 580172 353200 580224 353252
rect 272524 351160 272576 351212
rect 287704 351160 287756 351212
rect 410524 347012 410576 347064
rect 417516 347012 417568 347064
rect 56968 345652 57020 345704
rect 288532 345652 288584 345704
rect 242808 344972 242860 345024
rect 410524 344972 410576 345024
rect 76564 344292 76616 344344
rect 494704 344292 494756 344344
rect 263600 343952 263652 344004
rect 284300 343952 284352 344004
rect 256700 343884 256752 343936
rect 280252 343884 280304 343936
rect 253204 343816 253256 343868
rect 283196 343816 283248 343868
rect 255320 343748 255372 343800
rect 287520 343748 287572 343800
rect 220176 343680 220228 343732
rect 285956 343680 286008 343732
rect 144184 343612 144236 343664
rect 147588 343612 147640 343664
rect 220084 343612 220136 343664
rect 286048 343612 286100 343664
rect 251088 343068 251140 343120
rect 284392 343068 284444 343120
rect 249708 343000 249760 343052
rect 283288 343000 283340 343052
rect 245660 342932 245712 342984
rect 283104 342932 283156 342984
rect 247040 342864 247092 342916
rect 284484 342864 284536 342916
rect 243544 342796 243596 342848
rect 285680 342796 285732 342848
rect 244280 342728 244332 342780
rect 287612 342728 287664 342780
rect 240048 342660 240100 342712
rect 283012 342660 283064 342712
rect 231216 342592 231268 342644
rect 281540 342592 281592 342644
rect 231400 342524 231452 342576
rect 284944 342524 284996 342576
rect 226340 342456 226392 342508
rect 284852 342456 284904 342508
rect 223028 342388 223080 342440
rect 283564 342388 283616 342440
rect 226616 342320 226668 342372
rect 287428 342320 287480 342372
rect 220268 342252 220320 342304
rect 285864 342252 285916 342304
rect 240048 341776 240100 341828
rect 280620 341776 280672 341828
rect 237472 341708 237524 341760
rect 280344 341708 280396 341760
rect 58624 341640 58676 341692
rect 287060 341640 287112 341692
rect 236644 341572 236696 341624
rect 490748 341572 490800 341624
rect 236920 341504 236972 341556
rect 507308 341504 507360 341556
rect 237380 341436 237432 341488
rect 280712 341436 280764 341488
rect 240784 341368 240836 341420
rect 291844 341368 291896 341420
rect 227812 341300 227864 341352
rect 284760 341300 284812 341352
rect 225696 341232 225748 341284
rect 284576 341232 284628 341284
rect 223120 341164 223172 341216
rect 283472 341164 283524 341216
rect 224960 341096 225012 341148
rect 291384 341096 291436 341148
rect 225052 341028 225104 341080
rect 291292 341028 291344 341080
rect 227720 340960 227772 341012
rect 295340 340960 295392 341012
rect 225144 340892 225196 340944
rect 292580 340892 292632 340944
rect 147588 340824 147640 340876
rect 154488 340824 154540 340876
rect 239864 340348 239916 340400
rect 280988 340348 281040 340400
rect 238392 340280 238444 340332
rect 502984 340280 503036 340332
rect 237104 340212 237156 340264
rect 580356 340212 580408 340264
rect 79324 340144 79376 340196
rect 79784 340144 79836 340196
rect 503720 340144 503772 340196
rect 237472 340076 237524 340128
rect 280436 340076 280488 340128
rect 237564 340008 237616 340060
rect 280804 340008 280856 340060
rect 239956 339940 240008 339992
rect 285036 339940 285088 339992
rect 240048 339872 240100 339924
rect 285772 339872 285824 339924
rect 237380 339804 237432 339856
rect 284668 339804 284720 339856
rect 228456 339736 228508 339788
rect 281724 339736 281776 339788
rect 225880 339668 225932 339720
rect 283380 339668 283432 339720
rect 223488 339600 223540 339652
rect 283656 339600 283708 339652
rect 223396 339532 223448 339584
rect 283748 339532 283800 339584
rect 235724 339464 235776 339516
rect 580264 339464 580316 339516
rect 231308 339396 231360 339448
rect 281632 339396 281684 339448
rect 239128 338512 239180 338564
rect 239864 338512 239916 338564
rect 238024 337356 238076 337408
rect 238392 337356 238444 337408
rect 154488 336676 154540 336728
rect 158812 336676 158864 336728
rect 158812 332392 158864 332444
rect 162124 332392 162176 332444
rect 162124 321580 162176 321632
rect 166264 321580 166316 321632
rect 94044 312536 94096 312588
rect 158720 312536 158772 312588
rect 92388 311108 92440 311160
rect 154580 311108 154632 311160
rect 90732 309748 90784 309800
rect 150440 309748 150492 309800
rect 87420 308388 87472 308440
rect 143540 308388 143592 308440
rect 85764 307028 85816 307080
rect 140780 307028 140832 307080
rect 82452 304240 82504 304292
rect 132500 304240 132552 304292
rect 80796 302880 80848 302932
rect 129740 302880 129792 302932
rect 75828 300092 75880 300144
rect 119344 300092 119396 300144
rect 282184 299412 282236 299464
rect 285036 299412 285088 299464
rect 74172 297372 74224 297424
rect 115204 297372 115256 297424
rect 166264 292544 166316 292596
rect 169024 292544 169076 292596
rect 496728 291796 496780 291848
rect 503720 291796 503772 291848
rect 282184 289756 282236 289808
rect 284944 289756 284996 289808
rect 282092 288328 282144 288380
rect 284852 288328 284904 288380
rect 282736 288260 282788 288312
rect 286048 288260 286100 288312
rect 282644 286696 282696 286748
rect 285956 286696 286008 286748
rect 281540 285608 281592 285660
rect 283748 285608 283800 285660
rect 282644 285540 282696 285592
rect 285864 285540 285916 285592
rect 282092 284248 282144 284300
rect 284760 284248 284812 284300
rect 77484 282140 77536 282192
rect 122840 282140 122892 282192
rect 282000 281460 282052 281512
rect 284576 281460 284628 281512
rect 282000 280100 282052 280152
rect 284668 280100 284720 280152
rect 70860 279420 70912 279472
rect 108304 279420 108356 279472
rect 169024 279420 169076 279472
rect 182824 279420 182876 279472
rect 282828 277448 282880 277500
rect 288624 277448 288676 277500
rect 282828 276088 282880 276140
rect 288716 276088 288768 276140
rect 282736 276020 282788 276072
rect 289912 276020 289964 276072
rect 493968 275272 494020 275324
rect 506480 275272 506532 275324
rect 282828 274660 282880 274712
rect 287152 274660 287204 274712
rect 282828 273300 282880 273352
rect 287244 273300 287296 273352
rect 282736 273232 282788 273284
rect 290004 273232 290056 273284
rect 282828 271872 282880 271924
rect 287336 271872 287388 271924
rect 69204 271192 69256 271244
rect 105636 271192 105688 271244
rect 89076 271124 89128 271176
rect 147680 271124 147732 271176
rect 282828 270580 282880 270632
rect 291568 270580 291620 270632
rect 282736 270512 282788 270564
rect 291476 270512 291528 270564
rect 281908 270444 281960 270496
rect 284484 270444 284536 270496
rect 281908 267656 281960 267708
rect 284392 267656 284444 267708
rect 281816 266296 281868 266348
rect 284300 266296 284352 266348
rect 54668 262964 54720 263016
rect 72424 262964 72476 263016
rect 56324 262896 56376 262948
rect 76564 262896 76616 262948
rect 57888 262828 57940 262880
rect 79324 262828 79376 262880
rect 282828 262148 282880 262200
rect 287612 262148 287664 262200
rect 39948 261468 40000 261520
rect 233976 261468 234028 261520
rect 11704 260856 11756 260908
rect 102140 260856 102192 260908
rect 282552 260788 282604 260840
rect 285680 260788 285732 260840
rect 282552 257456 282604 257508
rect 285772 257456 285824 257508
rect 282828 256640 282880 256692
rect 287520 256640 287572 256692
rect 282828 253852 282880 253904
rect 287428 253852 287480 253904
rect 182824 249704 182876 249756
rect 189724 249704 189776 249756
rect 496728 245556 496780 245608
rect 580172 245556 580224 245608
rect 282828 242904 282880 242956
rect 288900 242904 288952 242956
rect 189724 235220 189776 235272
rect 207664 235220 207716 235272
rect 282184 229100 282236 229152
rect 284944 229100 284996 229152
rect 282276 227740 282328 227792
rect 285128 227740 285180 227792
rect 282828 219444 282880 219496
rect 290464 219444 290516 219496
rect 3424 215228 3476 215280
rect 11704 215228 11756 215280
rect 111064 214548 111116 214600
rect 158720 214548 158772 214600
rect 233884 213936 233936 213988
rect 237380 213936 237432 213988
rect 207664 211760 207716 211812
rect 218704 211760 218756 211812
rect 282828 211148 282880 211200
rect 288992 211148 289044 211200
rect 494704 206932 494756 206984
rect 580172 206932 580224 206984
rect 282828 204280 282880 204332
rect 291752 204280 291804 204332
rect 233976 201424 234028 201476
rect 237380 201424 237432 201476
rect 48228 200064 48280 200116
rect 110420 200064 110472 200116
rect 111064 200064 111116 200116
rect 218704 199996 218756 200048
rect 237380 199996 237432 200048
rect 104900 199928 104952 199980
rect 231032 199928 231084 199980
rect 106280 199860 106332 199912
rect 231308 199860 231360 199912
rect 95240 199792 95292 199844
rect 220084 199792 220136 199844
rect 100668 199724 100720 199776
rect 220176 199724 220228 199776
rect 103428 199656 103480 199708
rect 220268 199656 220320 199708
rect 94504 199588 94556 199640
rect 223028 199588 223080 199640
rect 107660 199520 107712 199572
rect 228456 199520 228508 199572
rect 88340 198636 88392 198688
rect 225880 198636 225932 198688
rect 86960 198568 87012 198620
rect 223488 198568 223540 198620
rect 98000 198500 98052 198552
rect 225696 198500 225748 198552
rect 96620 198432 96672 198484
rect 223120 198432 223172 198484
rect 104164 198364 104216 198416
rect 223396 198364 223448 198416
rect 85580 197684 85632 197736
rect 238668 197684 238720 197736
rect 78588 197616 78640 197668
rect 235448 197616 235500 197668
rect 79324 197548 79376 197600
rect 238484 197548 238536 197600
rect 70400 197480 70452 197532
rect 235356 197480 235408 197532
rect 73160 197412 73212 197464
rect 238300 197412 238352 197464
rect 71780 197344 71832 197396
rect 238208 197344 238260 197396
rect 287704 187688 287756 187740
rect 291200 187688 291252 187740
rect 282460 178032 282512 178084
rect 283748 178032 283800 178084
rect 282828 176672 282880 176724
rect 289176 176672 289228 176724
rect 282828 172456 282880 172508
rect 295340 172456 295392 172508
rect 282736 172388 282788 172440
rect 291384 172388 291436 172440
rect 282828 171028 282880 171080
rect 292580 171028 292632 171080
rect 282828 169668 282880 169720
rect 291292 169668 291344 169720
rect 282828 169532 282880 169584
rect 287060 169532 287112 169584
rect 282736 168308 282788 168360
rect 291200 168308 291252 168360
rect 282828 168240 282880 168292
rect 288532 168240 288584 168292
rect 493968 166948 494020 167000
rect 580172 166948 580224 167000
rect 232688 141992 232740 142044
rect 236828 141992 236880 142044
rect 238484 140632 238536 140684
rect 580448 140632 580500 140684
rect 237748 140564 237800 140616
rect 580356 140564 580408 140616
rect 238576 140496 238628 140548
rect 580264 140496 580316 140548
rect 239680 140428 239732 140480
rect 580540 140428 580592 140480
rect 239588 140360 239640 140412
rect 458824 140360 458876 140412
rect 235356 140292 235408 140344
rect 291568 140292 291620 140344
rect 235448 140224 235500 140276
rect 291476 140224 291528 140276
rect 235908 140156 235960 140208
rect 289176 140156 289228 140208
rect 238024 140088 238076 140140
rect 287244 140088 287296 140140
rect 238116 140020 238168 140072
rect 287336 140020 287388 140072
rect 266912 139952 266964 140004
rect 283748 139952 283800 140004
rect 238208 139340 238260 139392
rect 470876 139340 470928 139392
rect 240784 139272 240836 139324
rect 467288 139272 467340 139324
rect 205640 139204 205692 139256
rect 288992 139204 289044 139256
rect 215300 139136 215352 139188
rect 290464 139136 290516 139188
rect 218060 139068 218112 139120
rect 282184 139068 282236 139120
rect 235908 139000 235960 139052
rect 288716 139000 288768 139052
rect 235632 138932 235684 138984
rect 287152 138932 287204 138984
rect 233148 138864 233200 138916
rect 283380 138864 283432 138916
rect 238760 138796 238812 138848
rect 288900 138796 288952 138848
rect 235816 138728 235868 138780
rect 285128 138728 285180 138780
rect 235908 138660 235960 138712
rect 284944 138660 284996 138712
rect 235724 138592 235776 138644
rect 282092 138592 282144 138644
rect 251180 138524 251232 138576
rect 280344 138524 280396 138576
rect 237380 137912 237432 137964
rect 249800 137912 249852 137964
rect 262128 137912 262180 137964
rect 288624 137912 288676 137964
rect 66168 137844 66220 137896
rect 245016 137844 245068 137896
rect 247040 137844 247092 137896
rect 250996 137844 251048 137896
rect 115848 137776 115900 137828
rect 246212 137776 246264 137828
rect 118700 137708 118752 137760
rect 247408 137708 247460 137760
rect 233148 137640 233200 137692
rect 248604 137640 248656 137692
rect 44180 137572 44232 137624
rect 243820 137572 243872 137624
rect 271144 136620 271196 136672
rect 272524 136620 272576 136672
rect 73068 87320 73120 87372
rect 345664 87320 345716 87372
rect 74448 87252 74500 87304
rect 86316 87252 86368 87304
rect 66996 87184 67048 87236
rect 84936 87184 84988 87236
rect 70124 87116 70176 87168
rect 98736 87116 98788 87168
rect 76472 87048 76524 87100
rect 287704 87048 287756 87100
rect 82728 86980 82780 87032
rect 90456 86980 90508 87032
rect 84936 83444 84988 83496
rect 336280 83444 336332 83496
rect 84200 82764 84252 82816
rect 295984 82764 296036 82816
rect 86316 69640 86368 69692
rect 350448 69640 350500 69692
rect 88248 51688 88300 51740
rect 110420 51688 110472 51740
rect 90456 50328 90508 50380
rect 368204 50328 368256 50380
rect 572 40672 624 40724
rect 86960 40672 87012 40724
rect 98736 10276 98788 10328
rect 339868 10276 339920 10328
rect 291844 6808 291896 6860
rect 580172 6808 580224 6860
rect 287704 4768 287756 4820
rect 354036 4768 354088 4820
rect 345664 4156 345716 4208
rect 346952 4156 347004 4208
rect 241428 4088 241480 4140
rect 282920 4088 282972 4140
rect 264980 4020 265032 4072
rect 291752 4020 291804 4072
rect 295984 3408 296036 3460
rect 371700 3408 371752 3460
rect 442264 3408 442316 3460
rect 583392 3408 583444 3460
rect 438860 2796 438912 2848
rect 581000 2796 581052 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3424 632732 3476 632738
rect 3424 632674 3476 632680
rect 3436 632097 3464 632674
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 579698 3464 579935
rect 3424 579692 3476 579698
rect 3424 579634 3476 579640
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3424 476060 3476 476066
rect 3424 476002 3476 476008
rect 3436 475697 3464 476002
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 4066 410000 4122 410009
rect 4066 409935 4122 409944
rect 3974 398168 4030 398177
rect 3974 398103 4030 398112
rect 3988 382945 4016 398103
rect 3974 382936 4030 382945
rect 3974 382871 4030 382880
rect 4080 376145 4108 409935
rect 4066 376136 4122 376145
rect 4066 376071 4122 376080
rect 8128 316713 8156 703520
rect 24320 700369 24348 703520
rect 40512 701010 40540 703520
rect 40500 701004 40552 701010
rect 40500 700946 40552 700952
rect 59268 701004 59320 701010
rect 59268 700946 59320 700952
rect 24306 700360 24362 700369
rect 24306 700295 24362 700304
rect 32402 700360 32458 700369
rect 32402 700295 32458 700304
rect 28906 650040 28962 650049
rect 28906 649975 28962 649984
rect 26884 422340 26936 422346
rect 26884 422282 26936 422288
rect 26896 388482 26924 422282
rect 28920 395321 28948 649975
rect 31666 643648 31722 643657
rect 31666 643583 31722 643592
rect 31574 559736 31630 559745
rect 31574 559671 31630 559680
rect 31482 541104 31538 541113
rect 31482 541039 31538 541048
rect 30286 533352 30342 533361
rect 30286 533287 30342 533296
rect 28906 395312 28962 395321
rect 28906 395247 28962 395256
rect 26884 388476 26936 388482
rect 26884 388418 26936 388424
rect 30300 341601 30328 533287
rect 31390 522064 31446 522073
rect 31390 521999 31446 522008
rect 31404 501945 31432 521999
rect 31390 501936 31446 501945
rect 31390 501871 31446 501880
rect 31496 486713 31524 541039
rect 31588 487257 31616 559671
rect 31574 487248 31630 487257
rect 31574 487183 31630 487192
rect 31482 486704 31538 486713
rect 31482 486639 31538 486648
rect 31680 390425 31708 643583
rect 31666 390416 31722 390425
rect 31666 390351 31722 390360
rect 32416 341873 32444 700295
rect 59280 699825 59308 700946
rect 59266 699816 59322 699825
rect 59266 699751 59322 699760
rect 55220 683188 55272 683194
rect 55220 683130 55272 683136
rect 38566 650176 38622 650185
rect 38566 650111 38622 650120
rect 37186 648680 37242 648689
rect 37186 648615 37242 648624
rect 34426 648408 34482 648417
rect 34426 648343 34482 648352
rect 34334 551168 34390 551177
rect 34334 551103 34390 551112
rect 34242 545728 34298 545737
rect 34242 545663 34298 545672
rect 33046 534168 33102 534177
rect 33046 534103 33102 534112
rect 32862 527368 32918 527377
rect 32862 527303 32918 527312
rect 32876 503577 32904 527303
rect 32954 524512 33010 524521
rect 32954 524447 33010 524456
rect 32862 503568 32918 503577
rect 32862 503503 32918 503512
rect 32968 493785 32996 524447
rect 32954 493776 33010 493785
rect 32954 493711 33010 493720
rect 32402 341864 32458 341873
rect 32402 341799 32458 341808
rect 33060 341737 33088 534103
rect 34150 533080 34206 533089
rect 34150 533015 34206 533024
rect 34058 530632 34114 530641
rect 34058 530567 34114 530576
rect 34072 498137 34100 530567
rect 34058 498128 34114 498137
rect 34058 498063 34114 498072
rect 34164 427417 34192 533015
rect 34256 437209 34284 545663
rect 34242 437200 34298 437209
rect 34242 437135 34298 437144
rect 34348 428505 34376 551103
rect 34334 428496 34390 428505
rect 34334 428431 34390 428440
rect 34150 427408 34206 427417
rect 34150 427343 34206 427352
rect 34440 390969 34468 648343
rect 35806 647456 35862 647465
rect 35806 647391 35862 647400
rect 35714 645552 35770 645561
rect 35714 645487 35770 645496
rect 35622 641744 35678 641753
rect 35622 641679 35678 641688
rect 35438 552528 35494 552537
rect 35438 552463 35494 552472
rect 35346 545456 35402 545465
rect 35346 545391 35402 545400
rect 35360 462233 35388 545391
rect 35452 464409 35480 552463
rect 35530 539880 35586 539889
rect 35530 539815 35586 539824
rect 35438 464400 35494 464409
rect 35438 464335 35494 464344
rect 35346 462224 35402 462233
rect 35346 462159 35402 462168
rect 35544 426329 35572 539815
rect 35636 479641 35664 641679
rect 35728 481273 35756 645487
rect 35714 481264 35770 481273
rect 35714 481199 35770 481208
rect 35622 479632 35678 479641
rect 35622 479567 35678 479576
rect 35530 426320 35586 426329
rect 35530 426255 35586 426264
rect 35820 391513 35848 647391
rect 37002 645960 37058 645969
rect 37002 645895 37058 645904
rect 36910 645144 36966 645153
rect 36910 645079 36966 645088
rect 36818 641336 36874 641345
rect 36818 641271 36874 641280
rect 36634 548176 36690 548185
rect 36634 548111 36690 548120
rect 36648 464953 36676 548111
rect 36726 530224 36782 530233
rect 36726 530159 36782 530168
rect 36634 464944 36690 464953
rect 36634 464879 36690 464888
rect 36740 427961 36768 530159
rect 36832 511193 36860 641271
rect 36818 511184 36874 511193
rect 36818 511119 36874 511128
rect 36924 482361 36952 645079
rect 36910 482352 36966 482361
rect 36910 482287 36966 482296
rect 37016 480729 37044 645895
rect 37094 640520 37150 640529
rect 37094 640455 37150 640464
rect 37002 480720 37058 480729
rect 37002 480655 37058 480664
rect 37108 463321 37136 640455
rect 37094 463312 37150 463321
rect 37094 463247 37150 463256
rect 36726 427952 36782 427961
rect 36726 427887 36782 427896
rect 37200 392057 37228 648615
rect 38474 546544 38530 546553
rect 38474 546479 38530 546488
rect 38198 545184 38254 545193
rect 38198 545119 38254 545128
rect 38106 523288 38162 523297
rect 38106 523223 38162 523232
rect 37924 518968 37976 518974
rect 37924 518910 37976 518916
rect 37936 476066 37964 518910
rect 38120 492833 38148 523223
rect 38212 496505 38240 545119
rect 38382 540016 38438 540025
rect 38382 539951 38438 539960
rect 38290 530360 38346 530369
rect 38290 530295 38346 530304
rect 38198 496496 38254 496505
rect 38198 496431 38254 496440
rect 38106 492824 38162 492833
rect 38106 492759 38162 492768
rect 38304 477465 38332 530295
rect 38290 477456 38346 477465
rect 38290 477391 38346 477400
rect 37924 476060 37976 476066
rect 37924 476002 37976 476008
rect 38396 474745 38424 539951
rect 38382 474736 38438 474745
rect 38382 474671 38438 474680
rect 38488 398585 38516 546479
rect 38580 475833 38608 650111
rect 50802 646776 50858 646785
rect 50802 646711 50858 646720
rect 46846 644192 46902 644201
rect 46846 644127 46902 644136
rect 45282 644056 45338 644065
rect 45282 643991 45338 644000
rect 42614 642696 42670 642705
rect 42614 642631 42670 642640
rect 41326 639976 41382 639985
rect 41326 639911 41382 639920
rect 39854 637800 39910 637809
rect 39854 637735 39910 637744
rect 39762 551440 39818 551449
rect 39762 551375 39818 551384
rect 39670 542464 39726 542473
rect 39670 542399 39726 542408
rect 39394 533624 39450 533633
rect 39394 533559 39450 533568
rect 39408 478553 39436 533559
rect 39578 531584 39634 531593
rect 39578 531519 39634 531528
rect 39486 531312 39542 531321
rect 39486 531247 39542 531256
rect 39394 478544 39450 478553
rect 39394 478479 39450 478488
rect 38566 475824 38622 475833
rect 38566 475759 38622 475768
rect 39500 418713 39528 531247
rect 39486 418704 39542 418713
rect 39486 418639 39542 418648
rect 39592 411097 39620 531519
rect 39578 411088 39634 411097
rect 39578 411023 39634 411032
rect 39684 399129 39712 542399
rect 39670 399120 39726 399129
rect 39670 399055 39726 399064
rect 38474 398576 38530 398585
rect 38474 398511 38530 398520
rect 39776 396953 39804 551375
rect 39868 472025 39896 637735
rect 39948 635520 40000 635526
rect 39948 635462 40000 635468
rect 39854 472016 39910 472025
rect 39854 471951 39910 471960
rect 39762 396944 39818 396953
rect 39762 396879 39818 396888
rect 37186 392048 37242 392057
rect 37186 391983 37242 391992
rect 35806 391504 35862 391513
rect 35806 391439 35862 391448
rect 34426 390960 34482 390969
rect 34426 390895 34482 390904
rect 33046 341728 33102 341737
rect 33046 341663 33102 341672
rect 30286 341592 30342 341601
rect 30286 341527 30342 341536
rect 8114 316704 8170 316713
rect 8114 316639 8170 316648
rect 4802 262304 4858 262313
rect 4802 262239 4858 262248
rect 3424 215280 3476 215286
rect 3424 215222 3476 215228
rect 3436 214985 3464 215222
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 2870 91760 2926 91769
rect 2870 91695 2926 91704
rect 572 40724 624 40730
rect 572 40666 624 40672
rect 584 480 612 40666
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 480 1716 3431
rect 2884 480 2912 91695
rect 4816 32473 4844 262239
rect 39960 261526 39988 635462
rect 41050 545320 41106 545329
rect 41050 545255 41106 545264
rect 40774 531720 40830 531729
rect 40774 531655 40830 531664
rect 40590 526008 40646 526017
rect 40590 525943 40646 525952
rect 40498 522744 40554 522753
rect 40498 522679 40554 522688
rect 40512 498953 40540 522679
rect 40498 498944 40554 498953
rect 40498 498879 40554 498888
rect 40604 498817 40632 525943
rect 40682 519480 40738 519489
rect 40682 519415 40738 519424
rect 40590 498808 40646 498817
rect 40590 498743 40646 498752
rect 40696 479097 40724 519415
rect 40682 479088 40738 479097
rect 40682 479023 40738 479032
rect 40788 420345 40816 531655
rect 40958 531040 41014 531049
rect 40958 530975 41014 530984
rect 40866 524784 40922 524793
rect 40866 524719 40922 524728
rect 40774 420336 40830 420345
rect 40774 420271 40830 420280
rect 40880 408921 40908 524719
rect 40866 408912 40922 408921
rect 40866 408847 40922 408856
rect 40972 405657 41000 530975
rect 41064 407833 41092 545255
rect 41234 543960 41290 543969
rect 41234 543895 41290 543904
rect 41142 541240 41198 541249
rect 41142 541175 41198 541184
rect 41050 407824 41106 407833
rect 41050 407759 41106 407768
rect 40958 405648 41014 405657
rect 40958 405583 41014 405592
rect 41156 402937 41184 541175
rect 41142 402928 41198 402937
rect 41142 402863 41198 402872
rect 41248 399673 41276 543895
rect 41340 467129 41368 639911
rect 42430 549808 42486 549817
rect 42430 549743 42486 549752
rect 42154 525192 42210 525201
rect 42154 525127 42210 525136
rect 42062 523560 42118 523569
rect 42062 523495 42118 523504
rect 42076 499769 42104 523495
rect 42062 499760 42118 499769
rect 42062 499695 42118 499704
rect 42168 491201 42196 525127
rect 42246 523832 42302 523841
rect 42246 523767 42302 523776
rect 42154 491192 42210 491201
rect 42154 491127 42210 491136
rect 42260 482905 42288 523767
rect 42338 519344 42394 519353
rect 42338 519279 42394 519288
rect 42246 482896 42302 482905
rect 42246 482831 42302 482840
rect 42352 470393 42380 519279
rect 42338 470384 42394 470393
rect 42338 470319 42394 470328
rect 41326 467120 41382 467129
rect 41326 467055 41382 467064
rect 42444 426873 42472 549743
rect 42522 533488 42578 533497
rect 42522 533423 42578 533432
rect 42430 426864 42486 426873
rect 42430 426799 42486 426808
rect 42536 408377 42564 533423
rect 42628 509017 42656 642631
rect 42706 641472 42762 641481
rect 42706 641407 42762 641416
rect 42614 509008 42670 509017
rect 42614 508943 42670 508952
rect 42720 465497 42748 641407
rect 43994 635760 44050 635769
rect 43994 635695 44050 635704
rect 43534 556200 43590 556209
rect 43534 556135 43590 556144
rect 43442 537704 43498 537713
rect 43442 537639 43498 537648
rect 43350 518936 43406 518945
rect 43350 518871 43406 518880
rect 43364 476377 43392 518871
rect 43456 510513 43484 537639
rect 43442 510504 43498 510513
rect 43442 510439 43498 510448
rect 43548 497457 43576 556135
rect 43810 526144 43866 526153
rect 43810 526079 43866 526088
rect 43718 525328 43774 525337
rect 43718 525263 43774 525272
rect 43626 524920 43682 524929
rect 43626 524855 43682 524864
rect 43534 497448 43590 497457
rect 43534 497383 43590 497392
rect 43350 476368 43406 476377
rect 43350 476303 43406 476312
rect 43640 466041 43668 524855
rect 43626 466032 43682 466041
rect 43626 465967 43682 465976
rect 42706 465488 42762 465497
rect 42706 465423 42762 465432
rect 43732 459513 43760 525263
rect 43718 459504 43774 459513
rect 43718 459439 43774 459448
rect 42522 408368 42578 408377
rect 42522 408303 42578 408312
rect 43824 401849 43852 526079
rect 43902 520432 43958 520441
rect 43902 520367 43958 520376
rect 43810 401840 43866 401849
rect 43810 401775 43866 401784
rect 41234 399664 41290 399673
rect 41234 399599 41290 399608
rect 43916 395865 43944 520367
rect 44008 505209 44036 635695
rect 45006 548448 45062 548457
rect 45006 548383 45062 548392
rect 44086 547904 44142 547913
rect 44086 547839 44142 547848
rect 43994 505200 44050 505209
rect 43994 505135 44050 505144
rect 44100 402393 44128 547839
rect 44638 524648 44694 524657
rect 44638 524583 44694 524592
rect 44180 520124 44232 520130
rect 44180 520066 44232 520072
rect 44192 519489 44220 520066
rect 44178 519480 44234 519489
rect 44178 519415 44234 519424
rect 44652 504393 44680 524583
rect 44914 520024 44970 520033
rect 44914 519959 44970 519968
rect 44822 518120 44878 518129
rect 44822 518055 44878 518064
rect 44638 504384 44694 504393
rect 44638 504319 44694 504328
rect 44836 497729 44864 518055
rect 44822 497720 44878 497729
rect 44822 497655 44878 497664
rect 44928 469849 44956 519959
rect 45020 496369 45048 548383
rect 45190 537024 45246 537033
rect 45190 536959 45246 536968
rect 45098 519752 45154 519761
rect 45098 519687 45154 519696
rect 45006 496360 45062 496369
rect 45006 496295 45062 496304
rect 44914 469840 44970 469849
rect 44914 469775 44970 469784
rect 45112 460057 45140 519687
rect 45098 460048 45154 460057
rect 45098 459983 45154 459992
rect 45204 403481 45232 536959
rect 45190 403472 45246 403481
rect 45190 403407 45246 403416
rect 44086 402384 44142 402393
rect 44086 402319 44142 402328
rect 43902 395856 43958 395865
rect 43902 395791 43958 395800
rect 45296 394777 45324 643991
rect 46754 643512 46810 643521
rect 46754 643447 46810 643456
rect 45466 643240 45522 643249
rect 45466 643175 45522 643184
rect 45374 640792 45430 640801
rect 45374 640727 45430 640736
rect 45282 394768 45338 394777
rect 45282 394703 45338 394712
rect 45388 393145 45416 640727
rect 45480 393689 45508 643175
rect 46662 642152 46718 642161
rect 46662 642087 46718 642096
rect 46478 639432 46534 639441
rect 46478 639367 46534 639376
rect 46386 530088 46442 530097
rect 46386 530023 46442 530032
rect 46294 526416 46350 526425
rect 46294 526351 46350 526360
rect 46110 521928 46166 521937
rect 46110 521863 46166 521872
rect 46018 520840 46074 520849
rect 46018 520775 46074 520784
rect 45928 520192 45980 520198
rect 45928 520134 45980 520140
rect 45940 518945 45968 520134
rect 45926 518936 45982 518945
rect 45926 518871 45982 518880
rect 46032 506297 46060 520775
rect 46018 506288 46074 506297
rect 46018 506223 46074 506232
rect 46124 497865 46152 521863
rect 46110 497856 46166 497865
rect 46110 497791 46166 497800
rect 46308 417081 46336 526351
rect 46400 418169 46428 530023
rect 46492 498273 46520 639367
rect 46570 635352 46626 635361
rect 46570 635287 46626 635296
rect 46478 498264 46534 498273
rect 46478 498199 46534 498208
rect 46584 456929 46612 635287
rect 46676 458425 46704 642087
rect 46768 458969 46796 643447
rect 46754 458960 46810 458969
rect 46754 458895 46810 458904
rect 46662 458416 46718 458425
rect 46662 458351 46718 458360
rect 46570 456920 46626 456929
rect 46570 456855 46626 456864
rect 46386 418160 46442 418169
rect 46386 418095 46442 418104
rect 46294 417072 46350 417081
rect 46294 417007 46350 417016
rect 46860 394233 46888 644127
rect 48226 635080 48282 635089
rect 48226 635015 48282 635024
rect 48134 634536 48190 634545
rect 48134 634471 48190 634480
rect 48042 597408 48098 597417
rect 48042 597343 48098 597352
rect 47952 594856 48004 594862
rect 47952 594798 48004 594804
rect 47584 579692 47636 579698
rect 47584 579634 47636 579640
rect 47398 553752 47454 553761
rect 47398 553687 47454 553696
rect 47412 425241 47440 553687
rect 47596 552702 47624 579634
rect 47858 576736 47914 576745
rect 47858 576671 47914 576680
rect 47584 552696 47636 552702
rect 47584 552638 47636 552644
rect 47872 551313 47900 576671
rect 47964 558754 47992 594798
rect 47952 558748 48004 558754
rect 47952 558690 48004 558696
rect 48056 557025 48084 597343
rect 48042 557016 48098 557025
rect 48042 556951 48098 556960
rect 47950 552392 48006 552401
rect 47950 552327 48006 552336
rect 47858 551304 47914 551313
rect 47858 551239 47914 551248
rect 47766 551032 47822 551041
rect 47766 550967 47822 550976
rect 47674 539744 47730 539753
rect 47674 539679 47730 539688
rect 47582 520568 47638 520577
rect 47582 520503 47638 520512
rect 47490 517848 47546 517857
rect 47490 517783 47546 517792
rect 47504 507385 47532 517783
rect 47490 507376 47546 507385
rect 47490 507311 47546 507320
rect 47596 499225 47624 520503
rect 47582 499216 47638 499225
rect 47582 499151 47638 499160
rect 47398 425232 47454 425241
rect 47398 425167 47454 425176
rect 47688 424697 47716 539679
rect 47674 424688 47730 424697
rect 47674 424623 47730 424632
rect 47780 424153 47808 550967
rect 47766 424144 47822 424153
rect 47766 424079 47822 424088
rect 47964 423609 47992 552327
rect 48042 552256 48098 552265
rect 48042 552191 48098 552200
rect 47950 423600 48006 423609
rect 47950 423535 48006 423544
rect 48056 398041 48084 552191
rect 48148 455705 48176 634471
rect 48240 456793 48268 635015
rect 49606 618080 49662 618089
rect 49606 618015 49662 618024
rect 49422 580000 49478 580009
rect 49422 579935 49478 579944
rect 49436 555529 49464 579935
rect 49514 577824 49570 577833
rect 49514 577759 49570 577768
rect 49422 555520 49478 555529
rect 49422 555455 49478 555464
rect 49528 551993 49556 577759
rect 49514 551984 49570 551993
rect 49514 551919 49570 551928
rect 49514 549944 49570 549953
rect 49514 549879 49570 549888
rect 49422 545592 49478 545601
rect 49422 545527 49478 545536
rect 49146 544096 49202 544105
rect 49146 544031 49202 544040
rect 48870 542736 48926 542745
rect 48870 542671 48926 542680
rect 48226 456784 48282 456793
rect 48226 456719 48282 456728
rect 48134 455696 48190 455705
rect 48134 455631 48190 455640
rect 48884 422521 48912 542671
rect 49054 537296 49110 537305
rect 49054 537231 49110 537240
rect 48962 533760 49018 533769
rect 48962 533695 49018 533704
rect 48976 435577 49004 533695
rect 48962 435568 49018 435577
rect 48962 435503 49018 435512
rect 49068 434489 49096 537231
rect 49160 436665 49188 544031
rect 49238 541376 49294 541385
rect 49238 541311 49294 541320
rect 49146 436656 49202 436665
rect 49146 436591 49202 436600
rect 49054 434480 49110 434489
rect 49054 434415 49110 434424
rect 49252 432857 49280 541311
rect 49330 535936 49386 535945
rect 49330 535871 49386 535880
rect 49238 432848 49294 432857
rect 49238 432783 49294 432792
rect 48870 422512 48926 422521
rect 48870 422447 48926 422456
rect 49344 421977 49372 535871
rect 49436 431769 49464 545527
rect 49528 433401 49556 549879
rect 49620 542337 49648 618015
rect 50710 594144 50766 594153
rect 50710 594079 50766 594088
rect 50526 593056 50582 593065
rect 50526 592991 50582 593000
rect 50434 575648 50490 575657
rect 50434 575583 50490 575592
rect 50066 557696 50122 557705
rect 50066 557631 50122 557640
rect 49606 542328 49662 542337
rect 49606 542263 49662 542272
rect 49514 433392 49570 433401
rect 49514 433327 49570 433336
rect 49422 431760 49478 431769
rect 49422 431695 49478 431704
rect 50080 431225 50108 557631
rect 50448 551585 50476 575583
rect 50540 559065 50568 592991
rect 50620 590708 50672 590714
rect 50620 590650 50672 590656
rect 50526 559056 50582 559065
rect 50526 558991 50582 559000
rect 50632 556850 50660 590650
rect 50724 557433 50752 594079
rect 50710 557424 50766 557433
rect 50710 557359 50766 557368
rect 50620 556844 50672 556850
rect 50620 556786 50672 556792
rect 50434 551576 50490 551585
rect 50434 551511 50490 551520
rect 50710 548312 50766 548321
rect 50710 548247 50766 548256
rect 50526 546816 50582 546825
rect 50526 546751 50582 546760
rect 50342 538520 50398 538529
rect 50342 538455 50398 538464
rect 50250 532264 50306 532273
rect 50250 532199 50306 532208
rect 50160 520056 50212 520062
rect 50160 519998 50212 520004
rect 50172 519353 50200 519998
rect 50158 519344 50214 519353
rect 50158 519279 50214 519288
rect 50264 435033 50292 532199
rect 50356 437753 50384 538455
rect 50434 535800 50490 535809
rect 50434 535735 50490 535744
rect 50342 437744 50398 437753
rect 50342 437679 50398 437688
rect 50250 435024 50306 435033
rect 50250 434959 50306 434968
rect 50066 431216 50122 431225
rect 50066 431151 50122 431160
rect 49330 421968 49386 421977
rect 49330 421903 49386 421912
rect 50448 420889 50476 535735
rect 50540 423065 50568 546751
rect 50526 423056 50582 423065
rect 50526 422991 50582 423000
rect 50724 421433 50752 548247
rect 50816 481817 50844 646711
rect 53746 646640 53802 646649
rect 53746 646575 53802 646584
rect 52182 646504 52238 646513
rect 52182 646439 52238 646448
rect 52090 646232 52146 646241
rect 52090 646167 52146 646176
rect 50986 642016 51042 642025
rect 50986 641951 51042 641960
rect 50894 639024 50950 639033
rect 50894 638959 50950 638968
rect 50802 481808 50858 481817
rect 50802 481743 50858 481752
rect 50908 461689 50936 638959
rect 51000 462777 51028 641951
rect 51998 641200 52054 641209
rect 51998 641135 52054 641144
rect 51906 582176 51962 582185
rect 51906 582111 51962 582120
rect 51814 578912 51870 578921
rect 51814 578847 51870 578856
rect 51722 574560 51778 574569
rect 51722 574495 51778 574504
rect 51736 554033 51764 574495
rect 51722 554024 51778 554033
rect 51722 553959 51778 553968
rect 51828 552809 51856 578847
rect 51920 554169 51948 582111
rect 51906 554160 51962 554169
rect 51906 554095 51962 554104
rect 51906 553616 51962 553625
rect 51906 553551 51962 553560
rect 51814 552800 51870 552809
rect 51814 552735 51870 552744
rect 51814 546000 51870 546009
rect 51814 545935 51870 545944
rect 51722 529544 51778 529553
rect 51722 529479 51778 529488
rect 51538 528728 51594 528737
rect 51538 528663 51594 528672
rect 50986 462768 51042 462777
rect 50986 462703 51042 462712
rect 50894 461680 50950 461689
rect 50894 461615 50950 461624
rect 51552 432313 51580 528663
rect 51630 525056 51686 525065
rect 51630 524991 51686 525000
rect 51538 432304 51594 432313
rect 51538 432239 51594 432248
rect 51644 425785 51672 524991
rect 51630 425776 51686 425785
rect 51630 425711 51686 425720
rect 50710 421424 50766 421433
rect 50710 421359 50766 421368
rect 50434 420880 50490 420889
rect 50434 420815 50490 420824
rect 51736 417625 51764 529479
rect 51722 417616 51778 417625
rect 51722 417551 51778 417560
rect 51828 400217 51856 545935
rect 51920 400761 51948 553551
rect 52012 471481 52040 641135
rect 52104 473657 52132 646167
rect 52090 473648 52146 473657
rect 52090 473583 52146 473592
rect 52196 472569 52224 646439
rect 53654 646368 53710 646377
rect 53654 646303 53710 646312
rect 53470 646096 53526 646105
rect 53470 646031 53526 646040
rect 52366 643376 52422 643385
rect 52366 643311 52422 643320
rect 52274 640928 52330 640937
rect 52274 640863 52330 640872
rect 52182 472560 52238 472569
rect 52182 472495 52238 472504
rect 51998 471472 52054 471481
rect 51998 471407 52054 471416
rect 52288 461145 52316 640863
rect 52274 461136 52330 461145
rect 52274 461071 52330 461080
rect 52380 460601 52408 643311
rect 53286 636304 53342 636313
rect 53286 636239 53342 636248
rect 53194 587616 53250 587625
rect 53194 587551 53250 587560
rect 53102 573472 53158 573481
rect 53102 573407 53158 573416
rect 53116 555393 53144 573407
rect 53208 559609 53236 587551
rect 53194 559600 53250 559609
rect 53194 559535 53250 559544
rect 53102 555384 53158 555393
rect 53102 555319 53158 555328
rect 52460 552016 52512 552022
rect 52460 551958 52512 551964
rect 52472 551177 52500 551958
rect 52458 551168 52514 551177
rect 52458 551103 52514 551112
rect 53102 550896 53158 550905
rect 53102 550831 53158 550840
rect 53010 537160 53066 537169
rect 53010 537095 53066 537104
rect 52918 529952 52974 529961
rect 52918 529887 52974 529896
rect 52366 460592 52422 460601
rect 52366 460527 52422 460536
rect 52932 433945 52960 529887
rect 52918 433936 52974 433945
rect 52918 433871 52974 433880
rect 53024 412185 53052 537095
rect 53010 412176 53066 412185
rect 53010 412111 53066 412120
rect 53116 410553 53144 550831
rect 53194 549672 53250 549681
rect 53194 549607 53250 549616
rect 53102 410544 53158 410553
rect 53102 410479 53158 410488
rect 53208 409465 53236 549607
rect 53300 494193 53328 636239
rect 53380 589552 53432 589558
rect 53380 589494 53432 589500
rect 53392 558521 53420 589494
rect 53378 558512 53434 558521
rect 53378 558447 53434 558456
rect 53378 540424 53434 540433
rect 53378 540359 53434 540368
rect 53286 494184 53342 494193
rect 53286 494119 53342 494128
rect 53194 409456 53250 409465
rect 53194 409391 53250 409400
rect 51906 400752 51962 400761
rect 51906 400687 51962 400696
rect 51814 400208 51870 400217
rect 51814 400143 51870 400152
rect 48042 398032 48098 398041
rect 48042 397967 48098 397976
rect 53392 397497 53420 540359
rect 53484 478009 53512 646031
rect 53562 642832 53618 642841
rect 53562 642767 53618 642776
rect 53470 478000 53526 478009
rect 53470 477935 53526 477944
rect 53576 470937 53604 642767
rect 53668 474201 53696 646303
rect 53654 474192 53710 474201
rect 53654 474127 53710 474136
rect 53760 473113 53788 646575
rect 54298 644872 54354 644881
rect 54298 644807 54354 644816
rect 53840 635656 53892 635662
rect 53840 635598 53892 635604
rect 53852 635361 53880 635598
rect 53838 635352 53894 635361
rect 53838 635287 53894 635296
rect 53746 473104 53802 473113
rect 53746 473039 53802 473048
rect 53562 470928 53618 470937
rect 53562 470863 53618 470872
rect 54312 469305 54340 644807
rect 55034 639296 55090 639305
rect 55034 639231 55090 639240
rect 54850 636032 54906 636041
rect 54850 635967 54906 635976
rect 54666 635352 54722 635361
rect 54666 635287 54722 635296
rect 54680 601769 54708 635287
rect 54758 633448 54814 633457
rect 54758 633383 54814 633392
rect 54666 601760 54722 601769
rect 54666 601695 54722 601704
rect 54772 599593 54800 633383
rect 54864 600681 54892 635967
rect 54942 635488 54998 635497
rect 54942 635423 54998 635432
rect 54850 600672 54906 600681
rect 54850 600607 54906 600616
rect 54758 599584 54814 599593
rect 54758 599519 54814 599528
rect 54956 596329 54984 635423
rect 54942 596320 54998 596329
rect 54942 596255 54998 596264
rect 54850 591968 54906 591977
rect 54850 591903 54906 591912
rect 54758 586392 54814 586401
rect 54758 586327 54814 586336
rect 54666 585440 54722 585449
rect 54666 585375 54722 585384
rect 54482 584352 54538 584361
rect 54482 584287 54538 584296
rect 54496 555665 54524 584287
rect 54574 581088 54630 581097
rect 54574 581023 54630 581032
rect 54482 555656 54538 555665
rect 54482 555591 54538 555600
rect 54588 552945 54616 581023
rect 54680 555801 54708 585375
rect 54772 556753 54800 586327
rect 54864 559473 54892 591903
rect 54942 588704 54998 588713
rect 54942 588639 54998 588648
rect 54850 559464 54906 559473
rect 54850 559399 54906 559408
rect 54956 556889 54984 588639
rect 54942 556880 54998 556889
rect 54942 556815 54998 556824
rect 54758 556744 54814 556753
rect 54758 556679 54814 556688
rect 54666 555792 54722 555801
rect 54666 555727 54722 555736
rect 54574 552936 54630 552945
rect 54574 552871 54630 552880
rect 54758 548040 54814 548049
rect 54758 547975 54814 547984
rect 54666 542600 54722 542609
rect 54666 542535 54722 542544
rect 54574 539608 54630 539617
rect 54574 539543 54630 539552
rect 54482 535664 54538 535673
rect 54482 535599 54538 535608
rect 54390 532808 54446 532817
rect 54390 532743 54446 532752
rect 54298 469296 54354 469305
rect 54298 469231 54354 469240
rect 54404 410009 54432 532743
rect 54496 411641 54524 535599
rect 54482 411632 54538 411641
rect 54482 411567 54538 411576
rect 54390 410000 54446 410009
rect 54390 409935 54446 409944
rect 54588 404569 54616 539543
rect 54680 405113 54708 542535
rect 54772 407289 54800 547975
rect 54850 546680 54906 546689
rect 54850 546615 54906 546624
rect 54758 407280 54814 407289
rect 54758 407215 54814 407224
rect 54864 406201 54892 546615
rect 54942 543824 54998 543833
rect 54942 543759 54998 543768
rect 54850 406192 54906 406201
rect 54850 406127 54906 406136
rect 54666 405104 54722 405113
rect 54666 405039 54722 405048
rect 54574 404560 54630 404569
rect 54574 404495 54630 404504
rect 53378 397488 53434 397497
rect 53378 397423 53434 397432
rect 54956 396409 54984 543759
rect 55048 468217 55076 639231
rect 55126 583264 55182 583273
rect 55126 583199 55182 583208
rect 55140 558385 55168 583199
rect 55232 564369 55260 683130
rect 65246 647728 65302 647737
rect 65246 647663 65302 647672
rect 56506 640792 56562 640801
rect 56506 640727 56562 640736
rect 56520 640354 56548 640727
rect 56508 640348 56560 640354
rect 56508 640290 56560 640296
rect 58624 638988 58676 638994
rect 58624 638930 58676 638936
rect 55494 633312 55550 633321
rect 55494 633247 55550 633256
rect 55218 564360 55274 564369
rect 55218 564295 55274 564304
rect 55126 558376 55182 558385
rect 55126 558311 55182 558320
rect 55508 534993 55536 633247
rect 58636 632777 58664 638930
rect 63958 637256 64014 637265
rect 63958 637191 64014 637200
rect 62670 636712 62726 636721
rect 62670 636647 62726 636656
rect 62684 634916 62712 636647
rect 63972 634916 64000 637191
rect 65260 634916 65288 647663
rect 67822 639704 67878 639713
rect 67822 639639 67878 639648
rect 66534 637936 66590 637945
rect 66534 637871 66590 637880
rect 66548 634916 66576 637871
rect 67836 634916 67864 639639
rect 69110 638072 69166 638081
rect 69110 638007 69166 638016
rect 69124 634916 69152 638007
rect 71686 637392 71742 637401
rect 71686 637327 71742 637336
rect 70398 635896 70454 635905
rect 70398 635831 70454 635840
rect 70412 634916 70440 635831
rect 70582 635760 70638 635769
rect 70582 635695 70638 635704
rect 70596 634914 70624 635695
rect 71700 634916 71728 637327
rect 72988 635526 73016 703520
rect 89180 700369 89208 703520
rect 89166 700360 89222 700369
rect 105464 700330 105492 703520
rect 89166 700295 89222 700304
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 137284 700324 137336 700330
rect 137284 700266 137336 700272
rect 137296 658238 137324 700266
rect 137284 658232 137336 658238
rect 137284 658174 137336 658180
rect 103886 648136 103942 648145
rect 103886 648071 103942 648080
rect 96158 648000 96214 648009
rect 96158 647935 96214 647944
rect 91006 647864 91062 647873
rect 91006 647799 91062 647808
rect 86866 644192 86922 644201
rect 86866 644127 86922 644136
rect 80058 644056 80114 644065
rect 80058 643991 80114 644000
rect 85854 644056 85910 644065
rect 85854 643991 85910 644000
rect 80072 643278 80100 643991
rect 80702 643784 80758 643793
rect 80702 643719 80758 643728
rect 80060 643272 80112 643278
rect 80060 643214 80112 643220
rect 76838 638208 76894 638217
rect 76838 638143 76894 638152
rect 73160 637084 73212 637090
rect 73160 637026 73212 637032
rect 73172 636585 73200 637026
rect 75550 636984 75606 636993
rect 75550 636919 75606 636928
rect 73158 636576 73214 636585
rect 73158 636511 73214 636520
rect 74262 636440 74318 636449
rect 74262 636375 74318 636384
rect 72976 635520 73028 635526
rect 72976 635462 73028 635468
rect 71870 635216 71926 635225
rect 71870 635151 71926 635160
rect 72974 635216 73030 635225
rect 72974 635151 73030 635160
rect 71884 634982 71912 635151
rect 71872 634976 71924 634982
rect 71872 634918 71924 634924
rect 72988 634916 73016 635151
rect 74276 634916 74304 636375
rect 75564 634916 75592 636919
rect 75826 636848 75882 636857
rect 75826 636783 75882 636792
rect 75840 636410 75868 636783
rect 75828 636404 75880 636410
rect 75828 636346 75880 636352
rect 76852 634916 76880 638143
rect 78126 636984 78182 636993
rect 78126 636919 78182 636928
rect 78140 634916 78168 636919
rect 78588 636472 78640 636478
rect 78588 636414 78640 636420
rect 78600 636313 78628 636414
rect 78586 636304 78642 636313
rect 78586 636239 78642 636248
rect 79414 635760 79470 635769
rect 79324 635724 79376 635730
rect 79414 635695 79470 635704
rect 79324 635666 79376 635672
rect 79336 635089 79364 635666
rect 79322 635080 79378 635089
rect 79322 635015 79378 635024
rect 79428 634916 79456 635695
rect 80716 634916 80744 643719
rect 84566 642424 84622 642433
rect 84566 642359 84622 642368
rect 82818 639976 82874 639985
rect 82818 639911 82874 639920
rect 81438 639296 81494 639305
rect 82832 639266 82860 639911
rect 83278 639296 83334 639305
rect 81438 639231 81494 639240
rect 82820 639260 82872 639266
rect 81452 639198 81480 639231
rect 83278 639231 83334 639240
rect 82820 639202 82872 639208
rect 81440 639192 81492 639198
rect 81440 639134 81492 639140
rect 81990 639160 82046 639169
rect 81990 639095 82046 639104
rect 82004 634916 82032 639095
rect 83292 634916 83320 639231
rect 84580 634916 84608 642359
rect 85488 642116 85540 642122
rect 85488 642058 85540 642064
rect 85500 641753 85528 642058
rect 85486 641744 85542 641753
rect 85486 641679 85542 641688
rect 85868 634916 85896 643991
rect 86880 643346 86908 644127
rect 88430 643920 88486 643929
rect 88430 643855 88486 643864
rect 86868 643340 86920 643346
rect 86868 643282 86920 643288
rect 87142 638616 87198 638625
rect 87142 638551 87198 638560
rect 87156 634916 87184 638551
rect 88444 634916 88472 643855
rect 88984 643408 89036 643414
rect 88984 643350 89036 643356
rect 88996 643249 89024 643350
rect 88982 643240 89038 643249
rect 88982 643175 89038 643184
rect 89718 638344 89774 638353
rect 89718 638279 89774 638288
rect 89732 634916 89760 638279
rect 91020 634916 91048 647799
rect 92478 642560 92534 642569
rect 92478 642495 92534 642504
rect 93582 642560 93638 642569
rect 93582 642495 93638 642504
rect 92492 642190 92520 642495
rect 92480 642184 92532 642190
rect 92480 642126 92532 642132
rect 91098 641200 91154 641209
rect 91098 641135 91154 641144
rect 92294 641200 92350 641209
rect 92294 641135 92350 641144
rect 91112 640762 91140 641135
rect 91100 640756 91152 640762
rect 91100 640698 91152 640704
rect 92308 634916 92336 641135
rect 93596 634916 93624 642495
rect 94870 639976 94926 639985
rect 94870 639911 94926 639920
rect 94884 634916 94912 639911
rect 95146 639840 95202 639849
rect 95146 639775 95202 639784
rect 95160 639402 95188 639775
rect 95148 639396 95200 639402
rect 95148 639338 95200 639344
rect 96172 634916 96200 647935
rect 102598 645416 102654 645425
rect 102598 645351 102654 645360
rect 98734 645280 98790 645289
rect 98734 645215 98790 645224
rect 97828 635718 98132 635746
rect 97828 634930 97856 635718
rect 98104 635633 98132 635718
rect 97906 635624 97962 635633
rect 97906 635559 97962 635568
rect 98090 635624 98146 635633
rect 98090 635559 98146 635568
rect 97920 635322 97948 635559
rect 97908 635316 97960 635322
rect 97908 635258 97960 635264
rect 70584 634908 70636 634914
rect 97474 634902 97856 634930
rect 98748 634916 98776 645215
rect 102138 645144 102194 645153
rect 102138 645079 102194 645088
rect 102152 644706 102180 645079
rect 102140 644700 102192 644706
rect 102140 644642 102192 644648
rect 99378 637528 99434 637537
rect 99378 637463 99434 637472
rect 99392 636750 99420 637463
rect 100022 637120 100078 637129
rect 100022 637055 100078 637064
rect 99380 636744 99432 636750
rect 99380 636686 99432 636692
rect 100036 634916 100064 637055
rect 101312 636880 101364 636886
rect 101312 636822 101364 636828
rect 101324 634916 101352 636822
rect 102612 634916 102640 645351
rect 103900 634916 103928 648071
rect 106186 645552 106242 645561
rect 106186 645487 106242 645496
rect 105174 645144 105230 645153
rect 105174 645079 105230 645088
rect 105188 634916 105216 645079
rect 106200 644842 106228 645487
rect 106188 644836 106240 644842
rect 106188 644778 106240 644784
rect 125598 640112 125654 640121
rect 125598 640047 125654 640056
rect 121918 639568 121974 639577
rect 121918 639503 121974 639512
rect 109038 638752 109094 638761
rect 109038 638687 109094 638696
rect 107750 638480 107806 638489
rect 107750 638415 107806 638424
rect 106464 636540 106516 636546
rect 106464 636482 106516 636488
rect 106476 634916 106504 636482
rect 107764 634916 107792 638415
rect 108304 637968 108356 637974
rect 108304 637910 108356 637916
rect 108316 637809 108344 637910
rect 108302 637800 108358 637809
rect 108302 637735 108358 637744
rect 109052 637634 109080 638687
rect 110328 638036 110380 638042
rect 110328 637978 110380 637984
rect 109498 637664 109554 637673
rect 109040 637628 109092 637634
rect 109498 637599 109554 637608
rect 109040 637570 109092 637576
rect 109512 634930 109540 637599
rect 109066 634902 109540 634930
rect 110340 634916 110368 637978
rect 115480 637696 115532 637702
rect 115480 637638 115532 637644
rect 114192 636676 114244 636682
rect 114192 636618 114244 636624
rect 111616 636608 111668 636614
rect 111616 636550 111668 636556
rect 111628 634916 111656 636550
rect 112904 635520 112956 635526
rect 112904 635462 112956 635468
rect 112916 634916 112944 635462
rect 114204 634916 114232 636618
rect 115492 634916 115520 637638
rect 121366 635760 121422 635769
rect 121366 635695 121422 635704
rect 119986 635624 120042 635633
rect 119986 635559 120042 635568
rect 120000 635458 120028 635559
rect 119988 635452 120040 635458
rect 119988 635394 120040 635400
rect 121380 635390 121408 635695
rect 121368 635384 121420 635390
rect 121368 635326 121420 635332
rect 121090 635080 121146 635089
rect 121090 635015 121146 635024
rect 119342 634944 119398 634953
rect 121104 634930 121132 635015
rect 120658 634902 121132 634930
rect 121932 634916 121960 639503
rect 122748 639464 122800 639470
rect 122748 639406 122800 639412
rect 122760 639033 122788 639406
rect 125612 639130 125640 640047
rect 125600 639124 125652 639130
rect 125600 639066 125652 639072
rect 122746 639024 122802 639033
rect 122746 638959 122802 638968
rect 125782 639024 125838 639033
rect 125782 638959 125838 638968
rect 123484 638376 123536 638382
rect 123484 638318 123536 638324
rect 123206 637800 123262 637809
rect 123206 637735 123262 637744
rect 123220 634916 123248 637735
rect 123496 637673 123524 638318
rect 123482 637664 123538 637673
rect 123482 637599 123538 637608
rect 124218 637120 124274 637129
rect 124218 637055 124274 637064
rect 124232 636818 124260 637055
rect 124220 636812 124272 636818
rect 124220 636754 124272 636760
rect 124494 636304 124550 636313
rect 124494 636239 124550 636248
rect 124508 634916 124536 636239
rect 125796 634916 125824 638959
rect 129738 638480 129794 638489
rect 129738 638415 129740 638424
rect 129792 638415 129794 638424
rect 130934 638480 130990 638489
rect 130934 638415 130990 638424
rect 129740 638386 129792 638392
rect 129648 636268 129700 636274
rect 129648 636210 129700 636216
rect 129660 634916 129688 636210
rect 119342 634879 119398 634888
rect 70584 634850 70636 634856
rect 127070 634672 127126 634681
rect 127070 634607 127126 634616
rect 130948 634545 130976 638415
rect 136086 637392 136142 637401
rect 136086 637327 136142 637336
rect 131118 636984 131174 636993
rect 131118 636919 131174 636928
rect 131132 636342 131160 636919
rect 135996 636880 136048 636886
rect 134614 636848 134670 636857
rect 135996 636822 136048 636828
rect 134614 636783 134670 636792
rect 135904 636812 135956 636818
rect 132222 636576 132278 636585
rect 132222 636511 132278 636520
rect 131120 636336 131172 636342
rect 131120 636278 131172 636284
rect 132236 634916 132264 636511
rect 134628 634814 134656 636783
rect 135904 636754 135956 636760
rect 134708 636336 134760 636342
rect 134708 636278 134760 636284
rect 135258 636304 135314 636313
rect 134536 634786 134656 634814
rect 129830 634536 129886 634545
rect 129830 634471 129886 634480
rect 130934 634536 130990 634545
rect 130934 634471 130990 634480
rect 129844 634438 129872 634471
rect 129832 634432 129884 634438
rect 118054 634400 118110 634409
rect 129832 634374 129884 634380
rect 118054 634335 118110 634344
rect 116757 634208 116766 634264
rect 116822 634208 116831 634264
rect 128349 634208 128358 634264
rect 128414 634208 128423 634264
rect 55586 632768 55642 632777
rect 55586 632703 55588 632712
rect 55640 632703 55642 632712
rect 58622 632768 58678 632777
rect 58622 632703 58678 632712
rect 55588 632674 55640 632680
rect 55600 632097 55628 632674
rect 55586 632088 55642 632097
rect 55586 632023 55642 632032
rect 56322 629912 56378 629921
rect 56322 629847 56378 629856
rect 56138 609376 56194 609385
rect 56138 609311 56194 609320
rect 55954 570208 56010 570217
rect 55954 570143 56010 570152
rect 55678 563544 55734 563553
rect 55678 563479 55734 563488
rect 55692 554577 55720 563479
rect 55770 558920 55826 558929
rect 55770 558855 55826 558864
rect 55678 554568 55734 554577
rect 55678 554503 55734 554512
rect 55494 534984 55550 534993
rect 55494 534919 55550 534928
rect 55678 529816 55734 529825
rect 55678 529751 55734 529760
rect 55128 520260 55180 520266
rect 55128 520202 55180 520208
rect 55140 519625 55168 520202
rect 55126 519616 55182 519625
rect 55126 519551 55182 519560
rect 55128 519036 55180 519042
rect 55128 518978 55180 518984
rect 55140 518945 55168 518978
rect 55126 518936 55182 518945
rect 55126 518871 55182 518880
rect 55034 468208 55090 468217
rect 55034 468143 55090 468152
rect 54942 396400 54998 396409
rect 54942 396335 54998 396344
rect 46846 394224 46902 394233
rect 46846 394159 46902 394168
rect 45466 393680 45522 393689
rect 45466 393615 45522 393624
rect 45374 393136 45430 393145
rect 45374 393071 45430 393080
rect 55692 387161 55720 529751
rect 55784 524482 55812 558855
rect 55864 557456 55916 557462
rect 55864 557398 55916 557404
rect 55876 556617 55904 557398
rect 55862 556608 55918 556617
rect 55862 556543 55918 556552
rect 55968 552673 55996 570143
rect 56046 568032 56102 568041
rect 56046 567967 56102 567976
rect 55954 552664 56010 552673
rect 55954 552599 56010 552608
rect 56060 547505 56088 567967
rect 56046 547496 56102 547505
rect 56046 547431 56102 547440
rect 56152 539209 56180 609311
rect 56230 598496 56286 598505
rect 56230 598431 56286 598440
rect 56244 557297 56272 598431
rect 56230 557288 56286 557297
rect 56230 557223 56286 557232
rect 56230 554840 56286 554849
rect 56230 554775 56286 554784
rect 56138 539200 56194 539209
rect 56138 539135 56194 539144
rect 55954 538384 56010 538393
rect 55954 538319 56010 538328
rect 55862 532944 55918 532953
rect 55862 532879 55918 532888
rect 55772 524476 55824 524482
rect 55772 524418 55824 524424
rect 55770 523016 55826 523025
rect 55770 522951 55826 522960
rect 55784 467673 55812 522951
rect 55770 467664 55826 467673
rect 55770 467599 55826 467608
rect 55876 419257 55904 532879
rect 55862 419248 55918 419257
rect 55862 419183 55918 419192
rect 55968 412729 55996 538319
rect 56046 534168 56102 534177
rect 56046 534103 56102 534112
rect 55954 412720 56010 412729
rect 55954 412655 56010 412664
rect 56060 406745 56088 534103
rect 56140 519716 56192 519722
rect 56140 519658 56192 519664
rect 56046 406736 56102 406745
rect 56046 406671 56102 406680
rect 56152 387598 56180 519658
rect 56244 419801 56272 554775
rect 56336 542065 56364 629847
rect 56414 628824 56470 628833
rect 56414 628759 56470 628768
rect 56322 542056 56378 542065
rect 56322 541991 56378 542000
rect 56428 540841 56456 628759
rect 59174 625696 59230 625705
rect 59174 625631 59230 625640
rect 57610 624608 57666 624617
rect 57610 624543 57666 624552
rect 57518 615904 57574 615913
rect 57518 615839 57574 615848
rect 57334 612640 57390 612649
rect 57334 612575 57390 612584
rect 57242 607200 57298 607209
rect 57242 607135 57298 607144
rect 57058 605024 57114 605033
rect 57058 604959 57114 604968
rect 56966 595232 57022 595241
rect 56966 595167 57022 595176
rect 56980 594862 57008 595167
rect 56968 594856 57020 594862
rect 56968 594798 57020 594804
rect 56966 590880 57022 590889
rect 56966 590815 57022 590824
rect 56980 590714 57008 590815
rect 56968 590708 57020 590714
rect 56968 590650 57020 590656
rect 56966 589792 57022 589801
rect 56966 589727 57022 589736
rect 56980 589558 57008 589727
rect 56968 589552 57020 589558
rect 56968 589494 57020 589500
rect 56968 563236 57020 563242
rect 56968 563178 57020 563184
rect 56508 558816 56560 558822
rect 56508 558758 56560 558764
rect 56520 557705 56548 558758
rect 56980 558634 57008 563178
rect 57072 559881 57100 604959
rect 57150 602848 57206 602857
rect 57150 602783 57206 602792
rect 57058 559872 57114 559881
rect 57058 559807 57114 559816
rect 57058 558648 57114 558657
rect 56980 558606 57058 558634
rect 57058 558583 57114 558592
rect 56506 557696 56562 557705
rect 56506 557631 56562 557640
rect 56508 557524 56560 557530
rect 56508 557466 56560 557472
rect 56520 556209 56548 557466
rect 56506 556200 56562 556209
rect 56506 556135 56562 556144
rect 57164 555937 57192 602783
rect 57256 560017 57284 607135
rect 57348 560318 57376 612575
rect 57426 603936 57482 603945
rect 57426 603871 57482 603880
rect 57336 560312 57388 560318
rect 57336 560254 57388 560260
rect 57336 560176 57388 560182
rect 57336 560118 57388 560124
rect 57242 560008 57298 560017
rect 57242 559943 57298 559952
rect 57348 559337 57376 560118
rect 57334 559328 57390 559337
rect 57334 559263 57390 559272
rect 57150 555928 57206 555937
rect 57150 555863 57206 555872
rect 57152 555484 57204 555490
rect 57152 555426 57204 555432
rect 56414 540832 56470 540841
rect 56414 540767 56470 540776
rect 56414 538248 56470 538257
rect 56414 538183 56470 538192
rect 56322 535528 56378 535537
rect 56322 535463 56378 535472
rect 56230 419792 56286 419801
rect 56230 419727 56286 419736
rect 56336 401305 56364 535463
rect 56428 404025 56456 538183
rect 56874 528592 56930 528601
rect 56874 528527 56930 528536
rect 56508 522980 56560 522986
rect 56508 522922 56560 522928
rect 56520 522617 56548 522922
rect 56506 522608 56562 522617
rect 56506 522543 56562 522552
rect 56508 519580 56560 519586
rect 56508 519522 56560 519528
rect 56520 518974 56548 519522
rect 56508 518968 56560 518974
rect 56508 518910 56560 518916
rect 56520 516186 56548 518910
rect 56784 518220 56836 518226
rect 56784 518162 56836 518168
rect 56508 516180 56560 516186
rect 56508 516122 56560 516128
rect 56796 499610 56824 518162
rect 56888 515545 56916 528527
rect 56966 524240 57022 524249
rect 56966 524175 57022 524184
rect 56874 515536 56930 515545
rect 56874 515471 56930 515480
rect 56980 514457 57008 524175
rect 56966 514448 57022 514457
rect 56966 514383 57022 514392
rect 57164 513369 57192 555426
rect 57440 547233 57468 603871
rect 57532 563242 57560 615839
rect 57520 563236 57572 563242
rect 57520 563178 57572 563184
rect 57624 563122 57652 624543
rect 59082 622432 59138 622441
rect 59082 622367 59138 622376
rect 57794 621344 57850 621353
rect 57794 621279 57850 621288
rect 57702 613728 57758 613737
rect 57702 613663 57758 613672
rect 57532 563094 57652 563122
rect 57532 560289 57560 563094
rect 57518 560280 57574 560289
rect 57518 560215 57574 560224
rect 57612 560244 57664 560250
rect 57612 560186 57664 560192
rect 57520 560108 57572 560114
rect 57520 560050 57572 560056
rect 57532 559201 57560 560050
rect 57624 559745 57652 560186
rect 57610 559736 57666 559745
rect 57610 559671 57666 559680
rect 57518 559192 57574 559201
rect 57518 559127 57574 559136
rect 57612 558884 57664 558890
rect 57612 558826 57664 558832
rect 57624 557977 57652 558826
rect 57610 557968 57666 557977
rect 57610 557903 57666 557912
rect 57716 555218 57744 613663
rect 57704 555212 57756 555218
rect 57704 555154 57756 555160
rect 57808 555098 57836 621279
rect 58438 620256 58494 620265
rect 58438 620191 58494 620200
rect 57886 616992 57942 617001
rect 57886 616927 57942 616936
rect 57532 555070 57836 555098
rect 57532 550497 57560 555070
rect 57704 555008 57756 555014
rect 57610 554976 57666 554985
rect 57704 554950 57756 554956
rect 57610 554911 57666 554920
rect 57518 550488 57574 550497
rect 57518 550423 57574 550432
rect 57426 547224 57482 547233
rect 57426 547159 57482 547168
rect 57334 546952 57390 546961
rect 57334 546887 57390 546896
rect 57244 516180 57296 516186
rect 57244 516122 57296 516128
rect 57150 513360 57206 513369
rect 57150 513295 57206 513304
rect 56968 512032 57020 512038
rect 56968 511974 57020 511980
rect 56876 499724 56928 499730
rect 56876 499666 56928 499672
rect 56888 499610 56916 499666
rect 56796 499582 56916 499610
rect 56414 404016 56470 404025
rect 56414 403951 56470 403960
rect 56322 401296 56378 401305
rect 56322 401231 56378 401240
rect 56140 387592 56192 387598
rect 56140 387534 56192 387540
rect 55678 387152 55734 387161
rect 55678 387087 55734 387096
rect 56980 345710 57008 511974
rect 57152 499724 57204 499730
rect 57152 499666 57204 499672
rect 57058 496360 57114 496369
rect 57058 496295 57114 496304
rect 57072 490618 57100 496295
rect 57164 495553 57192 499666
rect 57150 495544 57206 495553
rect 57150 495479 57206 495488
rect 57150 492688 57206 492697
rect 57150 492623 57206 492632
rect 57060 490612 57112 490618
rect 57060 490554 57112 490560
rect 57164 480185 57192 492623
rect 57150 480176 57206 480185
rect 57150 480111 57206 480120
rect 57256 387734 57284 516122
rect 57348 516089 57376 546887
rect 57426 529136 57482 529145
rect 57426 529071 57482 529080
rect 57440 517177 57468 529071
rect 57518 527640 57574 527649
rect 57518 527575 57574 527584
rect 57426 517168 57482 517177
rect 57426 517103 57482 517112
rect 57428 517064 57480 517070
rect 57428 517006 57480 517012
rect 57334 516080 57390 516089
rect 57334 516015 57390 516024
rect 57440 505094 57468 517006
rect 57532 513913 57560 527575
rect 57518 513904 57574 513913
rect 57518 513839 57574 513848
rect 57624 512825 57652 554911
rect 57716 543697 57744 554950
rect 57796 553308 57848 553314
rect 57796 553250 57848 553256
rect 57808 552537 57836 553250
rect 57794 552528 57850 552537
rect 57794 552463 57850 552472
rect 57702 543688 57758 543697
rect 57702 543623 57758 543632
rect 57900 539481 57928 616927
rect 58346 565856 58402 565865
rect 58346 565791 58402 565800
rect 58072 560312 58124 560318
rect 58072 560254 58124 560260
rect 58084 559337 58112 560254
rect 58070 559328 58126 559337
rect 58070 559263 58126 559272
rect 58360 549137 58388 565791
rect 58346 549128 58402 549137
rect 58346 549063 58402 549072
rect 58452 543425 58480 620191
rect 58990 619168 59046 619177
rect 58990 619103 59046 619112
rect 58898 614816 58954 614825
rect 58898 614751 58954 614760
rect 58806 610464 58862 610473
rect 58806 610399 58862 610408
rect 58714 608288 58770 608297
rect 58714 608223 58770 608232
rect 58622 571296 58678 571305
rect 58622 571231 58678 571240
rect 58636 554810 58664 571231
rect 58624 554804 58676 554810
rect 58624 554746 58676 554752
rect 58728 554690 58756 608223
rect 58544 554662 58756 554690
rect 58544 551857 58572 554662
rect 58624 554600 58676 554606
rect 58624 554542 58676 554548
rect 58530 551848 58586 551857
rect 58530 551783 58586 551792
rect 58438 543416 58494 543425
rect 58438 543351 58494 543360
rect 58636 541521 58664 554542
rect 58716 552084 58768 552090
rect 58716 552026 58768 552032
rect 58728 548350 58756 552026
rect 58716 548344 58768 548350
rect 58716 548286 58768 548292
rect 58820 547874 58848 610399
rect 58728 547846 58848 547874
rect 58728 544785 58756 547846
rect 58714 544776 58770 544785
rect 58714 544711 58770 544720
rect 58622 541512 58678 541521
rect 58622 541447 58678 541456
rect 57886 539472 57942 539481
rect 57886 539407 57942 539416
rect 58912 530505 58940 614751
rect 59004 532545 59032 619103
rect 59096 536489 59124 622367
rect 59082 536480 59138 536489
rect 59082 536415 59138 536424
rect 59188 536058 59216 625631
rect 59818 623520 59874 623529
rect 59818 623455 59874 623464
rect 59832 615494 59860 623455
rect 59832 615466 59952 615494
rect 59726 611552 59782 611561
rect 59726 611487 59782 611496
rect 59542 569120 59598 569129
rect 59542 569055 59598 569064
rect 59266 566808 59322 566817
rect 59266 566743 59322 566752
rect 59280 554713 59308 566743
rect 59556 557161 59584 569055
rect 59636 558204 59688 558210
rect 59636 558146 59688 558152
rect 59542 557152 59598 557161
rect 59542 557087 59598 557096
rect 59266 554704 59322 554713
rect 59266 554639 59322 554648
rect 59268 551948 59320 551954
rect 59268 551890 59320 551896
rect 59280 551041 59308 551890
rect 59266 551032 59322 551041
rect 59266 550967 59322 550976
rect 59268 549024 59320 549030
rect 59268 548966 59320 548972
rect 59280 548457 59308 548966
rect 59266 548448 59322 548457
rect 59266 548383 59322 548392
rect 59268 548344 59320 548350
rect 59268 548286 59320 548292
rect 59096 536030 59216 536058
rect 59096 533905 59124 536030
rect 59176 533928 59228 533934
rect 59082 533896 59138 533905
rect 59176 533870 59228 533876
rect 59082 533831 59138 533840
rect 59188 533633 59216 533870
rect 59174 533624 59230 533633
rect 59174 533559 59230 533568
rect 58990 532536 59046 532545
rect 58990 532471 59046 532480
rect 59176 531072 59228 531078
rect 59176 531014 59228 531020
rect 58898 530496 58954 530505
rect 58898 530431 58954 530440
rect 59188 530369 59216 531014
rect 59174 530360 59230 530369
rect 59174 530295 59230 530304
rect 59176 529848 59228 529854
rect 59176 529790 59228 529796
rect 59082 529272 59138 529281
rect 59082 529207 59138 529216
rect 57794 528864 57850 528873
rect 57794 528799 57850 528808
rect 57702 520024 57758 520033
rect 57702 519959 57704 519968
rect 57756 519959 57758 519968
rect 57704 519930 57756 519936
rect 57704 517608 57756 517614
rect 57704 517550 57756 517556
rect 57610 512816 57666 512825
rect 57610 512751 57666 512760
rect 57518 506424 57574 506433
rect 57518 506359 57574 506368
rect 57348 505066 57468 505094
rect 57348 504529 57376 505066
rect 57334 504520 57390 504529
rect 57334 504455 57390 504464
rect 57532 500313 57560 506359
rect 57610 504384 57666 504393
rect 57610 504319 57666 504328
rect 57518 500304 57574 500313
rect 57518 500239 57574 500248
rect 57624 499361 57652 504319
rect 57716 500954 57744 517550
rect 57808 516633 57836 528799
rect 57886 527504 57942 527513
rect 57886 527439 57942 527448
rect 57794 516624 57850 516633
rect 57794 516559 57850 516568
rect 57900 512281 57928 527439
rect 58624 524476 58676 524482
rect 58624 524418 58676 524424
rect 57978 523832 58034 523841
rect 57978 523767 58034 523776
rect 57886 512272 57942 512281
rect 57886 512207 57942 512216
rect 57794 509960 57850 509969
rect 57794 509895 57850 509904
rect 57704 500948 57756 500954
rect 57704 500890 57756 500896
rect 57610 499352 57666 499361
rect 57610 499287 57666 499296
rect 57518 499216 57574 499225
rect 57518 499151 57574 499160
rect 57426 497856 57482 497865
rect 57426 497791 57482 497800
rect 57334 497720 57390 497729
rect 57334 497655 57390 497664
rect 57348 491609 57376 497655
rect 57440 493241 57468 497791
rect 57532 497049 57560 499151
rect 57610 498944 57666 498953
rect 57610 498879 57666 498888
rect 57624 497593 57652 498879
rect 57702 498808 57758 498817
rect 57702 498743 57758 498752
rect 57610 497584 57666 497593
rect 57610 497519 57666 497528
rect 57610 497448 57666 497457
rect 57610 497383 57666 497392
rect 57518 497040 57574 497049
rect 57518 496975 57574 496984
rect 57624 494329 57652 497383
rect 57716 495417 57744 498743
rect 57702 495408 57758 495417
rect 57702 495343 57758 495352
rect 57610 494320 57666 494329
rect 57610 494255 57666 494264
rect 57518 494184 57574 494193
rect 57518 494119 57574 494128
rect 57426 493232 57482 493241
rect 57426 493167 57482 493176
rect 57532 493082 57560 494119
rect 57440 493054 57560 493082
rect 57334 491600 57390 491609
rect 57334 491535 57390 491544
rect 57336 490612 57388 490618
rect 57336 490554 57388 490560
rect 57348 392601 57376 490554
rect 57440 468761 57468 493054
rect 57702 492960 57758 492969
rect 57702 492895 57758 492904
rect 57518 491328 57574 491337
rect 57518 491263 57574 491272
rect 57532 475289 57560 491263
rect 57610 489832 57666 489841
rect 57610 489767 57666 489776
rect 57518 475280 57574 475289
rect 57518 475215 57574 475224
rect 57426 468752 57482 468761
rect 57426 468687 57482 468696
rect 57624 463865 57652 489767
rect 57610 463856 57666 463865
rect 57610 463791 57666 463800
rect 57716 430681 57744 492895
rect 57702 430672 57758 430681
rect 57702 430607 57758 430616
rect 57334 392592 57390 392601
rect 57334 392527 57390 392536
rect 57244 387728 57296 387734
rect 57244 387670 57296 387676
rect 57808 386481 57836 509895
rect 57886 509144 57942 509153
rect 57886 509079 57942 509088
rect 57900 503033 57928 509079
rect 57886 503024 57942 503033
rect 57886 502959 57942 502968
rect 57992 491337 58020 523767
rect 58440 519648 58492 519654
rect 58440 519590 58492 519596
rect 58070 517576 58126 517585
rect 58070 517511 58126 517520
rect 57978 491328 58034 491337
rect 57978 491263 58034 491272
rect 58084 489841 58112 517511
rect 58452 512038 58480 519590
rect 58530 518800 58586 518809
rect 58530 518735 58586 518744
rect 58440 512032 58492 512038
rect 58440 511974 58492 511980
rect 58544 506433 58572 518735
rect 58530 506424 58586 506433
rect 58530 506359 58586 506368
rect 58070 489832 58126 489841
rect 58070 489767 58126 489776
rect 57794 386472 57850 386481
rect 57794 386407 57850 386416
rect 56968 345704 57020 345710
rect 56968 345646 57020 345652
rect 58636 341698 58664 524418
rect 59096 523682 59124 529207
rect 59188 528737 59216 529790
rect 59174 528728 59230 528737
rect 59174 528663 59230 528672
rect 59176 524408 59228 524414
rect 59176 524350 59228 524356
rect 59188 523977 59216 524350
rect 59174 523968 59230 523977
rect 59174 523903 59230 523912
rect 59096 523654 59216 523682
rect 59082 521656 59138 521665
rect 59082 521591 59138 521600
rect 58808 521008 58860 521014
rect 58808 520950 58860 520956
rect 58716 519036 58768 519042
rect 58716 518978 58768 518984
rect 58728 387666 58756 518978
rect 58820 517562 58848 520950
rect 58900 518900 58952 518906
rect 58900 518842 58952 518848
rect 58912 517857 58940 518842
rect 58992 518832 59044 518838
rect 58992 518774 59044 518780
rect 59004 517993 59032 518774
rect 58990 517984 59046 517993
rect 58990 517919 59046 517928
rect 58992 517880 59044 517886
rect 58898 517848 58954 517857
rect 58992 517822 59044 517828
rect 58898 517783 58954 517792
rect 58820 517534 58940 517562
rect 58912 511737 58940 517534
rect 58898 511728 58954 511737
rect 58898 511663 58954 511672
rect 59004 509153 59032 517822
rect 58990 509144 59046 509153
rect 58990 509079 59046 509088
rect 58990 504520 59046 504529
rect 58990 504455 59046 504464
rect 58808 500948 58860 500954
rect 58808 500890 58860 500896
rect 58820 389910 58848 500890
rect 58898 495544 58954 495553
rect 58898 495479 58954 495488
rect 58912 429049 58940 495479
rect 59004 492697 59032 504455
rect 58990 492688 59046 492697
rect 58990 492623 59046 492632
rect 59096 466585 59124 521591
rect 59188 502489 59216 523654
rect 59174 502480 59230 502489
rect 59174 502415 59230 502424
rect 59174 489832 59230 489841
rect 59174 489767 59230 489776
rect 59082 466576 59138 466585
rect 59082 466511 59138 466520
rect 58898 429040 58954 429049
rect 58898 428975 58954 428984
rect 58808 389904 58860 389910
rect 58808 389846 58860 389852
rect 59188 389201 59216 489767
rect 59174 389192 59230 389201
rect 59174 389127 59230 389136
rect 58716 387660 58768 387666
rect 58716 387602 58768 387608
rect 59280 387297 59308 548286
rect 59542 530768 59598 530777
rect 59542 530703 59598 530712
rect 59452 529916 59504 529922
rect 59452 529858 59504 529864
rect 59464 529145 59492 529858
rect 59450 529136 59506 529145
rect 59450 529071 59506 529080
rect 59556 523025 59584 530703
rect 59542 523016 59598 523025
rect 59542 522951 59598 522960
rect 59544 518288 59596 518294
rect 59544 518230 59596 518236
rect 59556 509969 59584 518230
rect 59542 509960 59598 509969
rect 59542 509895 59598 509904
rect 59648 492969 59676 558146
rect 59740 538121 59768 611487
rect 59818 606112 59874 606121
rect 59818 606047 59874 606056
rect 59726 538112 59782 538121
rect 59726 538047 59782 538056
rect 59832 531865 59860 606047
rect 59818 531856 59874 531865
rect 59818 531791 59874 531800
rect 59924 531706 59952 615466
rect 98736 560652 98788 560658
rect 98736 560594 98788 560600
rect 60738 560416 60794 560425
rect 60738 560351 60794 560360
rect 60002 560280 60058 560289
rect 60002 560215 60058 560224
rect 59832 531678 59952 531706
rect 59832 529802 59860 531678
rect 59912 531276 59964 531282
rect 59912 531218 59964 531224
rect 59924 529961 59952 531218
rect 59910 529952 59966 529961
rect 59910 529887 59966 529896
rect 59910 529816 59966 529825
rect 59832 529774 59910 529802
rect 59910 529751 59966 529760
rect 59912 522844 59964 522850
rect 59912 522786 59964 522792
rect 59924 522073 59952 522786
rect 59910 522064 59966 522073
rect 59910 521999 59966 522008
rect 59634 492960 59690 492969
rect 59634 492895 59690 492904
rect 59450 492688 59506 492697
rect 59450 492623 59506 492632
rect 59464 489841 59492 492623
rect 59450 489832 59506 489841
rect 59450 489767 59506 489776
rect 60016 402974 60044 560215
rect 60464 558408 60516 558414
rect 60464 558350 60516 558356
rect 60096 557388 60148 557394
rect 60096 557330 60148 557336
rect 60108 556345 60136 557330
rect 60094 556336 60150 556345
rect 60094 556271 60150 556280
rect 60096 551336 60148 551342
rect 60096 551278 60148 551284
rect 60108 430409 60136 551278
rect 60476 547874 60504 558350
rect 60556 558340 60608 558346
rect 60556 558282 60608 558288
rect 60568 557534 60596 558282
rect 60568 557506 60688 557534
rect 60556 552696 60608 552702
rect 60556 552638 60608 552644
rect 60384 547846 60504 547874
rect 60188 546440 60240 546446
rect 60188 546382 60240 546388
rect 60200 545737 60228 546382
rect 60384 545873 60412 547846
rect 60370 545864 60426 545873
rect 60370 545799 60426 545808
rect 60186 545728 60242 545737
rect 60186 545663 60242 545672
rect 60186 537432 60242 537441
rect 60186 537367 60242 537376
rect 60200 436393 60228 537367
rect 60278 534304 60334 534313
rect 60278 534239 60334 534248
rect 60186 436384 60242 436393
rect 60186 436319 60242 436328
rect 60094 430400 60150 430409
rect 60094 430335 60150 430344
rect 60292 429865 60320 534239
rect 60372 527876 60424 527882
rect 60372 527818 60424 527824
rect 60384 527202 60412 527818
rect 60372 527196 60424 527202
rect 60372 527138 60424 527144
rect 60384 518894 60412 527138
rect 60384 518866 60504 518894
rect 60372 517540 60424 517546
rect 60372 517482 60424 517488
rect 60278 429856 60334 429865
rect 60278 429791 60334 429800
rect 60016 402946 60320 402974
rect 59266 387288 59322 387297
rect 60292 387258 60320 402946
rect 60384 389842 60412 517482
rect 60372 389836 60424 389842
rect 60372 389778 60424 389784
rect 60476 387433 60504 518866
rect 60568 387530 60596 552638
rect 60660 387705 60688 557506
rect 60752 535650 60780 560351
rect 96526 560280 96582 560289
rect 96526 560215 96582 560224
rect 63774 560144 63830 560153
rect 60832 538212 60884 538218
rect 60832 538154 60884 538160
rect 60844 537713 60872 538154
rect 60830 537704 60886 537713
rect 60830 537639 60886 537648
rect 61488 537577 61516 560116
rect 61566 538792 61622 538801
rect 61566 538727 61622 538736
rect 61474 537568 61530 537577
rect 61474 537503 61530 537512
rect 60752 535622 60872 535650
rect 60740 534064 60792 534070
rect 60740 534006 60792 534012
rect 60752 533769 60780 534006
rect 60738 533760 60794 533769
rect 60738 533695 60794 533704
rect 60738 533216 60794 533225
rect 60844 533202 60872 535622
rect 60794 533174 60872 533202
rect 60738 533151 60794 533160
rect 60740 521620 60792 521626
rect 60740 521562 60792 521568
rect 60752 517546 60780 521562
rect 60832 521552 60884 521558
rect 60832 521494 60884 521500
rect 60844 517614 60872 521494
rect 60924 518152 60976 518158
rect 60924 518094 60976 518100
rect 60936 517682 60964 518094
rect 61580 517993 61608 538727
rect 62212 527196 62264 527202
rect 62212 527138 62264 527144
rect 62120 522776 62172 522782
rect 62120 522718 62172 522724
rect 62132 522209 62160 522718
rect 62118 522200 62174 522209
rect 62118 522135 62174 522144
rect 62224 521626 62252 527138
rect 62500 523025 62528 560116
rect 63512 538214 63540 560116
rect 94594 560144 94650 560153
rect 63774 560079 63830 560088
rect 63788 558958 63816 560079
rect 64326 559736 64382 559745
rect 64326 559671 64382 559680
rect 63776 558952 63828 558958
rect 63776 558894 63828 558900
rect 63512 538186 63724 538214
rect 62856 525768 62908 525774
rect 62856 525710 62908 525716
rect 62486 523016 62542 523025
rect 62486 522951 62542 522960
rect 62212 521620 62264 521626
rect 62212 521562 62264 521568
rect 62868 521558 62896 525710
rect 63500 524340 63552 524346
rect 63500 524282 63552 524288
rect 63512 524249 63540 524282
rect 63498 524240 63554 524249
rect 63498 524175 63554 524184
rect 63500 522912 63552 522918
rect 63696 522889 63724 538186
rect 63500 522854 63552 522860
rect 63682 522880 63738 522889
rect 63512 522753 63540 522854
rect 63682 522815 63738 522824
rect 63498 522744 63554 522753
rect 63498 522679 63554 522688
rect 62856 521552 62908 521558
rect 62856 521494 62908 521500
rect 61936 521144 61988 521150
rect 61936 521086 61988 521092
rect 61948 518158 61976 521086
rect 62028 521076 62080 521082
rect 62028 521018 62080 521024
rect 62040 518226 62068 521018
rect 62028 518220 62080 518226
rect 62028 518162 62080 518168
rect 61936 518152 61988 518158
rect 64340 518106 64368 559671
rect 64524 523977 64552 560116
rect 64788 530596 64840 530602
rect 64788 530538 64840 530544
rect 64800 527202 64828 530538
rect 64788 527196 64840 527202
rect 64788 527138 64840 527144
rect 64510 523968 64566 523977
rect 64510 523903 64566 523912
rect 65536 523841 65564 560116
rect 65890 558240 65946 558249
rect 65890 558175 65946 558184
rect 65522 523832 65578 523841
rect 65522 523767 65578 523776
rect 65904 518106 65932 558175
rect 66548 536625 66576 560116
rect 67454 555384 67510 555393
rect 67454 555319 67510 555328
rect 66534 536616 66590 536625
rect 66534 536551 66590 536560
rect 66168 527196 66220 527202
rect 66168 527138 66220 527144
rect 66180 525978 66208 527138
rect 66168 525972 66220 525978
rect 66168 525914 66220 525920
rect 66168 524272 66220 524278
rect 66168 524214 66220 524220
rect 66180 524113 66208 524214
rect 66166 524104 66222 524113
rect 66166 524039 66222 524048
rect 67468 518106 67496 555319
rect 67560 531298 67588 560116
rect 68284 558952 68336 558958
rect 68284 558894 68336 558900
rect 67916 532840 67968 532846
rect 67916 532782 67968 532788
rect 67560 531270 67680 531298
rect 67548 531208 67600 531214
rect 67652 531185 67680 531270
rect 67548 531150 67600 531156
rect 67638 531176 67694 531185
rect 67560 530233 67588 531150
rect 67638 531111 67694 531120
rect 67928 530602 67956 532782
rect 67916 530596 67968 530602
rect 67916 530538 67968 530544
rect 67546 530224 67602 530233
rect 67546 530159 67602 530168
rect 68296 520946 68324 558894
rect 68572 532137 68600 560116
rect 68926 554024 68982 554033
rect 68926 553959 68982 553968
rect 68558 532128 68614 532137
rect 68558 532063 68614 532072
rect 68652 529780 68704 529786
rect 68652 529722 68704 529728
rect 68664 527202 68692 529722
rect 68652 527196 68704 527202
rect 68652 527138 68704 527144
rect 68284 520940 68336 520946
rect 68284 520882 68336 520888
rect 61936 518094 61988 518100
rect 64264 518078 64368 518106
rect 65828 518078 65932 518106
rect 67392 518078 67496 518106
rect 68940 518106 68968 553959
rect 69584 524113 69612 560116
rect 70610 560102 70716 560130
rect 70582 551576 70638 551585
rect 70582 551511 70638 551520
rect 70492 534132 70544 534138
rect 70492 534074 70544 534080
rect 70400 533996 70452 534002
rect 70400 533938 70452 533944
rect 70412 533089 70440 533938
rect 70398 533080 70454 533089
rect 70398 533015 70454 533024
rect 70504 532794 70532 534074
rect 70320 532766 70532 532794
rect 70320 529786 70348 532766
rect 70308 529780 70360 529786
rect 70308 529722 70360 529728
rect 69664 524204 69716 524210
rect 69664 524146 69716 524152
rect 69570 524104 69626 524113
rect 69570 524039 69626 524048
rect 69676 523569 69704 524146
rect 69662 523560 69718 523569
rect 69662 523495 69718 523504
rect 70596 518106 70624 551511
rect 70688 533633 70716 560102
rect 71044 549296 71096 549302
rect 71044 549238 71096 549244
rect 70674 533624 70730 533633
rect 70674 533559 70730 533568
rect 71056 532846 71084 549238
rect 71608 538665 71636 560116
rect 71778 551712 71834 551721
rect 71778 551647 71834 551656
rect 71792 551313 71820 551647
rect 71778 551304 71834 551313
rect 71778 551239 71834 551248
rect 71792 547874 71820 551239
rect 71792 547846 72188 547874
rect 71594 538656 71650 538665
rect 71594 538591 71650 538600
rect 71044 532840 71096 532846
rect 71044 532782 71096 532788
rect 72160 518106 72188 547846
rect 72424 543720 72476 543726
rect 72424 543662 72476 543668
rect 72436 534138 72464 543662
rect 72620 543561 72648 560116
rect 73160 554736 73212 554742
rect 73160 554678 73212 554684
rect 73172 553761 73200 554678
rect 73632 554441 73660 560116
rect 73618 554432 73674 554441
rect 73618 554367 73674 554376
rect 73158 553752 73214 553761
rect 73158 553687 73214 553696
rect 73710 551984 73766 551993
rect 73710 551919 73766 551928
rect 72606 543552 72662 543561
rect 72606 543487 72662 543496
rect 72424 534132 72476 534138
rect 72424 534074 72476 534080
rect 73724 518106 73752 551919
rect 74644 540297 74672 560116
rect 75274 552800 75330 552809
rect 75274 552735 75330 552744
rect 74630 540288 74686 540297
rect 74630 540223 74686 540232
rect 75288 518106 75316 552735
rect 75656 549273 75684 560116
rect 76012 559564 76064 559570
rect 76012 559506 76064 559512
rect 76024 557534 76052 559506
rect 75840 557506 76052 557534
rect 75840 549302 75868 557506
rect 75828 549296 75880 549302
rect 75642 549264 75698 549273
rect 75828 549238 75880 549244
rect 75642 549199 75698 549208
rect 75828 549160 75880 549166
rect 75828 549102 75880 549108
rect 75840 548185 75868 549102
rect 75826 548176 75882 548185
rect 75826 548111 75882 548120
rect 75828 545216 75880 545222
rect 75828 545158 75880 545164
rect 75840 543794 75868 545158
rect 75828 543788 75880 543794
rect 75828 543730 75880 543736
rect 76668 541657 76696 560116
rect 76838 555520 76894 555529
rect 76838 555455 76894 555464
rect 76654 541648 76710 541657
rect 76654 541583 76710 541592
rect 75828 540796 75880 540802
rect 75828 540738 75880 540744
rect 75840 540025 75868 540738
rect 75826 540016 75882 540025
rect 75826 539951 75882 539960
rect 76852 518106 76880 555455
rect 77680 547369 77708 560116
rect 78402 553072 78458 553081
rect 78402 553007 78458 553016
rect 77666 547360 77722 547369
rect 77666 547295 77722 547304
rect 78416 518106 78444 553007
rect 78588 547868 78640 547874
rect 78588 547810 78640 547816
rect 78600 546961 78628 547810
rect 78586 546952 78642 546961
rect 78586 546887 78642 546896
rect 78692 545737 78720 560116
rect 79324 546304 79376 546310
rect 79324 546246 79376 546252
rect 78678 545728 78734 545737
rect 78678 545663 78734 545672
rect 79336 545601 79364 546246
rect 79322 545592 79378 545601
rect 79322 545527 79378 545536
rect 79704 544921 79732 560116
rect 79966 554160 80022 554169
rect 79966 554095 80022 554104
rect 79690 544912 79746 544921
rect 79690 544847 79746 544856
rect 79980 518106 80008 554095
rect 80716 522753 80744 560116
rect 81530 558376 81586 558385
rect 81530 558311 81586 558320
rect 81440 553376 81492 553382
rect 81440 553318 81492 553324
rect 81452 552401 81480 553318
rect 81438 552392 81494 552401
rect 81438 552327 81494 552336
rect 81440 551812 81492 551818
rect 81440 551754 81492 551760
rect 81452 550905 81480 551754
rect 81438 550896 81494 550905
rect 81438 550831 81494 550840
rect 80702 522744 80758 522753
rect 80060 522708 80112 522714
rect 80702 522679 80758 522688
rect 80060 522650 80112 522656
rect 80072 521937 80100 522650
rect 80058 521928 80114 521937
rect 80058 521863 80114 521872
rect 81544 518106 81572 558311
rect 81728 553217 81756 560116
rect 81714 553208 81770 553217
rect 81714 553143 81770 553152
rect 82740 551177 82768 560116
rect 83094 555656 83150 555665
rect 83094 555591 83150 555600
rect 82726 551168 82782 551177
rect 82726 551103 82782 551112
rect 81808 549296 81860 549302
rect 81808 549238 81860 549244
rect 81820 545222 81848 549238
rect 81808 545216 81860 545222
rect 81808 545158 81860 545164
rect 82820 538144 82872 538150
rect 82820 538086 82872 538092
rect 82832 537441 82860 538086
rect 82818 537432 82874 537441
rect 82818 537367 82874 537376
rect 83108 518106 83136 555591
rect 83752 537441 83780 560116
rect 84658 555792 84714 555801
rect 84658 555727 84714 555736
rect 83738 537432 83794 537441
rect 83738 537367 83794 537376
rect 84672 518106 84700 555727
rect 84764 550089 84792 560116
rect 85488 550588 85540 550594
rect 85488 550530 85540 550536
rect 84750 550080 84806 550089
rect 84750 550015 84806 550024
rect 85500 549953 85528 550530
rect 85486 549944 85542 549953
rect 85486 549879 85542 549888
rect 85776 548593 85804 560116
rect 86222 556744 86278 556753
rect 86222 556679 86278 556688
rect 85762 548584 85818 548593
rect 85762 548519 85818 548528
rect 86236 518106 86264 556679
rect 86788 539345 86816 560116
rect 87814 560102 87920 560130
rect 87786 559600 87842 559609
rect 87786 559535 87842 559544
rect 86960 556232 87012 556238
rect 86960 556174 87012 556180
rect 86972 550746 87000 556174
rect 86880 550718 87000 550746
rect 86880 549506 86908 550718
rect 86868 549500 86920 549506
rect 86868 549442 86920 549448
rect 86868 549228 86920 549234
rect 86868 549170 86920 549176
rect 86880 548321 86908 549170
rect 86866 548312 86922 548321
rect 86866 548247 86922 548256
rect 86868 539572 86920 539578
rect 86868 539514 86920 539520
rect 86774 539336 86830 539345
rect 86774 539271 86830 539280
rect 86880 538529 86908 539514
rect 86866 538520 86922 538529
rect 86866 538455 86922 538464
rect 86868 523048 86920 523054
rect 86868 522990 86920 522996
rect 86880 521150 86908 522990
rect 86868 521144 86920 521150
rect 86868 521086 86920 521092
rect 87800 518106 87828 559535
rect 87892 543017 87920 560102
rect 88812 554169 88840 560116
rect 89350 556880 89406 556889
rect 89350 556815 89406 556824
rect 88984 554668 89036 554674
rect 88984 554610 89036 554616
rect 88798 554160 88854 554169
rect 88798 554095 88854 554104
rect 88996 553625 89024 554610
rect 88982 553616 89038 553625
rect 88982 553551 89038 553560
rect 87878 543008 87934 543017
rect 87878 542943 87934 542952
rect 89364 518106 89392 556815
rect 89720 547800 89772 547806
rect 89720 547742 89772 547748
rect 89732 546825 89760 547742
rect 89824 547097 89852 560116
rect 89810 547088 89866 547097
rect 89810 547023 89866 547032
rect 89718 546816 89774 546825
rect 89718 546751 89774 546760
rect 89720 546168 89772 546174
rect 89720 546110 89772 546116
rect 89732 545465 89760 546110
rect 90836 545873 90864 560116
rect 90916 559632 90968 559638
rect 90916 559574 90968 559580
rect 90928 556238 90956 559574
rect 91006 558512 91062 558521
rect 91006 558447 91062 558456
rect 91020 557705 91048 558447
rect 91006 557696 91062 557705
rect 91006 557631 91062 557640
rect 90916 556232 90968 556238
rect 90916 556174 90968 556180
rect 91020 547874 91048 557631
rect 90928 547846 91048 547874
rect 90822 545864 90878 545873
rect 90822 545799 90878 545808
rect 89718 545456 89774 545465
rect 89718 545391 89774 545400
rect 90928 518106 90956 547846
rect 91848 540977 91876 560116
rect 92388 556844 92440 556850
rect 92388 556786 92440 556792
rect 91834 540968 91890 540977
rect 91100 540932 91152 540938
rect 91834 540903 91890 540912
rect 91100 540874 91152 540880
rect 91112 539889 91140 540874
rect 91098 539880 91154 539889
rect 91098 539815 91154 539824
rect 68940 518078 68984 518106
rect 61566 517984 61622 517993
rect 64264 517956 64292 518078
rect 65828 517956 65856 518078
rect 67392 517956 67420 518078
rect 68956 517956 68984 518078
rect 70520 518078 70624 518106
rect 72084 518078 72188 518106
rect 73648 518078 73752 518106
rect 75212 518078 75316 518106
rect 76776 518078 76880 518106
rect 78340 518078 78444 518106
rect 79904 518078 80008 518106
rect 81468 518078 81572 518106
rect 83032 518078 83136 518106
rect 84596 518078 84700 518106
rect 86160 518078 86264 518106
rect 87724 518078 87828 518106
rect 89288 518078 89392 518106
rect 90852 518078 90956 518106
rect 92400 518106 92428 556786
rect 92480 545080 92532 545086
rect 92480 545022 92532 545028
rect 92492 544241 92520 545022
rect 92860 544513 92888 560116
rect 93886 560102 94176 560130
rect 94148 556617 94176 560102
rect 94594 560079 94650 560088
rect 94608 559473 94636 560079
rect 94226 559464 94282 559473
rect 94226 559399 94282 559408
rect 94594 559464 94650 559473
rect 94594 559399 94650 559408
rect 94134 556608 94190 556617
rect 94134 556543 94190 556552
rect 94240 547874 94268 559399
rect 94056 547846 94268 547874
rect 92846 544504 92902 544513
rect 92846 544439 92902 544448
rect 92478 544232 92534 544241
rect 92478 544167 92534 544176
rect 92480 527944 92532 527950
rect 92480 527886 92532 527892
rect 92492 523054 92520 527886
rect 92480 523048 92532 523054
rect 92480 522990 92532 522996
rect 94056 518106 94084 547846
rect 94884 543153 94912 560116
rect 95606 559056 95662 559065
rect 95606 558991 95662 559000
rect 95148 557320 95200 557326
rect 95148 557262 95200 557268
rect 95160 556481 95188 557262
rect 95146 556472 95202 556481
rect 95146 556407 95202 556416
rect 95148 543720 95200 543726
rect 95148 543662 95200 543668
rect 94870 543144 94926 543153
rect 94870 543079 94926 543088
rect 95160 542745 95188 543662
rect 95146 542736 95202 542745
rect 95146 542671 95202 542680
rect 95620 518106 95648 558991
rect 95896 532001 95924 560116
rect 96540 559065 96568 560215
rect 96526 559056 96582 559065
rect 96526 558991 96582 559000
rect 96908 535401 96936 560116
rect 97722 559464 97778 559473
rect 97722 559399 97778 559408
rect 97736 557534 97764 559399
rect 97814 559328 97870 559337
rect 97814 559263 97870 559272
rect 97828 558958 97856 559263
rect 97816 558952 97868 558958
rect 97816 558894 97868 558900
rect 97184 557506 97764 557534
rect 97184 557433 97212 557506
rect 97170 557424 97226 557433
rect 97170 557359 97226 557368
rect 96894 535392 96950 535401
rect 96894 535327 96950 535336
rect 96528 532704 96580 532710
rect 96528 532646 96580 532652
rect 96540 532273 96568 532646
rect 96526 532264 96582 532273
rect 96526 532199 96582 532208
rect 95882 531992 95938 532001
rect 95882 531927 95938 531936
rect 97184 518106 97212 557359
rect 97920 538214 97948 560116
rect 98748 558754 98776 560594
rect 98736 558748 98788 558754
rect 98736 558690 98788 558696
rect 98644 553240 98696 553246
rect 98644 553182 98696 553188
rect 98656 552265 98684 553182
rect 98642 552256 98698 552265
rect 98642 552191 98698 552200
rect 97828 538186 97948 538214
rect 97828 536217 97856 538186
rect 97908 536784 97960 536790
rect 97908 536726 97960 536732
rect 97814 536208 97870 536217
rect 97814 536143 97870 536152
rect 97920 535945 97948 536726
rect 97906 535936 97962 535945
rect 97906 535871 97962 535880
rect 97908 535424 97960 535430
rect 97908 535366 97960 535372
rect 97920 534313 97948 535366
rect 97906 534304 97962 534313
rect 97906 534239 97962 534248
rect 98748 518106 98776 558690
rect 98932 552945 98960 560116
rect 98918 552936 98974 552945
rect 98918 552871 98974 552880
rect 99380 551880 99432 551886
rect 99380 551822 99432 551828
rect 99392 550769 99420 551822
rect 99944 551313 99972 560116
rect 100850 557016 100906 557025
rect 100850 556951 100906 556960
rect 100760 556164 100812 556170
rect 100760 556106 100812 556112
rect 100772 554985 100800 556106
rect 100864 556073 100892 556951
rect 100850 556064 100906 556073
rect 100850 555999 100906 556008
rect 100758 554976 100814 554985
rect 100758 554911 100814 554920
rect 99930 551304 99986 551313
rect 99930 551239 99986 551248
rect 99378 550760 99434 550769
rect 99378 550695 99434 550704
rect 100760 550520 100812 550526
rect 100760 550462 100812 550468
rect 100772 549817 100800 550462
rect 100956 549953 100984 560116
rect 101862 556064 101918 556073
rect 101862 555999 101918 556008
rect 100942 549944 100998 549953
rect 100942 549879 100998 549888
rect 100758 549808 100814 549817
rect 100758 549743 100814 549752
rect 100760 525768 100812 525774
rect 100760 525710 100812 525716
rect 100772 525201 100800 525710
rect 100758 525192 100814 525201
rect 100758 525127 100814 525136
rect 99380 521620 99432 521626
rect 99380 521562 99432 521568
rect 99392 520849 99420 521562
rect 100298 521520 100354 521529
rect 100298 521455 100354 521464
rect 99378 520840 99434 520849
rect 99378 520775 99434 520784
rect 100312 518106 100340 521455
rect 101876 518106 101904 555999
rect 101968 525609 101996 560116
rect 102138 557288 102194 557297
rect 102138 557223 102194 557232
rect 102152 557025 102180 557223
rect 102138 557016 102194 557025
rect 102138 556951 102194 556960
rect 101954 525600 102010 525609
rect 101954 525535 102010 525544
rect 102140 525496 102192 525502
rect 102140 525438 102192 525444
rect 102152 525337 102180 525438
rect 102980 525337 103008 560116
rect 103426 557016 103482 557025
rect 103426 556951 103482 556960
rect 102138 525328 102194 525337
rect 102138 525263 102194 525272
rect 102966 525328 103022 525337
rect 102966 525263 103022 525272
rect 103440 518106 103468 556951
rect 103992 527105 104020 560116
rect 105018 560102 105124 560130
rect 104990 557288 105046 557297
rect 104990 557223 105046 557232
rect 103978 527096 104034 527105
rect 103978 527031 104034 527040
rect 105004 518106 105032 557223
rect 105096 526289 105124 560102
rect 106016 526969 106044 560116
rect 106554 553888 106610 553897
rect 106554 553823 106610 553832
rect 106002 526960 106058 526969
rect 106002 526895 106058 526904
rect 105082 526280 105138 526289
rect 105082 526215 105138 526224
rect 106568 518106 106596 553823
rect 107028 526833 107056 560116
rect 107568 554600 107620 554606
rect 107568 554542 107620 554548
rect 107580 553489 107608 554542
rect 107566 553480 107622 553489
rect 107566 553415 107622 553424
rect 107568 527060 107620 527066
rect 107568 527002 107620 527008
rect 107014 526824 107070 526833
rect 107014 526759 107070 526768
rect 107580 526425 107608 527002
rect 108040 526697 108068 560116
rect 108302 554568 108358 554577
rect 108302 554503 108358 554512
rect 108118 553752 108174 553761
rect 108118 553687 108174 553696
rect 108026 526688 108082 526697
rect 108026 526623 108082 526632
rect 107566 526416 107622 526425
rect 107566 526351 107622 526360
rect 108132 518106 108160 553687
rect 108316 553450 108344 554503
rect 108304 553444 108356 553450
rect 108304 553386 108356 553392
rect 109052 538214 109080 560116
rect 109132 558748 109184 558754
rect 109132 558690 109184 558696
rect 109144 557569 109172 558690
rect 109682 558512 109738 558521
rect 109682 558447 109738 558456
rect 109130 557560 109186 557569
rect 109130 557495 109186 557504
rect 109052 538186 109356 538214
rect 108304 527128 108356 527134
rect 108304 527070 108356 527076
rect 108316 526017 108344 527070
rect 109040 526992 109092 526998
rect 109040 526934 109092 526940
rect 109052 526153 109080 526934
rect 109132 526924 109184 526930
rect 109132 526866 109184 526872
rect 109038 526144 109094 526153
rect 109038 526079 109094 526088
rect 108302 526008 108358 526017
rect 108302 525943 108358 525952
rect 109144 525881 109172 526866
rect 109328 526561 109356 538186
rect 109314 526552 109370 526561
rect 109314 526487 109370 526496
rect 109130 525872 109186 525881
rect 109130 525807 109186 525816
rect 109696 518106 109724 558447
rect 110064 526425 110092 560116
rect 111076 526522 111104 560116
rect 111800 542360 111852 542366
rect 111800 542302 111852 542308
rect 111812 541385 111840 542302
rect 111798 541376 111854 541385
rect 111798 541311 111854 541320
rect 111800 531140 111852 531146
rect 111800 531082 111852 531088
rect 111812 530097 111840 531082
rect 112088 530913 112116 560116
rect 112810 557424 112866 557433
rect 112810 557359 112866 557368
rect 112074 530904 112130 530913
rect 112074 530839 112130 530848
rect 111798 530088 111854 530097
rect 111798 530023 111854 530032
rect 111064 526516 111116 526522
rect 111064 526458 111116 526464
rect 110050 526416 110106 526425
rect 110050 526351 110106 526360
rect 111246 521656 111302 521665
rect 111246 521591 111302 521600
rect 110420 521552 110472 521558
rect 110420 521494 110472 521500
rect 110432 520713 110460 521494
rect 110418 520704 110474 520713
rect 110418 520639 110474 520648
rect 111260 518106 111288 521591
rect 112824 518106 112852 557359
rect 113100 541793 113128 560116
rect 113086 541784 113142 541793
rect 113086 541719 113142 541728
rect 113180 530596 113232 530602
rect 113180 530538 113232 530544
rect 113192 527950 113220 530538
rect 113180 527944 113232 527950
rect 113180 527886 113232 527892
rect 114112 522209 114140 560116
rect 114468 522640 114520 522646
rect 114468 522582 114520 522588
rect 114098 522200 114154 522209
rect 114098 522135 114154 522144
rect 114480 521801 114508 522582
rect 114466 521792 114522 521801
rect 114466 521727 114522 521736
rect 114468 521484 114520 521490
rect 114468 521426 114520 521432
rect 114374 520840 114430 520849
rect 114374 520775 114430 520784
rect 114388 518106 114416 520775
rect 114480 520577 114508 521426
rect 115124 521393 115152 560116
rect 115846 554704 115902 554713
rect 115846 554639 115902 554648
rect 115754 554568 115810 554577
rect 115754 554503 115810 554512
rect 115768 547874 115796 554503
rect 115860 553518 115888 554639
rect 115848 553512 115900 553518
rect 115848 553454 115900 553460
rect 115768 547846 115888 547874
rect 115756 521416 115808 521422
rect 115110 521384 115166 521393
rect 115756 521358 115808 521364
rect 115110 521319 115166 521328
rect 114466 520568 114522 520577
rect 114466 520503 114522 520512
rect 115768 520305 115796 521358
rect 115754 520296 115810 520305
rect 115754 520231 115810 520240
rect 92400 518078 92444 518106
rect 70520 517956 70548 518078
rect 72084 517956 72112 518078
rect 73648 517956 73676 518078
rect 75212 517956 75240 518078
rect 76776 517956 76804 518078
rect 78340 517956 78368 518078
rect 79904 517956 79932 518078
rect 81468 517956 81496 518078
rect 83032 517956 83060 518078
rect 84596 517956 84624 518078
rect 86160 517956 86188 518078
rect 87724 517956 87752 518078
rect 89288 517956 89316 518078
rect 90852 517956 90880 518078
rect 92416 517956 92444 518078
rect 93980 518078 94084 518106
rect 95544 518078 95648 518106
rect 97108 518078 97212 518106
rect 98672 518078 98776 518106
rect 100236 518078 100340 518106
rect 101800 518078 101904 518106
rect 103364 518078 103468 518106
rect 104928 518078 105032 518106
rect 106492 518078 106596 518106
rect 108056 518078 108160 518106
rect 109620 518078 109724 518106
rect 111184 518078 111288 518106
rect 112748 518078 112852 518106
rect 114312 518078 114416 518106
rect 115860 518106 115888 547846
rect 116136 521257 116164 560116
rect 117148 532273 117176 560116
rect 117778 558784 117834 558793
rect 117778 558719 117834 558728
rect 117502 558104 117558 558113
rect 117502 558039 117558 558048
rect 117228 532636 117280 532642
rect 117228 532578 117280 532584
rect 117134 532264 117190 532273
rect 117134 532199 117190 532208
rect 117240 531729 117268 532578
rect 117226 531720 117282 531729
rect 117226 531655 117282 531664
rect 117228 521348 117280 521354
rect 117228 521290 117280 521296
rect 116122 521248 116178 521257
rect 116122 521183 116178 521192
rect 117240 520441 117268 521290
rect 117226 520432 117282 520441
rect 117226 520367 117282 520376
rect 117516 518106 117544 558039
rect 117792 557598 117820 558719
rect 117962 558648 118018 558657
rect 117962 558583 118018 558592
rect 117976 557734 118004 558583
rect 118160 557977 118188 560116
rect 119066 558920 119122 558929
rect 119066 558855 119122 558864
rect 118146 557968 118202 557977
rect 118146 557903 118202 557912
rect 117964 557728 118016 557734
rect 117964 557670 118016 557676
rect 117780 557592 117832 557598
rect 117780 557534 117832 557540
rect 118700 539504 118752 539510
rect 118700 539446 118752 539452
rect 118712 538393 118740 539446
rect 118698 538384 118754 538393
rect 118698 538319 118754 538328
rect 118700 525428 118752 525434
rect 118700 525370 118752 525376
rect 118712 524929 118740 525370
rect 118698 524920 118754 524929
rect 118698 524855 118754 524864
rect 119080 518106 119108 558855
rect 119172 525201 119200 560116
rect 120184 558793 120212 560116
rect 120170 558784 120226 558793
rect 120170 558719 120226 558728
rect 120080 558680 120132 558686
rect 120080 558622 120132 558628
rect 120170 558648 120226 558657
rect 119342 557968 119398 557977
rect 119342 557903 119398 557912
rect 119356 538937 119384 557903
rect 120092 557705 120120 558622
rect 120170 558583 120226 558592
rect 120814 558648 120870 558657
rect 120814 558583 120870 558592
rect 120078 557696 120134 557705
rect 120184 557666 120212 558583
rect 120078 557631 120134 557640
rect 120172 557660 120224 557666
rect 120172 557602 120224 557608
rect 120828 547874 120856 558583
rect 120644 547846 120856 547874
rect 119342 538928 119398 538937
rect 119342 538863 119398 538872
rect 120080 525700 120132 525706
rect 120080 525642 120132 525648
rect 119158 525192 119214 525201
rect 119158 525127 119214 525136
rect 120092 525065 120120 525642
rect 120078 525056 120134 525065
rect 120078 524991 120134 525000
rect 120644 518106 120672 547846
rect 121196 525065 121224 560116
rect 122222 560102 122328 560130
rect 122102 558784 122158 558793
rect 122102 558719 122158 558728
rect 121460 556096 121512 556102
rect 121460 556038 121512 556044
rect 121472 554849 121500 556038
rect 121458 554840 121514 554849
rect 121458 554775 121514 554784
rect 121460 546236 121512 546242
rect 121460 546178 121512 546184
rect 121472 545329 121500 546178
rect 121458 545320 121514 545329
rect 121458 545255 121514 545264
rect 121460 540864 121512 540870
rect 121460 540806 121512 540812
rect 121472 539753 121500 540806
rect 122116 540705 122144 558719
rect 122194 555248 122250 555257
rect 122194 555183 122250 555192
rect 122102 540696 122158 540705
rect 122102 540631 122158 540640
rect 121458 539744 121514 539753
rect 121458 539679 121514 539688
rect 121182 525056 121238 525065
rect 121182 524991 121238 525000
rect 122208 518106 122236 555183
rect 122300 545601 122328 560102
rect 122286 545592 122342 545601
rect 122286 545527 122342 545536
rect 123220 537849 123248 560116
rect 124232 558929 124260 560116
rect 124218 558920 124274 558929
rect 124218 558855 124274 558864
rect 123772 556022 124260 556050
rect 123206 537840 123262 537849
rect 123206 537775 123262 537784
rect 123772 518106 123800 556022
rect 124126 555928 124182 555937
rect 124232 555914 124260 556022
rect 124402 555928 124458 555937
rect 124232 555886 124402 555914
rect 124126 555863 124182 555872
rect 124402 555863 124458 555872
rect 124140 554810 124168 555863
rect 124128 554804 124180 554810
rect 124128 554746 124180 554752
rect 124864 551404 124916 551410
rect 124864 551346 124916 551352
rect 124128 538076 124180 538082
rect 124128 538018 124180 538024
rect 124140 537305 124168 538018
rect 124126 537296 124182 537305
rect 124126 537231 124182 537240
rect 124876 530602 124904 551346
rect 125244 543289 125272 560116
rect 126256 546961 126284 560116
rect 126334 558920 126390 558929
rect 126334 558855 126390 558864
rect 126348 548729 126376 558855
rect 126888 549092 126940 549098
rect 126888 549034 126940 549040
rect 126334 548720 126390 548729
rect 126334 548655 126390 548664
rect 126900 548049 126928 549034
rect 126886 548040 126942 548049
rect 126886 547975 126942 547984
rect 126888 547732 126940 547738
rect 126888 547674 126940 547680
rect 126242 546952 126298 546961
rect 126242 546887 126298 546896
rect 126900 546689 126928 547674
rect 126886 546680 126942 546689
rect 126886 546615 126942 546624
rect 125508 543652 125560 543658
rect 125508 543594 125560 543600
rect 125230 543280 125286 543289
rect 125230 543215 125286 543224
rect 125520 542609 125548 543594
rect 125506 542600 125562 542609
rect 125506 542535 125562 542544
rect 125322 537568 125378 537577
rect 125322 537503 125378 537512
rect 124864 530596 124916 530602
rect 124864 530538 124916 530544
rect 125336 518106 125364 537503
rect 127268 529689 127296 560116
rect 128280 547874 128308 560116
rect 128188 547846 128308 547874
rect 127624 545012 127676 545018
rect 127624 544954 127676 544960
rect 127636 544105 127664 544954
rect 128188 544649 128216 547846
rect 128174 544640 128230 544649
rect 128174 544575 128230 544584
rect 127622 544096 127678 544105
rect 127622 544031 127678 544040
rect 128360 536716 128412 536722
rect 128360 536658 128412 536664
rect 128372 535809 128400 536658
rect 129292 536353 129320 560116
rect 129278 536344 129334 536353
rect 129278 536279 129334 536288
rect 128358 535800 128414 535809
rect 128358 535735 128414 535744
rect 127624 529780 127676 529786
rect 127624 529722 127676 529728
rect 127254 529680 127310 529689
rect 127254 529615 127310 529624
rect 127636 528873 127664 529722
rect 127622 528864 127678 528873
rect 127622 528799 127678 528808
rect 130304 523977 130332 560116
rect 131120 539436 131172 539442
rect 131120 539378 131172 539384
rect 131132 538257 131160 539378
rect 131316 539073 131344 560116
rect 131302 539064 131358 539073
rect 131302 538999 131358 539008
rect 131118 538248 131174 538257
rect 131118 538183 131174 538192
rect 131120 532568 131172 532574
rect 131120 532510 131172 532516
rect 131132 531593 131160 532510
rect 132328 532409 132356 560116
rect 133142 536616 133198 536625
rect 133142 536551 133198 536560
rect 132314 532400 132370 532409
rect 132314 532335 132370 532344
rect 131118 531584 131174 531593
rect 131118 531519 131174 531528
rect 130014 523968 130070 523977
rect 130014 523903 130070 523912
rect 130290 523968 130346 523977
rect 130290 523903 130346 523912
rect 126886 523016 126942 523025
rect 126886 522951 126942 522960
rect 126900 518106 126928 522951
rect 128450 522880 128506 522889
rect 128450 522815 128506 522824
rect 128464 518106 128492 522815
rect 130028 518106 130056 523903
rect 131578 523832 131634 523841
rect 131578 523767 131634 523776
rect 131592 518106 131620 523767
rect 133156 518106 133184 536551
rect 133340 524929 133368 560116
rect 134536 529009 134564 634786
rect 134720 625154 134748 636278
rect 135258 636239 135314 636248
rect 134628 625126 134748 625154
rect 134628 549982 134656 625126
rect 134798 604480 134854 604489
rect 134798 604415 134854 604424
rect 134708 575544 134760 575550
rect 134708 575486 134760 575492
rect 134720 551410 134748 575486
rect 134708 551404 134760 551410
rect 134708 551346 134760 551352
rect 134616 549976 134668 549982
rect 134616 549918 134668 549924
rect 134706 531176 134762 531185
rect 134706 531111 134762 531120
rect 134522 529000 134578 529009
rect 134522 528935 134578 528944
rect 133788 525564 133840 525570
rect 133788 525506 133840 525512
rect 133326 524920 133382 524929
rect 133326 524855 133382 524864
rect 133800 524793 133828 525506
rect 133786 524784 133842 524793
rect 133786 524719 133842 524728
rect 134720 518106 134748 531111
rect 134812 521529 134840 604415
rect 135166 561640 135222 561649
rect 135166 561575 135222 561584
rect 135180 559570 135208 561575
rect 135168 559564 135220 559570
rect 135168 559506 135220 559512
rect 135272 558793 135300 636239
rect 135350 634944 135406 634953
rect 135350 634879 135406 634888
rect 135258 558784 135314 558793
rect 135258 558719 135314 558728
rect 135364 557433 135392 634879
rect 135350 557424 135406 557433
rect 135350 557359 135406 557368
rect 134982 556608 135038 556617
rect 134982 556543 135038 556552
rect 134996 521529 135024 556543
rect 135916 541890 135944 636754
rect 136008 547330 136036 636822
rect 136100 554062 136128 637327
rect 136914 635488 136970 635497
rect 136914 635423 136970 635432
rect 136638 635080 136694 635089
rect 136638 635015 136694 635024
rect 136088 554056 136140 554062
rect 136088 553998 136140 554004
rect 135996 547324 136048 547330
rect 135996 547266 136048 547272
rect 135904 541884 135956 541890
rect 135904 541826 135956 541832
rect 136270 532128 136326 532137
rect 136270 532063 136326 532072
rect 135168 529712 135220 529718
rect 135168 529654 135220 529660
rect 135180 528737 135208 529654
rect 135166 528728 135222 528737
rect 135166 528663 135222 528672
rect 134798 521520 134854 521529
rect 134798 521455 134854 521464
rect 134982 521520 135038 521529
rect 134982 521455 135038 521464
rect 136284 518106 136312 532063
rect 136652 520849 136680 635015
rect 136822 633992 136878 634001
rect 136822 633927 136878 633936
rect 136730 633856 136786 633865
rect 136730 633791 136786 633800
rect 136744 521665 136772 633791
rect 136836 558521 136864 633927
rect 136928 605169 136956 635423
rect 137282 619712 137338 619721
rect 137282 619647 137338 619656
rect 136914 605160 136970 605169
rect 136914 605095 136970 605104
rect 136928 604489 136956 605095
rect 136914 604480 136970 604489
rect 136914 604415 136970 604424
rect 136822 558512 136878 558521
rect 136822 558447 136878 558456
rect 137296 555558 137324 619647
rect 137466 598360 137522 598369
rect 137466 598295 137522 598304
rect 137374 576872 137430 576881
rect 137374 576807 137430 576816
rect 137284 555552 137336 555558
rect 137284 555494 137336 555500
rect 137388 523841 137416 576807
rect 137480 557025 137508 598295
rect 137650 597680 137706 597689
rect 137650 597615 137706 597624
rect 137560 585200 137612 585206
rect 137560 585142 137612 585148
rect 137572 575550 137600 585142
rect 137560 575544 137612 575550
rect 137560 575486 137612 575492
rect 137558 572928 137614 572937
rect 137558 572863 137614 572872
rect 137466 557016 137522 557025
rect 137466 556951 137522 556960
rect 137572 524385 137600 572863
rect 137664 560969 137692 597615
rect 137650 560960 137706 560969
rect 137650 560895 137706 560904
rect 137558 524376 137614 524385
rect 137558 524311 137614 524320
rect 137742 524104 137798 524113
rect 137742 524039 137798 524048
rect 137374 523832 137430 523841
rect 137374 523767 137430 523776
rect 136730 521656 136786 521665
rect 136730 521591 136786 521600
rect 136638 520840 136694 520849
rect 136638 520775 136694 520784
rect 115860 518078 115904 518106
rect 93980 517956 94008 518078
rect 95544 517956 95572 518078
rect 97108 517956 97136 518078
rect 98672 517956 98700 518078
rect 100236 517956 100264 518078
rect 101800 517956 101828 518078
rect 103364 517956 103392 518078
rect 104928 517956 104956 518078
rect 106492 517956 106520 518078
rect 108056 517956 108084 518078
rect 109620 517956 109648 518078
rect 111184 517956 111212 518078
rect 112748 517956 112776 518078
rect 114312 517956 114340 518078
rect 115876 517956 115904 518078
rect 117440 518078 117544 518106
rect 119004 518078 119108 518106
rect 120568 518078 120672 518106
rect 122132 518078 122236 518106
rect 123696 518078 123800 518106
rect 125260 518078 125364 518106
rect 126824 518078 126928 518106
rect 128388 518078 128492 518106
rect 129952 518078 130056 518106
rect 131516 518078 131620 518106
rect 133080 518078 133184 518106
rect 134644 518078 134748 518106
rect 136208 518078 136312 518106
rect 137756 518106 137784 524039
rect 137848 520266 137876 703520
rect 141422 699816 141478 699825
rect 141422 699751 141478 699760
rect 138020 658232 138072 658238
rect 138020 658174 138072 658180
rect 138032 657286 138060 658174
rect 141436 657558 141464 699751
rect 144184 683188 144236 683194
rect 144184 683130 144236 683136
rect 144196 657626 144224 683130
rect 153198 681864 153254 681873
rect 153198 681799 153254 681808
rect 153212 678994 153240 681799
rect 152476 678966 153240 678994
rect 152476 660929 152504 678966
rect 150530 660920 150586 660929
rect 150530 660855 150586 660864
rect 152462 660920 152518 660929
rect 152462 660855 152518 660864
rect 144184 657620 144236 657626
rect 144184 657562 144236 657568
rect 141424 657552 141476 657558
rect 141424 657494 141476 657500
rect 138020 657280 138072 657286
rect 138020 657222 138072 657228
rect 137836 520260 137888 520266
rect 137836 520202 137888 520208
rect 138032 519722 138060 657222
rect 148324 655580 148376 655586
rect 148324 655522 148376 655528
rect 140778 639568 140834 639577
rect 140778 639503 140834 639512
rect 138110 639024 138166 639033
rect 138110 638959 138166 638968
rect 139032 638988 139084 638994
rect 138124 558657 138152 638959
rect 139032 638930 139084 638936
rect 138664 636676 138716 636682
rect 138664 636618 138716 636624
rect 138110 558648 138166 558657
rect 138110 558583 138166 558592
rect 138676 539034 138704 636618
rect 138756 636608 138808 636614
rect 138756 636550 138808 636556
rect 138768 543114 138796 636550
rect 138846 635352 138902 635361
rect 138846 635287 138902 635296
rect 138860 602993 138888 635287
rect 138938 633448 138994 633457
rect 139044 633418 139072 638930
rect 139398 637800 139454 637809
rect 139398 637735 139454 637744
rect 138938 633383 138994 633392
rect 139032 633412 139084 633418
rect 138846 602984 138902 602993
rect 138846 602919 138902 602928
rect 138860 553761 138888 602919
rect 138952 600273 138980 633383
rect 139032 633354 139084 633360
rect 138938 600264 138994 600273
rect 138938 600199 138994 600208
rect 138952 557297 138980 600199
rect 139412 565842 139440 637735
rect 140042 636032 140098 636041
rect 140042 635967 140098 635976
rect 139490 634264 139546 634273
rect 139490 634199 139546 634208
rect 139504 566114 139532 634199
rect 140056 601633 140084 635967
rect 140042 601624 140098 601633
rect 140042 601559 140098 601568
rect 139504 566086 139716 566114
rect 139582 565856 139638 565865
rect 139412 565814 139532 565842
rect 139504 558113 139532 565814
rect 139582 565791 139638 565800
rect 139596 559638 139624 565791
rect 139584 559632 139636 559638
rect 139584 559574 139636 559580
rect 139490 558104 139546 558113
rect 139490 558039 139546 558048
rect 138938 557288 138994 557297
rect 138938 557223 138994 557232
rect 139688 555937 139716 566086
rect 139674 555928 139730 555937
rect 139674 555863 139730 555872
rect 140056 553897 140084 601559
rect 140792 554577 140820 639503
rect 140870 634672 140926 634681
rect 140870 634607 140926 634616
rect 140884 555257 140912 634607
rect 140962 634536 141018 634545
rect 140962 634471 141018 634480
rect 140976 559745 141004 634471
rect 144182 633448 144238 633457
rect 148336 633418 148364 655522
rect 150544 654134 150572 660855
rect 151084 654492 151136 654498
rect 151084 654434 151136 654440
rect 149808 654106 150572 654134
rect 149702 649904 149758 649913
rect 149702 649839 149758 649848
rect 144182 633383 144238 633392
rect 148324 633412 148376 633418
rect 142802 625152 142858 625161
rect 142802 625087 142858 625096
rect 141422 590608 141478 590617
rect 141422 590543 141478 590552
rect 141436 565865 141464 590543
rect 142158 569936 142214 569945
rect 142158 569871 142214 569880
rect 141422 565856 141478 565865
rect 141422 565791 141478 565800
rect 142172 561785 142200 569871
rect 142158 561776 142214 561785
rect 142158 561711 142214 561720
rect 140962 559736 141018 559745
rect 140962 559671 141018 559680
rect 140870 555248 140926 555257
rect 140870 555183 140926 555192
rect 140778 554568 140834 554577
rect 140778 554503 140834 554512
rect 142816 553897 142844 625087
rect 144196 590617 144224 633383
rect 148324 633354 148376 633360
rect 149716 629241 149744 649839
rect 149808 633457 149836 654106
rect 149794 633448 149850 633457
rect 149794 633383 149850 633392
rect 148414 629232 148470 629241
rect 148414 629167 148470 629176
rect 149702 629232 149758 629241
rect 149702 629167 149758 629176
rect 148322 623384 148378 623393
rect 148322 623319 148378 623328
rect 146942 621208 146998 621217
rect 146942 621143 146998 621152
rect 146298 603256 146354 603265
rect 146298 603191 146354 603200
rect 146312 598890 146340 603191
rect 145576 598862 146340 598890
rect 144276 590708 144328 590714
rect 144276 590650 144328 590656
rect 144182 590608 144238 590617
rect 144182 590543 144238 590552
rect 144182 585304 144238 585313
rect 144182 585239 144238 585248
rect 144196 569945 144224 585239
rect 144288 585206 144316 590650
rect 145576 585313 145604 598862
rect 145562 585304 145618 585313
rect 145562 585239 145618 585248
rect 144276 585200 144328 585206
rect 144276 585142 144328 585148
rect 144182 569936 144238 569945
rect 144182 569871 144238 569880
rect 146956 561105 146984 621143
rect 147404 594108 147456 594114
rect 147404 594050 147456 594056
rect 147416 590714 147444 594050
rect 147404 590708 147456 590714
rect 147404 590650 147456 590656
rect 146942 561096 146998 561105
rect 146942 561031 146998 561040
rect 144090 554432 144146 554441
rect 144090 554367 144146 554376
rect 140042 553888 140098 553897
rect 140042 553823 140098 553832
rect 142802 553888 142858 553897
rect 142802 553823 142858 553832
rect 138846 553752 138902 553761
rect 138846 553687 138902 553696
rect 142526 543552 142582 543561
rect 142526 543487 142582 543496
rect 138756 543108 138808 543114
rect 138756 543050 138808 543056
rect 138664 539028 138716 539034
rect 138664 538970 138716 538976
rect 140962 538656 141018 538665
rect 140962 538591 141018 538600
rect 139306 533624 139362 533633
rect 139306 533559 139362 533568
rect 138020 519716 138072 519722
rect 138020 519658 138072 519664
rect 139320 518106 139348 533559
rect 140976 518106 141004 538591
rect 142540 518106 142568 543487
rect 144104 518106 144132 554367
rect 147218 549264 147274 549273
rect 147218 549199 147274 549208
rect 145654 540288 145710 540297
rect 145654 540223 145710 540232
rect 145668 518106 145696 540223
rect 147232 518106 147260 549199
rect 148336 532137 148364 623319
rect 148428 603265 148456 629167
rect 148414 603256 148470 603265
rect 148414 603191 148470 603200
rect 151096 552702 151124 654434
rect 153566 652896 153622 652905
rect 153566 652831 153622 652840
rect 153580 649913 153608 652831
rect 153566 649904 153622 649913
rect 153566 649839 153622 649848
rect 152554 639840 152610 639849
rect 152554 639775 152610 639784
rect 152462 637256 152518 637265
rect 152462 637191 152518 637200
rect 151084 552696 151136 552702
rect 151084 552638 151136 552644
rect 150346 547360 150402 547369
rect 150346 547295 150402 547304
rect 148782 541648 148838 541657
rect 148782 541583 148838 541592
rect 148322 532128 148378 532137
rect 148322 532063 148378 532072
rect 148796 518106 148824 541583
rect 150360 518106 150388 547295
rect 151910 545728 151966 545737
rect 151910 545663 151966 545672
rect 151924 518106 151952 545663
rect 152476 538665 152504 637191
rect 152568 544241 152596 639775
rect 152646 622704 152702 622713
rect 152646 622639 152702 622648
rect 152660 561241 152688 622639
rect 152646 561232 152702 561241
rect 152646 561167 152702 561176
rect 153108 544944 153160 544950
rect 153108 544886 153160 544892
rect 153474 544912 153530 544921
rect 152554 544232 152610 544241
rect 152554 544167 152610 544176
rect 153120 543969 153148 544886
rect 153474 544847 153530 544856
rect 153106 543960 153162 543969
rect 153106 543895 153162 543904
rect 152462 538656 152518 538665
rect 152462 538591 152518 538600
rect 153488 518106 153516 544847
rect 154132 519654 154160 703520
rect 160098 700360 160154 700369
rect 160098 700295 160154 700304
rect 160112 698329 160140 700295
rect 156602 698320 156658 698329
rect 156602 698255 156658 698264
rect 160098 698320 160154 698329
rect 160098 698255 160154 698264
rect 156616 681873 156644 698255
rect 167642 687168 167698 687177
rect 167642 687103 167698 687112
rect 156602 681864 156658 681873
rect 156602 681799 156658 681808
rect 167656 679017 167684 687103
rect 167642 679008 167698 679017
rect 167642 678943 167698 678952
rect 158902 678192 158958 678201
rect 158902 678127 158958 678136
rect 158916 675889 158944 678127
rect 157982 675880 158038 675889
rect 157982 675815 158038 675824
rect 158902 675880 158958 675889
rect 158902 675815 158958 675824
rect 157996 666505 158024 675815
rect 155314 666496 155370 666505
rect 155314 666431 155370 666440
rect 157982 666496 158038 666505
rect 157982 666431 158038 666440
rect 155224 655648 155276 655654
rect 155224 655590 155276 655596
rect 155236 527882 155264 655590
rect 155328 652905 155356 666431
rect 170324 658238 170352 703520
rect 176934 700496 176990 700505
rect 176934 700431 176990 700440
rect 176948 698329 176976 700431
rect 202800 700369 202828 703520
rect 218992 700505 219020 703520
rect 218978 700496 219034 700505
rect 218978 700431 219034 700440
rect 202786 700360 202842 700369
rect 202786 700295 202842 700304
rect 173162 698320 173218 698329
rect 173162 698255 173218 698264
rect 176934 698320 176990 698329
rect 176934 698255 176990 698264
rect 173176 687313 173204 698255
rect 173162 687304 173218 687313
rect 173162 687239 173218 687248
rect 232504 668636 232556 668642
rect 232504 668578 232556 668584
rect 170312 658232 170364 658238
rect 170312 658174 170364 658180
rect 171140 658232 171192 658238
rect 171140 658174 171192 658180
rect 172428 658232 172480 658238
rect 172428 658174 172480 658180
rect 162124 657008 162176 657014
rect 162124 656950 162176 656956
rect 155314 652896 155370 652905
rect 155314 652831 155370 652840
rect 159364 648644 159416 648650
rect 159364 648586 159416 648592
rect 155314 639296 155370 639305
rect 155314 639231 155370 639240
rect 155328 528465 155356 639231
rect 155498 639160 155554 639169
rect 155498 639095 155554 639104
rect 155406 638616 155462 638625
rect 155406 638551 155462 638560
rect 155420 542881 155448 638551
rect 155406 542872 155462 542881
rect 155406 542807 155462 542816
rect 155512 534585 155540 639095
rect 157064 597508 157116 597514
rect 157064 597450 157116 597456
rect 157076 594114 157104 597450
rect 157064 594108 157116 594114
rect 157064 594050 157116 594056
rect 157982 581224 158038 581233
rect 157982 581159 158038 581168
rect 157996 554305 158024 581159
rect 158166 579728 158222 579737
rect 158166 579663 158222 579672
rect 158074 578368 158130 578377
rect 158074 578303 158130 578312
rect 157982 554296 158038 554305
rect 157982 554231 158038 554240
rect 156602 553208 156658 553217
rect 156602 553143 156658 553152
rect 155868 535356 155920 535362
rect 155868 535298 155920 535304
rect 155498 534576 155554 534585
rect 155498 534511 155554 534520
rect 155880 534177 155908 535298
rect 155866 534168 155922 534177
rect 155866 534103 155922 534112
rect 155314 528456 155370 528465
rect 155314 528391 155370 528400
rect 155224 527876 155276 527882
rect 155224 527818 155276 527824
rect 155038 522744 155094 522753
rect 155038 522679 155094 522688
rect 154120 519648 154172 519654
rect 154120 519590 154172 519596
rect 155052 518106 155080 522679
rect 156616 518106 156644 553143
rect 158088 552809 158116 578303
rect 158180 555529 158208 579663
rect 158350 576872 158406 576881
rect 158350 576807 158406 576816
rect 158166 555520 158222 555529
rect 158166 555455 158222 555464
rect 158074 552800 158130 552809
rect 158074 552735 158130 552744
rect 158364 551993 158392 576807
rect 158534 575512 158590 575521
rect 158534 575447 158590 575456
rect 158350 551984 158406 551993
rect 158350 551919 158406 551928
rect 158548 551721 158576 575447
rect 158534 551712 158590 551721
rect 158534 551647 158590 551656
rect 158166 551168 158222 551177
rect 158166 551103 158222 551112
rect 158180 518106 158208 551103
rect 159376 549030 159404 648586
rect 159454 636440 159510 636449
rect 159454 636375 159510 636384
rect 159364 549024 159416 549030
rect 159364 548966 159416 548972
rect 159468 545057 159496 636375
rect 159548 612060 159600 612066
rect 159548 612002 159600 612008
rect 159560 597514 159588 612002
rect 159548 597508 159600 597514
rect 159548 597450 159600 597456
rect 160834 594824 160890 594833
rect 160834 594759 160890 594768
rect 160742 593464 160798 593473
rect 160742 593399 160798 593408
rect 159546 581088 159602 581097
rect 159546 581023 159602 581032
rect 159560 553081 159588 581023
rect 160756 559473 160784 593399
rect 160848 560658 160876 594759
rect 160926 592104 160982 592113
rect 160926 592039 160982 592048
rect 160836 560652 160888 560658
rect 160836 560594 160888 560600
rect 160940 560289 160968 592039
rect 161110 590744 161166 590753
rect 161110 590679 161166 590688
rect 161018 575648 161074 575657
rect 161018 575583 161074 575592
rect 160926 560280 160982 560289
rect 160926 560215 160982 560224
rect 160742 559464 160798 559473
rect 160742 559399 160798 559408
rect 159546 553072 159602 553081
rect 159546 553007 159602 553016
rect 161032 551585 161060 575583
rect 161124 560153 161152 590679
rect 161202 570480 161258 570489
rect 161202 570415 161258 570424
rect 161110 560144 161166 560153
rect 161110 560079 161166 560088
rect 161018 551576 161074 551585
rect 161018 551511 161074 551520
rect 161216 546689 161244 570415
rect 161294 550080 161350 550089
rect 161294 550015 161350 550024
rect 161202 546680 161258 546689
rect 161202 546615 161258 546624
rect 159454 545048 159510 545057
rect 159454 544983 159510 544992
rect 159730 537432 159786 537441
rect 159730 537367 159786 537376
rect 159744 518106 159772 537367
rect 161308 518106 161336 550015
rect 162136 519586 162164 656950
rect 163594 636576 163650 636585
rect 162308 636540 162360 636546
rect 163594 636511 163650 636520
rect 162308 636482 162360 636488
rect 162214 624336 162270 624345
rect 162214 624271 162270 624280
rect 162228 533769 162256 624271
rect 162320 548690 162348 636482
rect 163502 625968 163558 625977
rect 163502 625903 163558 625912
rect 162308 548684 162360 548690
rect 162308 548626 162360 548632
rect 162766 548584 162822 548593
rect 162766 548519 162822 548528
rect 162214 533760 162270 533769
rect 162214 533695 162270 533704
rect 162124 519580 162176 519586
rect 162124 519522 162176 519528
rect 137756 518078 137800 518106
rect 139320 518078 139364 518106
rect 117440 517956 117468 518078
rect 119004 517956 119032 518078
rect 120568 517956 120596 518078
rect 122132 517956 122160 518078
rect 123696 517956 123724 518078
rect 125260 517956 125288 518078
rect 126824 517956 126852 518078
rect 128388 517956 128416 518078
rect 129952 517956 129980 518078
rect 131516 517956 131544 518078
rect 133080 517956 133108 518078
rect 134644 517956 134672 518078
rect 136208 517956 136236 518078
rect 137772 517956 137800 518078
rect 139336 517956 139364 518078
rect 140900 518078 141004 518106
rect 142464 518078 142568 518106
rect 144028 518078 144132 518106
rect 145592 518078 145696 518106
rect 147156 518078 147260 518106
rect 148720 518078 148824 518106
rect 150284 518078 150388 518106
rect 151848 518078 151952 518106
rect 153412 518078 153516 518106
rect 154976 518078 155080 518106
rect 156540 518078 156644 518106
rect 158104 518078 158208 518106
rect 159668 518078 159772 518106
rect 161232 518078 161336 518106
rect 162780 518106 162808 548519
rect 163516 534449 163544 625903
rect 163608 552401 163636 636511
rect 170404 635588 170456 635594
rect 170404 635530 170456 635536
rect 170416 622470 170444 635530
rect 164976 622464 165028 622470
rect 164976 622406 165028 622412
rect 170404 622464 170456 622470
rect 170404 622406 170456 622412
rect 164882 619440 164938 619449
rect 164882 619375 164938 619384
rect 163778 591016 163834 591025
rect 163778 590951 163834 590960
rect 163686 568848 163742 568857
rect 163686 568783 163742 568792
rect 163594 552392 163650 552401
rect 163594 552327 163650 552336
rect 163502 534440 163558 534449
rect 163502 534375 163558 534384
rect 163700 520010 163728 568783
rect 163792 556850 163820 590951
rect 163870 589384 163926 589393
rect 163870 589319 163926 589328
rect 163884 558686 163912 589319
rect 163962 588296 164018 588305
rect 163962 588231 164018 588240
rect 163872 558680 163924 558686
rect 163872 558622 163924 558628
rect 163976 556889 164004 588231
rect 164054 574560 164110 574569
rect 164054 574495 164110 574504
rect 163962 556880 164018 556889
rect 163780 556844 163832 556850
rect 163962 556815 164018 556824
rect 163780 556786 163832 556792
rect 164068 554033 164096 574495
rect 164054 554024 164110 554033
rect 164054 553959 164110 553968
rect 164422 539336 164478 539345
rect 164422 539271 164478 539280
rect 164146 535392 164202 535401
rect 164146 535327 164202 535336
rect 164160 534274 164188 535327
rect 164148 534268 164200 534274
rect 164148 534210 164200 534216
rect 163700 519982 164280 520010
rect 164148 519852 164200 519858
rect 164148 519794 164200 519800
rect 164160 519761 164188 519794
rect 164146 519752 164202 519761
rect 164252 519738 164280 519982
rect 164330 519752 164386 519761
rect 164252 519710 164330 519738
rect 164146 519687 164202 519696
rect 164330 519687 164386 519696
rect 164436 518106 164464 539271
rect 164896 527921 164924 619375
rect 164988 612066 165016 622406
rect 169022 618624 169078 618633
rect 169022 618559 169078 618568
rect 166354 616992 166410 617001
rect 166354 616927 166410 616936
rect 166262 612912 166318 612921
rect 166262 612847 166318 612856
rect 164976 612060 165028 612066
rect 164976 612002 165028 612008
rect 164974 601488 165030 601497
rect 164974 601423 165030 601432
rect 164988 537577 165016 601423
rect 165986 543008 166042 543017
rect 165986 542943 166042 542952
rect 164974 537568 165030 537577
rect 164974 537503 165030 537512
rect 164882 527912 164938 527921
rect 164882 527847 164938 527856
rect 166000 518106 166028 542943
rect 166276 538214 166304 612847
rect 166368 555529 166396 616927
rect 167642 616176 167698 616185
rect 167642 616111 167698 616120
rect 166446 596592 166502 596601
rect 166446 596527 166502 596536
rect 166354 555520 166410 555529
rect 166354 555455 166410 555464
rect 166460 541657 166488 596527
rect 166538 585440 166594 585449
rect 166538 585375 166594 585384
rect 166552 555801 166580 585375
rect 166998 582176 167054 582185
rect 166998 582111 167054 582120
rect 167012 581233 167040 582111
rect 166998 581224 167054 581233
rect 166998 581159 167054 581168
rect 166906 575376 166962 575385
rect 166906 575311 166962 575320
rect 166722 573472 166778 573481
rect 166722 573407 166778 573416
rect 166632 569832 166684 569838
rect 166632 569774 166684 569780
rect 166644 556753 166672 569774
rect 166630 556744 166686 556753
rect 166630 556679 166686 556688
rect 166538 555792 166594 555801
rect 166538 555727 166594 555736
rect 166736 555393 166764 573407
rect 166816 559972 166868 559978
rect 166816 559914 166868 559920
rect 166828 559609 166856 559914
rect 166814 559600 166870 559609
rect 166814 559535 166870 559544
rect 166920 556753 166948 575311
rect 166906 556744 166962 556753
rect 166906 556679 166962 556688
rect 166722 555384 166778 555393
rect 166722 555319 166778 555328
rect 167550 554160 167606 554169
rect 167550 554095 167606 554104
rect 166446 541648 166502 541657
rect 166446 541583 166502 541592
rect 166184 538186 166304 538214
rect 166184 528714 166212 538186
rect 167000 533860 167052 533866
rect 167000 533802 167052 533808
rect 167012 532953 167040 533802
rect 166998 532944 167054 532953
rect 166998 532879 167054 532888
rect 166264 529644 166316 529650
rect 166264 529586 166316 529592
rect 166276 529417 166304 529586
rect 166262 529408 166318 529417
rect 166262 529343 166318 529352
rect 166262 528728 166318 528737
rect 166184 528686 166262 528714
rect 166262 528663 166318 528672
rect 167564 518106 167592 554095
rect 167656 543017 167684 616111
rect 167734 603936 167790 603945
rect 167734 603871 167790 603880
rect 167642 543008 167698 543017
rect 167642 542943 167698 542952
rect 167748 540297 167776 603871
rect 167918 597408 167974 597417
rect 167918 597343 167974 597352
rect 167826 595776 167882 595785
rect 167826 595711 167882 595720
rect 167734 540288 167790 540297
rect 167734 540223 167790 540232
rect 167840 533633 167868 595711
rect 167932 548593 167960 597343
rect 168286 582176 168342 582185
rect 168286 582111 168342 582120
rect 168194 579728 168250 579737
rect 168194 579663 168250 579672
rect 168010 574424 168066 574433
rect 168010 574359 168066 574368
rect 168024 556889 168052 574359
rect 168010 556880 168066 556889
rect 168010 556815 168066 556824
rect 168208 553081 168236 579663
rect 168194 553072 168250 553081
rect 168194 553007 168250 553016
rect 168300 550633 168328 582111
rect 168286 550624 168342 550633
rect 168286 550559 168342 550568
rect 167918 548584 167974 548593
rect 167918 548519 167974 548528
rect 169036 540394 169064 618559
rect 169298 608832 169354 608841
rect 169298 608767 169354 608776
rect 169206 603120 169262 603129
rect 169206 603055 169262 603064
rect 169114 583808 169170 583817
rect 169114 583743 169170 583752
rect 169128 555665 169156 583743
rect 169114 555656 169170 555665
rect 169114 555591 169170 555600
rect 169114 547088 169170 547097
rect 169114 547023 169170 547032
rect 169024 540388 169076 540394
rect 169024 540330 169076 540336
rect 167826 533624 167882 533633
rect 167826 533559 167882 533568
rect 169128 518106 169156 547023
rect 169220 528057 169248 603055
rect 169312 545737 169340 608767
rect 170494 605568 170550 605577
rect 170494 605503 170550 605512
rect 170402 594960 170458 594969
rect 170402 594895 170458 594904
rect 169758 593056 169814 593065
rect 169758 592991 169814 593000
rect 169772 592113 169800 592991
rect 169758 592104 169814 592113
rect 169758 592039 169814 592048
rect 169390 582448 169446 582457
rect 169390 582383 169446 582392
rect 169404 560046 169432 582383
rect 169758 578912 169814 578921
rect 169758 578847 169814 578856
rect 170310 578912 170366 578921
rect 170310 578847 170366 578856
rect 169772 578377 169800 578847
rect 169758 578368 169814 578377
rect 169758 578303 169814 578312
rect 170218 575648 170274 575657
rect 170218 575583 170274 575592
rect 169482 572928 169538 572937
rect 169482 572863 169538 572872
rect 169392 560040 169444 560046
rect 169392 559982 169444 559988
rect 169404 558385 169432 559982
rect 169390 558376 169446 558385
rect 169390 558311 169446 558320
rect 169496 557025 169524 572863
rect 169482 557016 169538 557025
rect 169482 556951 169538 556960
rect 169758 553208 169814 553217
rect 169758 553143 169814 553152
rect 169772 552090 169800 553143
rect 169760 552084 169812 552090
rect 169760 552026 169812 552032
rect 170232 551993 170260 575583
rect 170218 551984 170274 551993
rect 170218 551919 170274 551928
rect 169760 550384 169812 550390
rect 169760 550326 169812 550332
rect 169772 549681 169800 550326
rect 169758 549672 169814 549681
rect 169758 549607 169814 549616
rect 170324 549273 170352 578847
rect 170310 549264 170366 549273
rect 170310 549199 170366 549208
rect 169298 545728 169354 545737
rect 169298 545663 169354 545672
rect 170416 528193 170444 594895
rect 170508 537305 170536 605503
rect 170586 599856 170642 599865
rect 170586 599791 170642 599800
rect 170600 550089 170628 599791
rect 170678 597408 170734 597417
rect 170678 597343 170734 597352
rect 170692 556073 170720 597343
rect 170954 593328 171010 593337
rect 170954 593263 171010 593272
rect 170862 589248 170918 589257
rect 170862 589183 170918 589192
rect 170770 569664 170826 569673
rect 170770 569599 170826 569608
rect 170678 556064 170734 556073
rect 170678 555999 170734 556008
rect 170586 550080 170642 550089
rect 170586 550015 170642 550024
rect 170678 545864 170734 545873
rect 170678 545799 170734 545808
rect 170494 537296 170550 537305
rect 170494 537231 170550 537240
rect 170402 528184 170458 528193
rect 170402 528119 170458 528128
rect 169206 528048 169262 528057
rect 169206 527983 169262 527992
rect 169758 527912 169814 527921
rect 169758 527847 169814 527856
rect 169772 527202 169800 527847
rect 169760 527196 169812 527202
rect 169760 527138 169812 527144
rect 169760 524136 169812 524142
rect 169760 524078 169812 524084
rect 169772 523433 169800 524078
rect 169758 523424 169814 523433
rect 169758 523359 169814 523368
rect 170692 518106 170720 545799
rect 170784 524249 170812 569599
rect 170876 546281 170904 589183
rect 170968 556617 170996 593263
rect 171046 593056 171102 593065
rect 171046 592991 171102 593000
rect 171060 558793 171088 592991
rect 171046 558784 171102 558793
rect 171046 558719 171102 558728
rect 170954 556608 171010 556617
rect 170954 556543 171010 556552
rect 170862 546272 170918 546281
rect 170862 546207 170918 546216
rect 171046 537432 171102 537441
rect 171046 537367 171102 537376
rect 171060 536858 171088 537367
rect 171048 536852 171100 536858
rect 171048 536794 171100 536800
rect 170770 524240 170826 524249
rect 170770 524175 170826 524184
rect 171152 518294 171180 658174
rect 172440 657082 172468 658174
rect 172428 657076 172480 657082
rect 172428 657018 172480 657024
rect 204902 648408 204958 648417
rect 204902 648343 204958 648352
rect 193034 648272 193090 648281
rect 193034 648207 193090 648216
rect 186596 645992 186648 645998
rect 186596 645934 186648 645940
rect 176658 643648 176714 643657
rect 176658 643583 176660 643592
rect 176712 643583 176714 643592
rect 177670 643648 177726 643657
rect 177670 643583 177726 643592
rect 176660 643554 176712 643560
rect 177578 637120 177634 637129
rect 177578 637055 177634 637064
rect 176566 636848 176622 636857
rect 176566 636783 176622 636792
rect 174542 621888 174598 621897
rect 174542 621823 174598 621832
rect 173254 617808 173310 617817
rect 173254 617743 173310 617752
rect 171782 614544 171838 614553
rect 171782 614479 171838 614488
rect 171796 543734 171824 614479
rect 173162 607200 173218 607209
rect 173162 607135 173218 607144
rect 171874 606384 171930 606393
rect 171874 606319 171930 606328
rect 171704 543706 171824 543734
rect 171888 543734 171916 606319
rect 171966 600672 172022 600681
rect 171966 600607 172022 600616
rect 171980 544921 172008 600607
rect 172334 595232 172390 595241
rect 172334 595167 172390 595176
rect 172058 591696 172114 591705
rect 172058 591631 172114 591640
rect 171966 544912 172022 544921
rect 171966 544847 172022 544856
rect 171888 543706 172008 543734
rect 171704 536738 171732 543706
rect 171980 538286 172008 543706
rect 171968 538280 172020 538286
rect 171968 538222 172020 538228
rect 171784 538008 171836 538014
rect 171784 537950 171836 537956
rect 171796 537169 171824 537950
rect 172072 537713 172100 591631
rect 172242 586392 172298 586401
rect 172242 586327 172298 586336
rect 172150 572112 172206 572121
rect 172150 572047 172206 572056
rect 172164 557297 172192 572047
rect 172256 569838 172284 586327
rect 172244 569832 172296 569838
rect 172244 569774 172296 569780
rect 172150 557288 172206 557297
rect 172150 557223 172206 557232
rect 172256 554577 172284 569774
rect 172348 561649 172376 595167
rect 172426 586800 172482 586809
rect 172426 586735 172482 586744
rect 172334 561640 172390 561649
rect 172334 561575 172390 561584
rect 172242 554568 172298 554577
rect 172242 554503 172298 554512
rect 172440 547874 172468 586735
rect 172518 577824 172574 577833
rect 172518 577759 172574 577768
rect 172532 576881 172560 577759
rect 172518 576872 172574 576881
rect 172574 576826 173020 576854
rect 172518 576807 172574 576816
rect 172992 554441 173020 576826
rect 173072 560040 173124 560046
rect 173072 559982 173124 559988
rect 173084 557433 173112 559982
rect 173070 557424 173126 557433
rect 173070 557359 173126 557368
rect 172978 554432 173034 554441
rect 172978 554367 173034 554376
rect 172348 547846 172468 547874
rect 172348 540977 172376 547846
rect 172428 544876 172480 544882
rect 172428 544818 172480 544824
rect 172440 543833 172468 544818
rect 172426 543824 172482 543833
rect 172426 543759 172482 543768
rect 172518 543008 172574 543017
rect 172518 542943 172574 542952
rect 172532 542434 172560 542943
rect 172520 542428 172572 542434
rect 172520 542370 172572 542376
rect 172520 542224 172572 542230
rect 172520 542166 172572 542172
rect 172532 541249 172560 542166
rect 172518 541240 172574 541249
rect 172518 541175 172574 541184
rect 172150 540968 172206 540977
rect 172334 540968 172390 540977
rect 172206 540926 172284 540954
rect 172150 540903 172206 540912
rect 172058 537704 172114 537713
rect 172058 537639 172114 537648
rect 171782 537160 171838 537169
rect 171782 537095 171838 537104
rect 171782 536752 171838 536761
rect 171704 536710 171782 536738
rect 171782 536687 171838 536696
rect 171140 518288 171192 518294
rect 171140 518230 171192 518236
rect 172256 518106 172284 540926
rect 172334 540903 172390 540912
rect 173176 531185 173204 607135
rect 173268 551177 173296 617743
rect 174358 593464 174414 593473
rect 174358 593399 174414 593408
rect 173806 591968 173862 591977
rect 173806 591903 173862 591912
rect 173820 590753 173848 591903
rect 173806 590744 173862 590753
rect 173728 590702 173806 590730
rect 173438 590064 173494 590073
rect 173438 589999 173494 590008
rect 173346 588432 173402 588441
rect 173346 588367 173402 588376
rect 173254 551168 173310 551177
rect 173254 551103 173310 551112
rect 173360 542201 173388 588367
rect 173452 547369 173480 589999
rect 173530 581904 173586 581913
rect 173530 581839 173586 581848
rect 173438 547360 173494 547369
rect 173438 547295 173494 547304
rect 173544 543561 173572 581839
rect 173622 576192 173678 576201
rect 173622 576127 173678 576136
rect 173530 543552 173586 543561
rect 173530 543487 173586 543496
rect 173346 542192 173402 542201
rect 173346 542127 173402 542136
rect 173636 539345 173664 576127
rect 173728 560153 173756 590702
rect 173806 590679 173862 590688
rect 173806 587616 173862 587625
rect 173806 587551 173862 587560
rect 173714 560144 173770 560153
rect 173714 560079 173770 560088
rect 173820 559978 173848 587551
rect 173808 559972 173860 559978
rect 173808 559914 173860 559920
rect 173820 556073 173848 559914
rect 174372 559473 174400 593399
rect 174450 583808 174506 583817
rect 174450 583743 174506 583752
rect 174358 559464 174414 559473
rect 174358 559399 174414 559408
rect 174464 557705 174492 583743
rect 174450 557696 174506 557705
rect 174450 557631 174506 557640
rect 173806 556064 173862 556073
rect 173806 555999 173862 556008
rect 173806 552800 173862 552809
rect 173806 552735 173862 552744
rect 173820 552430 173848 552735
rect 173808 552424 173860 552430
rect 173808 552366 173860 552372
rect 173806 547768 173862 547777
rect 173806 547703 173862 547712
rect 173820 546514 173848 547703
rect 173808 546508 173860 546514
rect 173808 546450 173860 546456
rect 173714 544504 173770 544513
rect 173714 544439 173770 544448
rect 173728 543734 173756 544439
rect 173728 543706 173848 543734
rect 173622 539336 173678 539345
rect 173622 539271 173678 539280
rect 173162 531176 173218 531185
rect 173162 531111 173218 531120
rect 172426 526144 172482 526153
rect 172426 526079 172482 526088
rect 172440 525842 172468 526079
rect 172428 525836 172480 525842
rect 172428 525778 172480 525784
rect 173820 518106 173848 543706
rect 174556 540974 174584 621823
rect 174634 610464 174690 610473
rect 174634 610399 174690 610408
rect 174372 540946 174584 540974
rect 173990 536752 174046 536761
rect 173990 536687 174046 536696
rect 174004 535566 174032 536687
rect 173992 535560 174044 535566
rect 173992 535502 174044 535508
rect 174372 531314 174400 540946
rect 174648 532030 174676 610399
rect 174818 609648 174874 609657
rect 174818 609583 174874 609592
rect 174726 587480 174782 587489
rect 174726 587415 174782 587424
rect 174636 532024 174688 532030
rect 174636 531966 174688 531972
rect 174372 531286 174584 531314
rect 174556 523025 174584 531286
rect 174740 528329 174768 587415
rect 174832 555665 174860 609583
rect 176580 602993 176608 636783
rect 177592 626793 177620 637055
rect 177578 626784 177634 626793
rect 177578 626719 177634 626728
rect 177684 625705 177712 643583
rect 179326 643240 179382 643249
rect 179326 643175 179382 643184
rect 179340 643142 179368 643175
rect 179328 643136 179380 643142
rect 179328 643078 179380 643084
rect 179328 642048 179380 642054
rect 179328 641990 179380 641996
rect 177948 641980 178000 641986
rect 177948 641922 178000 641928
rect 177764 641912 177816 641918
rect 177764 641854 177816 641860
rect 177776 633321 177804 641854
rect 177856 641844 177908 641850
rect 177856 641786 177908 641792
rect 177762 633312 177818 633321
rect 177762 633247 177818 633256
rect 177868 631145 177896 641786
rect 177960 641753 177988 641922
rect 179340 641753 179368 641990
rect 177946 641744 178002 641753
rect 177946 641679 178002 641688
rect 179326 641744 179382 641753
rect 179326 641679 179382 641688
rect 185676 640484 185728 640490
rect 185676 640426 185728 640432
rect 184294 639160 184350 639169
rect 184294 639095 184350 639104
rect 183190 637800 183246 637809
rect 183112 637758 183190 637786
rect 179050 635624 179106 635633
rect 179050 635559 179106 635568
rect 177946 634672 178002 634681
rect 177946 634607 178002 634616
rect 177854 631136 177910 631145
rect 177854 631071 177910 631080
rect 177960 627881 177988 634607
rect 178958 633584 179014 633593
rect 178958 633519 179014 633528
rect 177946 627872 178002 627881
rect 177946 627807 178002 627816
rect 177670 625696 177726 625705
rect 177670 625631 177726 625640
rect 177302 612776 177358 612785
rect 177302 612711 177358 612720
rect 177210 610736 177266 610745
rect 177210 610671 177266 610680
rect 176566 602984 176622 602993
rect 176566 602919 176622 602928
rect 176198 602304 176254 602313
rect 176198 602239 176254 602248
rect 175922 599040 175978 599049
rect 175922 598975 175978 598984
rect 175094 594008 175150 594017
rect 175094 593943 175150 593952
rect 174910 590880 174966 590889
rect 174910 590815 174966 590824
rect 174818 555656 174874 555665
rect 174818 555591 174874 555600
rect 174924 544513 174952 590815
rect 175002 581360 175058 581369
rect 175002 581295 175058 581304
rect 174910 544504 174966 544513
rect 174910 544439 174966 544448
rect 175016 536625 175044 581295
rect 175108 556850 175136 593943
rect 175830 585440 175886 585449
rect 175830 585375 175886 585384
rect 175738 576736 175794 576745
rect 175738 576671 175794 576680
rect 175752 575521 175780 576671
rect 175738 575512 175794 575521
rect 175738 575447 175794 575456
rect 175462 571296 175518 571305
rect 175462 571231 175518 571240
rect 175476 567194 175504 571231
rect 175476 567166 175780 567194
rect 175370 561096 175426 561105
rect 175370 561031 175426 561040
rect 175186 560280 175242 560289
rect 175186 560215 175242 560224
rect 175096 556844 175148 556850
rect 175096 556786 175148 556792
rect 175002 536616 175058 536625
rect 175002 536551 175058 536560
rect 175200 534750 175228 560215
rect 175278 544912 175334 544921
rect 175278 544847 175334 544856
rect 175292 543794 175320 544847
rect 175280 543788 175332 543794
rect 175280 543730 175332 543736
rect 175280 543584 175332 543590
rect 175280 543526 175332 543532
rect 175292 542473 175320 543526
rect 175278 542464 175334 542473
rect 175278 542399 175334 542408
rect 175188 534744 175240 534750
rect 175188 534686 175240 534692
rect 175188 528488 175240 528494
rect 175188 528430 175240 528436
rect 174726 528320 174782 528329
rect 174726 528255 174782 528264
rect 175200 527649 175228 528430
rect 175186 527640 175242 527649
rect 175186 527575 175242 527584
rect 175186 525736 175242 525745
rect 175186 525671 175242 525680
rect 175200 524482 175228 525671
rect 175188 524476 175240 524482
rect 175188 524418 175240 524424
rect 174542 523016 174598 523025
rect 174542 522951 174598 522960
rect 175384 518106 175412 561031
rect 175752 544921 175780 567166
rect 175844 559201 175872 585375
rect 175830 559192 175886 559201
rect 175830 559127 175886 559136
rect 175830 553208 175886 553217
rect 175830 553143 175886 553152
rect 175844 552158 175872 553143
rect 175832 552152 175884 552158
rect 175832 552094 175884 552100
rect 175738 544912 175794 544921
rect 175738 544847 175794 544856
rect 175832 533792 175884 533798
rect 175832 533734 175884 533740
rect 175844 532817 175872 533734
rect 175830 532808 175886 532817
rect 175830 532743 175886 532752
rect 175832 528556 175884 528562
rect 175832 528498 175884 528504
rect 175844 527513 175872 528498
rect 175830 527504 175886 527513
rect 175830 527439 175886 527448
rect 175936 526454 175964 598975
rect 176014 584216 176070 584225
rect 176014 584151 176070 584160
rect 175924 526448 175976 526454
rect 175924 526390 175976 526396
rect 175924 525632 175976 525638
rect 175924 525574 175976 525580
rect 175936 524657 175964 525574
rect 175922 524648 175978 524657
rect 175922 524583 175978 524592
rect 176028 522753 176056 584151
rect 176106 582720 176162 582729
rect 176106 582655 176162 582664
rect 176120 525473 176148 582655
rect 176212 553217 176240 602239
rect 176580 601905 176608 602919
rect 176566 601896 176622 601905
rect 176566 601831 176622 601840
rect 176566 589792 176622 589801
rect 176566 589727 176622 589736
rect 176580 589393 176608 589727
rect 176566 589384 176622 589393
rect 176566 589319 176622 589328
rect 176474 585984 176530 585993
rect 176474 585919 176530 585928
rect 176290 579456 176346 579465
rect 176290 579391 176346 579400
rect 176198 553208 176254 553217
rect 176198 553143 176254 553152
rect 176304 534041 176332 579391
rect 176382 575512 176438 575521
rect 176382 575447 176438 575456
rect 176396 560561 176424 575447
rect 176382 560552 176438 560561
rect 176382 560487 176438 560496
rect 176488 559745 176516 585919
rect 176474 559736 176530 559745
rect 176474 559671 176530 559680
rect 176580 558657 176608 589319
rect 177118 569936 177174 569945
rect 177118 569871 177174 569880
rect 176566 558648 176622 558657
rect 176566 558583 176622 558592
rect 177132 548554 177160 569871
rect 177224 559570 177252 610671
rect 177212 559564 177264 559570
rect 177212 559506 177264 559512
rect 177316 549914 177344 612711
rect 177946 611688 178002 611697
rect 177946 611623 178002 611632
rect 177670 611416 177726 611425
rect 177670 611351 177726 611360
rect 177394 607064 177450 607073
rect 177394 606999 177450 607008
rect 177578 607064 177634 607073
rect 177578 606999 177634 607008
rect 177304 549908 177356 549914
rect 177304 549850 177356 549856
rect 177120 548548 177172 548554
rect 177120 548490 177172 548496
rect 177408 543046 177436 606999
rect 177592 605834 177620 606999
rect 177500 605806 177620 605834
rect 177396 543040 177448 543046
rect 177396 542982 177448 542988
rect 177500 540326 177528 605806
rect 177578 601760 177634 601769
rect 177578 601695 177634 601704
rect 177488 540320 177540 540326
rect 177488 540262 177540 540268
rect 176290 534032 176346 534041
rect 176290 533967 176346 533976
rect 177592 533458 177620 601695
rect 177580 533452 177632 533458
rect 177580 533394 177632 533400
rect 177684 530602 177712 611351
rect 177854 609784 177910 609793
rect 177854 609719 177910 609728
rect 177762 604480 177818 604489
rect 177762 604415 177818 604424
rect 177672 530596 177724 530602
rect 177672 530538 177724 530544
rect 177776 530482 177804 604415
rect 177592 530454 177804 530482
rect 177486 529408 177542 529417
rect 177486 529343 177542 529352
rect 177500 528630 177528 529343
rect 177488 528624 177540 528630
rect 177488 528566 177540 528572
rect 176106 525464 176162 525473
rect 176106 525399 176162 525408
rect 177592 523025 177620 530454
rect 177868 528554 177896 609719
rect 177684 528526 177896 528554
rect 176934 523016 176990 523025
rect 176934 522951 176990 522960
rect 177578 523016 177634 523025
rect 177578 522951 177634 522960
rect 176014 522744 176070 522753
rect 176014 522679 176070 522688
rect 175922 522200 175978 522209
rect 175922 522135 175978 522144
rect 175936 520849 175964 522135
rect 175922 520840 175978 520849
rect 175922 520775 175978 520784
rect 176948 518106 176976 522951
rect 177684 522209 177712 528526
rect 177670 522200 177726 522209
rect 177670 522135 177726 522144
rect 177960 519518 177988 611623
rect 178682 608016 178738 608025
rect 178682 607951 178738 607960
rect 178038 601624 178094 601633
rect 178038 601559 178094 601568
rect 178052 600681 178080 601559
rect 178038 600672 178094 600681
rect 178038 600607 178094 600616
rect 178590 590880 178646 590889
rect 178590 590815 178646 590824
rect 178406 572384 178462 572393
rect 178406 572319 178462 572328
rect 178420 558249 178448 572319
rect 178498 561232 178554 561241
rect 178498 561167 178554 561176
rect 178406 558240 178462 558249
rect 178406 558175 178462 558184
rect 178038 556608 178094 556617
rect 178038 556543 178094 556552
rect 178052 556238 178080 556543
rect 178040 556232 178092 556238
rect 178040 556174 178092 556180
rect 178420 555937 178448 558175
rect 178406 555928 178462 555937
rect 178406 555863 178462 555872
rect 178038 551032 178094 551041
rect 178038 550967 178094 550976
rect 178052 550662 178080 550967
rect 178040 550656 178092 550662
rect 178040 550598 178092 550604
rect 178040 536648 178092 536654
rect 178040 536590 178092 536596
rect 178052 535673 178080 536590
rect 178038 535664 178094 535673
rect 178038 535599 178094 535608
rect 178040 532500 178092 532506
rect 178040 532442 178092 532448
rect 178052 531457 178080 532442
rect 178038 531448 178094 531457
rect 178038 531383 178094 531392
rect 178040 524068 178092 524074
rect 178040 524010 178092 524016
rect 178052 523297 178080 524010
rect 178038 523288 178094 523297
rect 178038 523223 178094 523232
rect 177948 519512 178000 519518
rect 177948 519454 178000 519460
rect 178512 518106 178540 561167
rect 178604 560658 178632 590815
rect 178592 560652 178644 560658
rect 178592 560594 178644 560600
rect 178696 532098 178724 607951
rect 178972 599593 179000 633519
rect 179064 600681 179092 635559
rect 179234 635488 179290 635497
rect 179234 635423 179290 635432
rect 179142 634536 179198 634545
rect 179142 634471 179198 634480
rect 179050 600672 179106 600681
rect 179050 600607 179106 600616
rect 178958 599584 179014 599593
rect 178958 599519 179014 599528
rect 179156 598505 179184 634471
rect 179142 598496 179198 598505
rect 179142 598431 179198 598440
rect 179248 597417 179276 635423
rect 179326 635352 179382 635361
rect 179326 635287 179382 635296
rect 179340 605169 179368 635287
rect 183112 634930 183140 637758
rect 183190 637735 183246 637744
rect 184308 634930 184336 639095
rect 185688 634930 185716 640426
rect 186608 635202 186636 645934
rect 191748 644632 191800 644638
rect 191748 644574 191800 644580
rect 189172 644564 189224 644570
rect 189172 644506 189224 644512
rect 187884 644496 187936 644502
rect 187884 644438 187936 644444
rect 187896 635202 187924 644438
rect 189184 635202 189212 644506
rect 190736 640416 190788 640422
rect 190736 640358 190788 640364
rect 182712 634902 183140 634930
rect 184000 634902 184336 634930
rect 185288 634902 185716 634930
rect 186562 635174 186636 635202
rect 187850 635174 187924 635202
rect 189138 635174 189212 635202
rect 186562 634916 186590 635174
rect 187850 634916 187878 635174
rect 189138 634916 189166 635174
rect 190748 634930 190776 640358
rect 191760 635202 191788 644574
rect 193048 635202 193076 648207
rect 202050 647592 202106 647601
rect 202050 647527 202106 647536
rect 194324 645924 194376 645930
rect 194324 645866 194376 645872
rect 194336 635202 194364 645866
rect 199750 640112 199806 640121
rect 199750 640047 199806 640056
rect 198646 639568 198702 639577
rect 198568 639526 198646 639554
rect 197266 639024 197322 639033
rect 197266 638959 197322 638968
rect 195886 637664 195942 637673
rect 195886 637599 195942 637608
rect 190440 634902 190776 634930
rect 191714 635174 191788 635202
rect 193002 635174 193076 635202
rect 194290 635174 194364 635202
rect 191714 634916 191742 635174
rect 193002 634916 193030 635174
rect 194290 634916 194318 635174
rect 195900 634930 195928 637599
rect 197280 634930 197308 638959
rect 198568 634930 198596 639526
rect 198646 639503 198702 639512
rect 199764 634930 199792 640047
rect 201130 635760 201186 635769
rect 201130 635695 201186 635704
rect 201144 634930 201172 635695
rect 202064 635202 202092 647527
rect 204916 647494 204944 648343
rect 208398 648272 208454 648281
rect 208398 648207 208454 648216
rect 204904 647488 204956 647494
rect 202786 647456 202842 647465
rect 204904 647430 204956 647436
rect 202786 647391 202788 647400
rect 202840 647391 202842 647400
rect 202788 647362 202840 647368
rect 204626 647320 204682 647329
rect 208412 647290 208440 648207
rect 208490 647456 208546 647465
rect 208490 647391 208546 647400
rect 204626 647255 204682 647264
rect 208400 647284 208452 647290
rect 204166 643648 204222 643657
rect 204166 643583 204222 643592
rect 203798 643240 203854 643249
rect 195592 634902 195928 634930
rect 196880 634902 197308 634930
rect 198168 634902 198596 634930
rect 199456 634902 199792 634930
rect 200744 634902 201172 634930
rect 202018 635174 202092 635202
rect 203720 643198 203798 643226
rect 202018 634916 202046 635174
rect 203720 634930 203748 643198
rect 204180 643210 204208 643583
rect 203798 643175 203854 643184
rect 204168 643204 204220 643210
rect 204168 643146 204220 643152
rect 204640 635202 204668 647255
rect 208400 647226 208452 647232
rect 207478 643648 207534 643657
rect 207478 643583 207534 643592
rect 207020 643476 207072 643482
rect 207020 643418 207072 643424
rect 207032 643249 207060 643418
rect 207018 643240 207074 643249
rect 207018 643175 207074 643184
rect 206374 639976 206430 639985
rect 203320 634902 203748 634930
rect 204594 635174 204668 635202
rect 206296 639934 206374 639962
rect 204594 634916 204622 635174
rect 206296 634930 206324 639934
rect 206374 639911 206430 639920
rect 207492 634930 207520 643583
rect 208504 635202 208532 647391
rect 212354 646912 212410 646921
rect 212354 646847 212410 646856
rect 211068 640552 211120 640558
rect 211068 640494 211120 640500
rect 210146 638616 210202 638625
rect 210146 638551 210202 638560
rect 205896 634902 206324 634930
rect 207184 634902 207520 634930
rect 208458 635174 208532 635202
rect 208458 634916 208486 635174
rect 210160 634930 210188 638551
rect 211080 638330 211108 640494
rect 210988 638302 211108 638330
rect 210988 635202 211016 638302
rect 211068 638240 211120 638246
rect 211068 638182 211120 638188
rect 211080 637809 211108 638182
rect 211066 637800 211122 637809
rect 211066 637735 211122 637744
rect 212368 635202 212396 646847
rect 212446 646776 212502 646785
rect 212446 646711 212502 646720
rect 212460 646066 212488 646711
rect 232516 646542 232544 668578
rect 235184 657529 235212 703520
rect 267660 700330 267688 703520
rect 257344 700324 257396 700330
rect 257344 700266 257396 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 257356 687954 257384 700266
rect 247684 687948 247736 687954
rect 247684 687890 247736 687896
rect 257344 687948 257396 687954
rect 257344 687890 257396 687896
rect 247696 676190 247724 687890
rect 283852 681737 283880 703520
rect 283838 681728 283894 681737
rect 283838 681663 283894 681672
rect 288346 681728 288402 681737
rect 288346 681663 288402 681672
rect 288360 678745 288388 681663
rect 288346 678736 288402 678745
rect 288346 678671 288402 678680
rect 290462 678736 290518 678745
rect 290462 678671 290518 678680
rect 244556 676184 244608 676190
rect 244556 676126 244608 676132
rect 247684 676184 247736 676190
rect 247684 676126 247736 676132
rect 244568 668642 244596 676126
rect 244556 668636 244608 668642
rect 244556 668578 244608 668584
rect 290476 657801 290504 678671
rect 290462 657792 290518 657801
rect 290462 657727 290518 657736
rect 298744 657688 298796 657694
rect 300136 657665 300164 703520
rect 332520 694822 332548 703520
rect 348804 700330 348832 703520
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 332508 694816 332560 694822
rect 332508 694758 332560 694764
rect 338764 694816 338816 694822
rect 338764 694758 338816 694764
rect 338776 682446 338804 694758
rect 338764 682440 338816 682446
rect 338764 682382 338816 682388
rect 358728 682440 358780 682446
rect 358728 682382 358780 682388
rect 358740 680338 358768 682382
rect 358728 680332 358780 680338
rect 358728 680274 358780 680280
rect 309782 657792 309838 657801
rect 309782 657727 309838 657736
rect 298744 657630 298796 657636
rect 300122 657656 300178 657665
rect 235170 657520 235226 657529
rect 235170 657455 235226 657464
rect 280802 648136 280858 648145
rect 280802 648071 280858 648080
rect 275282 647728 275338 647737
rect 275282 647663 275338 647672
rect 233146 647592 233202 647601
rect 233422 647592 233478 647601
rect 233146 647527 233202 647536
rect 233252 647550 233422 647578
rect 233160 647358 233188 647527
rect 233148 647352 233200 647358
rect 233148 647294 233200 647300
rect 233252 647170 233280 647550
rect 233422 647527 233478 647536
rect 232976 647142 233280 647170
rect 222844 646536 222896 646542
rect 222844 646478 222896 646484
rect 232504 646536 232556 646542
rect 232504 646478 232556 646484
rect 212448 646060 212500 646066
rect 212448 646002 212500 646008
rect 216218 645552 216274 645561
rect 216218 645487 216274 645496
rect 215300 644972 215352 644978
rect 215300 644914 215352 644920
rect 215312 644881 215340 644914
rect 215298 644872 215354 644881
rect 215298 644807 215354 644816
rect 214564 640824 214616 640830
rect 214564 640766 214616 640772
rect 214576 640393 214604 640766
rect 214562 640384 214618 640393
rect 214562 640319 214618 640328
rect 215206 640384 215262 640393
rect 215206 640319 215262 640328
rect 213826 639296 213882 639305
rect 210988 635174 211062 635202
rect 209760 634902 210188 634930
rect 211034 634916 211062 635174
rect 212322 635174 212396 635202
rect 213748 639254 213826 639282
rect 212322 634916 212350 635174
rect 213748 634930 213776 639254
rect 213826 639231 213882 639240
rect 213826 639160 213882 639169
rect 213826 639095 213882 639104
rect 213840 638994 213868 639095
rect 213828 638988 213880 638994
rect 213828 638930 213880 638936
rect 215220 634930 215248 640319
rect 216232 635202 216260 645487
rect 218058 641472 218114 641481
rect 218058 641407 218114 641416
rect 218072 640898 218100 641407
rect 218060 640892 218112 640898
rect 218060 640834 218112 640840
rect 217966 640792 218022 640801
rect 217888 640750 217966 640778
rect 216772 640620 216824 640626
rect 216772 640562 216824 640568
rect 216784 640393 216812 640562
rect 216770 640384 216826 640393
rect 216770 640319 216826 640328
rect 213624 634902 213776 634930
rect 214912 634902 215248 634930
rect 216186 635174 216260 635202
rect 216186 634916 216214 635174
rect 217888 634930 217916 640750
rect 217966 640727 218022 640736
rect 219070 640656 219126 640665
rect 219070 640591 219126 640600
rect 219084 634930 219112 640591
rect 220728 639600 220780 639606
rect 220728 639542 220780 639548
rect 220358 639296 220414 639305
rect 220358 639231 220414 639240
rect 220372 634930 220400 639231
rect 220740 639033 220768 639542
rect 220726 639024 220782 639033
rect 220726 638959 220782 638968
rect 221830 636576 221886 636585
rect 221752 636534 221830 636562
rect 221752 634930 221780 636534
rect 221830 636511 221886 636520
rect 222856 635594 222884 646478
rect 227718 645552 227774 645561
rect 227718 645487 227774 645496
rect 227732 644774 227760 645487
rect 231766 645008 231822 645017
rect 232042 645008 232098 645017
rect 231766 644943 231822 644952
rect 231872 644966 232042 644994
rect 231780 644910 231808 644943
rect 231768 644904 231820 644910
rect 227810 644872 227866 644881
rect 231768 644846 231820 644852
rect 227810 644807 227866 644816
rect 227720 644768 227772 644774
rect 227720 644710 227772 644716
rect 223486 642832 223542 642841
rect 223486 642767 223542 642776
rect 223500 642258 223528 642767
rect 223488 642252 223540 642258
rect 223488 642194 223540 642200
rect 222934 641880 222990 641889
rect 222934 641815 222990 641824
rect 222844 635588 222896 635594
rect 222844 635530 222896 635536
rect 222948 634930 222976 641815
rect 224224 637832 224276 637838
rect 224224 637774 224276 637780
rect 224314 637800 224370 637809
rect 224236 637673 224264 637774
rect 224314 637735 224370 637744
rect 224222 637664 224278 637673
rect 224222 637599 224278 637608
rect 224328 634930 224356 637735
rect 225694 636304 225750 636313
rect 225616 636262 225694 636290
rect 225616 634930 225644 636262
rect 225694 636239 225750 636248
rect 227824 635202 227852 644807
rect 231872 644722 231900 644966
rect 232042 644943 232098 644952
rect 231688 644694 231900 644722
rect 230386 640792 230442 640801
rect 230662 640792 230718 640801
rect 230386 640727 230442 640736
rect 230492 640750 230662 640778
rect 230400 640694 230428 640727
rect 230388 640688 230440 640694
rect 230388 640630 230440 640636
rect 230492 640506 230520 640750
rect 230662 640727 230718 640736
rect 230308 640478 230520 640506
rect 229558 637664 229614 637673
rect 227778 635174 227852 635202
rect 229480 637622 229558 637650
rect 226338 635080 226394 635089
rect 226338 635015 226340 635024
rect 226392 635015 226394 635024
rect 226340 634986 226392 634992
rect 217488 634902 217916 634930
rect 218776 634902 219112 634930
rect 220064 634902 220400 634930
rect 221352 634902 221780 634930
rect 222640 634902 222976 634930
rect 223928 634902 224356 634930
rect 225216 634902 225644 634930
rect 226476 634944 226532 634953
rect 227778 634916 227806 635174
rect 229480 634930 229508 637622
rect 229558 637599 229614 637608
rect 230308 635202 230336 640478
rect 230386 638616 230442 638625
rect 230386 638551 230442 638560
rect 230400 637770 230428 638551
rect 230388 637764 230440 637770
rect 230388 637706 230440 637712
rect 231688 635202 231716 644694
rect 232976 635202 233004 647142
rect 233882 643648 233938 643657
rect 233882 643583 233938 643592
rect 234526 643648 234582 643657
rect 234526 643583 234582 643592
rect 233896 643550 233924 643583
rect 233884 643544 233936 643550
rect 233884 643486 233936 643492
rect 230308 635174 230382 635202
rect 229080 634902 229508 634930
rect 230354 634916 230382 635174
rect 231642 635174 231716 635202
rect 232930 635174 233004 635202
rect 231642 634916 231670 635174
rect 232930 634916 232958 635174
rect 234540 634930 234568 643583
rect 249708 641776 249760 641782
rect 249708 641718 249760 641724
rect 234618 639568 234674 639577
rect 234618 639503 234674 639512
rect 235906 639568 235962 639577
rect 235906 639503 235962 639512
rect 234632 639062 234660 639503
rect 234620 639056 234672 639062
rect 234620 638998 234672 639004
rect 235920 634930 235948 639503
rect 247500 637900 247552 637906
rect 247500 637842 247552 637848
rect 245014 637256 245070 637265
rect 244936 637214 245014 637242
rect 241060 637016 241112 637022
rect 241060 636958 241112 636964
rect 238392 636812 238444 636818
rect 238392 636754 238444 636760
rect 237104 636540 237156 636546
rect 237104 636482 237156 636488
rect 237116 634930 237144 636482
rect 238404 634930 238432 636754
rect 239680 636608 239732 636614
rect 239680 636550 239732 636556
rect 239692 634930 239720 636550
rect 241072 634930 241100 636958
rect 243636 636676 243688 636682
rect 243636 636618 243688 636624
rect 243648 634930 243676 636618
rect 244278 635760 244334 635769
rect 244278 635695 244334 635704
rect 244292 635118 244320 635695
rect 244280 635112 244332 635118
rect 244280 635054 244332 635060
rect 244936 634930 244964 637214
rect 245014 637191 245070 637200
rect 247512 634930 247540 637842
rect 249614 637256 249670 637265
rect 249614 637191 249670 637200
rect 249628 636886 249656 637191
rect 249616 636880 249668 636886
rect 249616 636822 249668 636828
rect 248786 636304 248842 636313
rect 249720 636274 249748 641718
rect 251086 640112 251142 640121
rect 251086 640047 251142 640056
rect 250994 639840 251050 639849
rect 250994 639775 251050 639784
rect 251008 638489 251036 639775
rect 251100 639334 251128 640047
rect 251088 639328 251140 639334
rect 251088 639270 251140 639276
rect 250994 638480 251050 638489
rect 250994 638415 251050 638424
rect 248786 636239 248842 636248
rect 249708 636268 249760 636274
rect 248800 634930 248828 636239
rect 249708 636210 249760 636216
rect 249720 635202 249748 636210
rect 251008 635202 251036 638415
rect 273996 636948 274048 636954
rect 273996 636890 274048 636896
rect 268384 636880 268436 636886
rect 268384 636822 268436 636828
rect 254582 636712 254638 636721
rect 254582 636647 254638 636656
rect 252466 636168 252522 636177
rect 252466 636103 252522 636112
rect 252480 635254 252508 636103
rect 234232 634902 234568 634930
rect 235520 634902 235948 634930
rect 236808 634902 237144 634930
rect 238096 634902 238432 634930
rect 239384 634902 239720 634930
rect 240672 634902 241100 634930
rect 243248 634902 243676 634930
rect 244536 634902 244964 634930
rect 247112 634902 247540 634930
rect 248400 634902 248828 634930
rect 249674 635174 249748 635202
rect 250962 635174 251036 635202
rect 252468 635248 252520 635254
rect 252468 635190 252520 635196
rect 249674 634916 249702 635174
rect 250962 634916 250990 635174
rect 252466 635080 252522 635089
rect 252466 635015 252522 635024
rect 252480 634930 252508 635015
rect 252264 634902 252508 634930
rect 226476 634879 226532 634888
rect 246132 634846 246160 634877
rect 246120 634840 246172 634846
rect 245824 634788 246120 634794
rect 245824 634782 246172 634788
rect 245824 634766 246160 634782
rect 241923 634208 241932 634264
rect 241988 634208 241997 634264
rect 179326 605160 179382 605169
rect 179326 605095 179382 605104
rect 179234 597408 179290 597417
rect 179234 597343 179290 597352
rect 179340 596329 179368 605095
rect 179326 596320 179382 596329
rect 179326 596255 179382 596264
rect 179234 592512 179290 592521
rect 179234 592447 179290 592456
rect 179142 585168 179198 585177
rect 179142 585103 179198 585112
rect 178866 583536 178922 583545
rect 178866 583471 178922 583480
rect 178774 577688 178830 577697
rect 178774 577623 178830 577632
rect 178684 532092 178736 532098
rect 178684 532034 178736 532040
rect 178788 524113 178816 577623
rect 178880 532166 178908 583471
rect 179050 580272 179106 580281
rect 179050 580207 179106 580216
rect 178958 578640 179014 578649
rect 178958 578575 179014 578584
rect 178972 532681 179000 578575
rect 179064 536761 179092 580207
rect 179156 551721 179184 585103
rect 179248 560386 179276 592447
rect 179326 588704 179382 588713
rect 179326 588639 179382 588648
rect 179236 560380 179288 560386
rect 179236 560322 179288 560328
rect 179234 560280 179290 560289
rect 179234 560215 179290 560224
rect 179142 551712 179198 551721
rect 179142 551647 179198 551656
rect 179050 536752 179106 536761
rect 179050 536687 179106 536696
rect 179248 534818 179276 560215
rect 179340 556617 179368 588639
rect 179878 581088 179934 581097
rect 179878 581023 179934 581032
rect 179892 576854 179920 581023
rect 179892 576826 180012 576854
rect 179878 574560 179934 574569
rect 179878 574495 179934 574504
rect 179786 573472 179842 573481
rect 179786 573407 179842 573416
rect 179602 562184 179658 562193
rect 179602 562119 179658 562128
rect 179418 561640 179474 561649
rect 179418 561575 179474 561584
rect 179432 560590 179460 561575
rect 179420 560584 179472 560590
rect 179420 560526 179472 560532
rect 179512 560380 179564 560386
rect 179512 560322 179564 560328
rect 179524 559609 179552 560322
rect 179510 559600 179566 559609
rect 179510 559535 179566 559544
rect 179326 556608 179382 556617
rect 179326 556543 179382 556552
rect 179420 553172 179472 553178
rect 179420 553114 179472 553120
rect 179432 552129 179460 553114
rect 179418 552120 179474 552129
rect 179418 552055 179474 552064
rect 179420 550452 179472 550458
rect 179420 550394 179472 550400
rect 179432 549545 179460 550394
rect 179418 549536 179474 549545
rect 179418 549471 179474 549480
rect 179616 536110 179644 562119
rect 179694 560960 179750 560969
rect 179694 560895 179750 560904
rect 179604 536104 179656 536110
rect 179604 536046 179656 536052
rect 179236 534812 179288 534818
rect 179236 534754 179288 534760
rect 178958 532672 179014 532681
rect 178958 532607 179014 532616
rect 178868 532160 178920 532166
rect 178868 532102 178920 532108
rect 178774 524104 178830 524113
rect 178774 524039 178830 524048
rect 179708 521665 179736 560895
rect 179800 552809 179828 573407
rect 179786 552800 179842 552809
rect 179786 552735 179842 552744
rect 179892 549817 179920 574495
rect 179984 555801 180012 576826
rect 254596 561649 254624 636647
rect 262862 636304 262918 636313
rect 262862 636239 262918 636248
rect 256146 635896 256202 635905
rect 256146 635831 256202 635840
rect 255962 635216 256018 635225
rect 255962 635151 256018 635160
rect 254582 561640 254638 561649
rect 254582 561575 254638 561584
rect 229742 560552 229798 560561
rect 229742 560487 229798 560496
rect 181502 559858 181530 560116
rect 182514 559858 182542 560116
rect 183526 559858 183554 560116
rect 184538 559858 184566 560116
rect 185550 559858 185578 560116
rect 186562 559858 186590 560116
rect 187574 559858 187602 560116
rect 188586 559858 188614 560116
rect 189598 559858 189626 560116
rect 190624 560102 190960 560130
rect 181502 559830 181576 559858
rect 182514 559830 182588 559858
rect 183526 559830 183600 559858
rect 184538 559830 184612 559858
rect 185550 559830 185624 559858
rect 186562 559830 186636 559858
rect 187574 559830 187648 559858
rect 188586 559830 188660 559858
rect 189598 559830 189672 559858
rect 179970 555792 180026 555801
rect 179970 555727 180026 555736
rect 179878 549808 179934 549817
rect 179878 549743 179934 549752
rect 180062 532128 180118 532137
rect 180062 532063 180118 532072
rect 179694 521656 179750 521665
rect 179694 521591 179750 521600
rect 180076 518106 180104 532063
rect 181548 529242 181576 559830
rect 182560 541686 182588 559830
rect 183190 553888 183246 553897
rect 183190 553823 183246 553832
rect 182548 541680 182600 541686
rect 182548 541622 182600 541628
rect 181626 533760 181682 533769
rect 181626 533695 181682 533704
rect 181536 529236 181588 529242
rect 181536 529178 181588 529184
rect 180246 525736 180302 525745
rect 180246 525671 180302 525680
rect 180260 524550 180288 525671
rect 180248 524544 180300 524550
rect 180248 524486 180300 524492
rect 181640 518106 181668 533695
rect 183204 518106 183232 553823
rect 183572 540258 183600 559830
rect 183560 540252 183612 540258
rect 183560 540194 183612 540200
rect 184584 533769 184612 559830
rect 185596 534449 185624 559830
rect 184754 534440 184810 534449
rect 184754 534375 184810 534384
rect 185582 534440 185638 534449
rect 185582 534375 185638 534384
rect 184570 533760 184626 533769
rect 184570 533695 184626 533704
rect 184768 518106 184796 534375
rect 186608 527882 186636 559830
rect 187620 541754 187648 559830
rect 188632 547194 188660 559830
rect 188620 547188 188672 547194
rect 188620 547130 188672 547136
rect 189644 546378 189672 559830
rect 190932 553897 190960 560102
rect 191622 559858 191650 560116
rect 192634 559858 192662 560116
rect 193646 559858 193674 560116
rect 194658 559858 194686 560116
rect 195684 560102 195836 560130
rect 191622 559830 191696 559858
rect 192634 559830 192708 559858
rect 193646 559830 193720 559858
rect 194658 559830 194732 559858
rect 190918 553888 190974 553897
rect 190918 553823 190974 553832
rect 189632 546372 189684 546378
rect 189632 546314 189684 546320
rect 187882 543144 187938 543153
rect 187882 543079 187938 543088
rect 187608 541748 187660 541754
rect 187608 541690 187660 541696
rect 186596 527876 186648 527882
rect 186596 527818 186648 527824
rect 186226 521520 186282 521529
rect 186226 521455 186282 521464
rect 162780 518078 162824 518106
rect 140900 517956 140928 518078
rect 142464 517956 142492 518078
rect 144028 517956 144056 518078
rect 145592 517956 145620 518078
rect 147156 517956 147184 518078
rect 148720 517956 148748 518078
rect 150284 517956 150312 518078
rect 151848 517956 151876 518078
rect 153412 517956 153440 518078
rect 154976 517956 155004 518078
rect 156540 517956 156568 518078
rect 158104 517956 158132 518078
rect 159668 517956 159696 518078
rect 161232 517956 161260 518078
rect 162796 517956 162824 518078
rect 164360 518078 164464 518106
rect 165924 518078 166028 518106
rect 167488 518078 167592 518106
rect 169052 518078 169156 518106
rect 170616 518078 170720 518106
rect 172180 518078 172284 518106
rect 173744 518078 173848 518106
rect 175308 518078 175412 518106
rect 176872 518078 176976 518106
rect 178436 518078 178540 518106
rect 180000 518078 180104 518106
rect 181564 518078 181668 518106
rect 183128 518078 183232 518106
rect 184692 518078 184796 518106
rect 186240 518106 186268 521455
rect 187896 518106 187924 543079
rect 191010 536208 191066 536217
rect 191010 536143 191066 536152
rect 189446 531992 189502 532001
rect 189446 531927 189502 531936
rect 189460 518106 189488 531927
rect 191024 518106 191052 536143
rect 191668 533882 191696 559830
rect 192574 552936 192630 552945
rect 192574 552871 192630 552880
rect 191668 533854 191880 533882
rect 191746 533760 191802 533769
rect 191852 533746 191880 533854
rect 191930 533760 191986 533769
rect 191852 533718 191930 533746
rect 191746 533695 191802 533704
rect 191930 533695 191986 533704
rect 191760 532778 191788 533695
rect 191748 532772 191800 532778
rect 191748 532714 191800 532720
rect 192588 518106 192616 552871
rect 192680 536217 192708 559830
rect 192666 536208 192722 536217
rect 192666 536143 192722 536152
rect 193692 535401 193720 559830
rect 194138 551304 194194 551313
rect 194138 551239 194194 551248
rect 193678 535392 193734 535401
rect 193678 535327 193734 535336
rect 194152 518106 194180 551239
rect 194704 538898 194732 559830
rect 195702 549944 195758 549953
rect 195702 549879 195758 549888
rect 194692 538892 194744 538898
rect 194692 538834 194744 538840
rect 194506 534440 194562 534449
rect 194506 534375 194562 534384
rect 194520 534138 194548 534375
rect 194508 534132 194560 534138
rect 194508 534074 194560 534080
rect 195716 518106 195744 549879
rect 195808 537538 195836 560102
rect 196682 559858 196710 560116
rect 197694 559858 197722 560116
rect 198706 559858 198734 560116
rect 199718 559858 199746 560116
rect 200730 559858 200758 560116
rect 201742 559858 201770 560116
rect 202754 559858 202782 560116
rect 203766 559858 203794 560116
rect 204778 559858 204806 560116
rect 205804 560102 206140 560130
rect 196682 559830 196756 559858
rect 197694 559830 197768 559858
rect 198706 559830 198780 559858
rect 199718 559830 199792 559858
rect 200730 559830 200804 559858
rect 201742 559830 201816 559858
rect 202754 559830 202828 559858
rect 203766 559830 203840 559858
rect 204778 559830 204852 559858
rect 196728 541822 196756 559830
rect 196716 541816 196768 541822
rect 196716 541758 196768 541764
rect 195796 537532 195848 537538
rect 195796 537474 195848 537480
rect 197740 531729 197768 559830
rect 198752 532001 198780 559830
rect 199764 544406 199792 559830
rect 199752 544400 199804 544406
rect 199752 544342 199804 544348
rect 200776 543153 200804 559830
rect 200762 543144 200818 543153
rect 200762 543079 200818 543088
rect 198738 531992 198794 532001
rect 198738 531927 198794 531936
rect 197726 531720 197782 531729
rect 197726 531655 197782 531664
rect 200394 527096 200450 527105
rect 200394 527031 200450 527040
rect 197266 525600 197322 525609
rect 197266 525535 197322 525544
rect 197280 518106 197308 525535
rect 198830 525328 198886 525337
rect 198830 525263 198886 525272
rect 198844 518106 198872 525263
rect 200408 518106 200436 527031
rect 201788 526153 201816 559830
rect 202800 548622 202828 559830
rect 202788 548616 202840 548622
rect 202788 548558 202840 548564
rect 203812 537606 203840 559830
rect 204824 550225 204852 559830
rect 206112 551313 206140 560102
rect 206802 559858 206830 560116
rect 207814 559858 207842 560116
rect 208826 559858 208854 560116
rect 209838 559858 209866 560116
rect 210850 559858 210878 560116
rect 211862 559858 211890 560116
rect 212874 559858 212902 560116
rect 213886 559858 213914 560116
rect 214898 559858 214926 560116
rect 215910 559858 215938 560116
rect 216922 559858 216950 560116
rect 217934 559858 217962 560116
rect 218946 559858 218974 560116
rect 219958 559858 219986 560116
rect 220970 559858 220998 560116
rect 221982 559858 222010 560116
rect 222994 559858 223022 560116
rect 224006 559858 224034 560116
rect 225018 559858 225046 560116
rect 226030 559858 226058 560116
rect 227042 559858 227070 560116
rect 228068 560102 228404 560130
rect 229080 560102 229416 560130
rect 206802 559830 206876 559858
rect 207814 559830 207888 559858
rect 208826 559830 208900 559858
rect 209838 559830 209912 559858
rect 210850 559830 210924 559858
rect 211862 559830 211936 559858
rect 212874 559830 212948 559858
rect 213886 559830 213960 559858
rect 214898 559830 214972 559858
rect 215910 559830 215984 559858
rect 216922 559830 216996 559858
rect 217934 559830 218008 559858
rect 218946 559830 219020 559858
rect 219958 559830 220032 559858
rect 220970 559830 221044 559858
rect 221982 559830 222056 559858
rect 222994 559830 223068 559858
rect 224006 559830 224080 559858
rect 225018 559830 225092 559858
rect 226030 559830 226104 559858
rect 227042 559830 227116 559858
rect 206098 551304 206154 551313
rect 206098 551239 206154 551248
rect 204810 550216 204866 550225
rect 204810 550151 204866 550160
rect 203800 537600 203852 537606
rect 203800 537542 203852 537548
rect 206848 536217 206876 559830
rect 207860 545766 207888 559830
rect 207848 545760 207900 545766
rect 207848 545702 207900 545708
rect 208872 540462 208900 559830
rect 208860 540456 208912 540462
rect 208860 540398 208912 540404
rect 209884 538966 209912 559830
rect 209872 538960 209924 538966
rect 209872 538902 209924 538908
rect 210896 538214 210924 559830
rect 210896 538186 211108 538214
rect 205638 536208 205694 536217
rect 205638 536143 205694 536152
rect 206834 536208 206890 536217
rect 206834 536143 206890 536152
rect 205652 535498 205680 536143
rect 205640 535492 205692 535498
rect 205640 535434 205692 535440
rect 211080 531457 211108 538186
rect 211908 534449 211936 559830
rect 212446 535392 212502 535401
rect 212446 535327 212502 535336
rect 211894 534440 211950 534449
rect 211894 534375 211950 534384
rect 212460 534206 212488 535327
rect 212448 534200 212500 534206
rect 212448 534142 212500 534148
rect 212920 532137 212948 559830
rect 213932 541385 213960 559830
rect 214470 541784 214526 541793
rect 214470 541719 214526 541728
rect 213918 541376 213974 541385
rect 213918 541311 213974 541320
rect 212906 532128 212962 532137
rect 212906 532063 212962 532072
rect 213826 531720 213882 531729
rect 213826 531655 213882 531664
rect 211066 531448 211122 531457
rect 211066 531383 211122 531392
rect 213840 531350 213868 531655
rect 213828 531344 213880 531350
rect 211066 531312 211122 531321
rect 213828 531286 213880 531292
rect 211066 531247 211122 531256
rect 211080 531010 211108 531247
rect 211068 531004 211120 531010
rect 211068 530946 211120 530952
rect 212906 530904 212962 530913
rect 212906 530839 212962 530848
rect 203522 526960 203578 526969
rect 203522 526895 203578 526904
rect 201958 526280 202014 526289
rect 201958 526215 202014 526224
rect 201774 526144 201830 526153
rect 201774 526079 201830 526088
rect 201972 518106 202000 526215
rect 203536 518106 203564 526895
rect 205086 526824 205142 526833
rect 205086 526759 205142 526768
rect 205100 518106 205128 526759
rect 206650 526688 206706 526697
rect 206650 526623 206706 526632
rect 206664 518106 206692 526623
rect 208214 526552 208270 526561
rect 208214 526487 208270 526496
rect 211344 526516 211396 526522
rect 208228 518106 208256 526487
rect 211344 526458 211396 526464
rect 209686 526416 209742 526425
rect 209686 526351 209742 526360
rect 186240 518078 186284 518106
rect 164360 517956 164388 518078
rect 165924 517956 165952 518078
rect 167488 517956 167516 518078
rect 169052 517956 169080 518078
rect 170616 517956 170644 518078
rect 172180 517956 172208 518078
rect 173744 517956 173772 518078
rect 175308 517956 175336 518078
rect 176872 517956 176900 518078
rect 178436 517956 178464 518078
rect 180000 517956 180028 518078
rect 181564 517956 181592 518078
rect 183128 517956 183156 518078
rect 184692 517956 184720 518078
rect 186256 517956 186284 518078
rect 187820 518078 187924 518106
rect 189384 518078 189488 518106
rect 190948 518078 191052 518106
rect 192512 518078 192616 518106
rect 194076 518078 194180 518106
rect 195640 518078 195744 518106
rect 197204 518078 197308 518106
rect 198768 518078 198872 518106
rect 200332 518078 200436 518106
rect 201896 518078 202000 518106
rect 203460 518078 203564 518106
rect 205024 518078 205128 518106
rect 206588 518078 206692 518106
rect 208152 518078 208256 518106
rect 209700 518106 209728 526351
rect 211066 524920 211122 524929
rect 211066 524855 211122 524864
rect 211080 521529 211108 524855
rect 211066 521520 211122 521529
rect 211066 521455 211122 521464
rect 211356 518106 211384 526458
rect 212920 518106 212948 530839
rect 214484 518106 214512 541719
rect 214944 526561 214972 559830
rect 215956 544474 215984 559830
rect 216128 557728 216180 557734
rect 216128 557670 216180 557676
rect 215944 544468 215996 544474
rect 215944 544410 215996 544416
rect 214930 526552 214986 526561
rect 214930 526487 214986 526496
rect 216140 521150 216168 557670
rect 216680 547664 216732 547670
rect 216680 547606 216732 547612
rect 216692 546553 216720 547606
rect 216968 547097 216996 559830
rect 216954 547088 217010 547097
rect 216954 547023 217010 547032
rect 216678 546544 216734 546553
rect 216678 546479 216734 546488
rect 217980 526425 218008 559830
rect 218992 536217 219020 559830
rect 218058 536208 218114 536217
rect 218058 536143 218114 536152
rect 218978 536208 219034 536217
rect 218978 536143 219034 536152
rect 218072 535634 218100 536143
rect 218060 535628 218112 535634
rect 218060 535570 218112 535576
rect 218702 532400 218758 532409
rect 218702 532335 218758 532344
rect 217966 526416 218022 526425
rect 217966 526351 218022 526360
rect 218716 521393 218744 532335
rect 220004 527921 220032 559830
rect 220726 532264 220782 532273
rect 220726 532199 220782 532208
rect 220636 528420 220688 528426
rect 220636 528362 220688 528368
rect 219990 527912 220046 527921
rect 219990 527847 220046 527856
rect 220648 527377 220676 528362
rect 220634 527368 220690 527377
rect 220634 527303 220690 527312
rect 217506 521384 217562 521393
rect 217506 521319 217562 521328
rect 218702 521384 218758 521393
rect 218702 521319 218758 521328
rect 216128 521144 216180 521150
rect 216128 521086 216180 521092
rect 215942 520840 215998 520849
rect 215942 520775 215998 520784
rect 209700 518078 209744 518106
rect 187820 517956 187848 518078
rect 189384 517956 189412 518078
rect 190948 517956 190976 518078
rect 192512 517956 192540 518078
rect 194076 517956 194104 518078
rect 195640 517956 195668 518078
rect 197204 517956 197232 518078
rect 198768 517956 198796 518078
rect 200332 517956 200360 518078
rect 201896 517956 201924 518078
rect 203460 517956 203488 518078
rect 205024 517956 205052 518078
rect 206588 517956 206616 518078
rect 208152 517956 208180 518078
rect 209716 517956 209744 518078
rect 211280 518078 211384 518106
rect 212844 518078 212948 518106
rect 214408 518078 214512 518106
rect 215956 518106 215984 520775
rect 217520 518106 217548 521319
rect 219070 521248 219126 521257
rect 219070 521183 219126 521192
rect 219084 518106 219112 521183
rect 220740 518106 220768 532199
rect 221016 530913 221044 559830
rect 221002 530904 221058 530913
rect 221002 530839 221058 530848
rect 222028 526697 222056 559830
rect 223040 545873 223068 559830
rect 223488 546100 223540 546106
rect 223488 546042 223540 546048
rect 223026 545864 223082 545873
rect 223026 545799 223082 545808
rect 223500 545193 223528 546042
rect 223486 545184 223542 545193
rect 223486 545119 223542 545128
rect 224052 541793 224080 559830
rect 224958 550216 225014 550225
rect 224958 550151 225014 550160
rect 224972 549302 225000 550151
rect 225064 549953 225092 559830
rect 225050 549944 225106 549953
rect 225050 549879 225106 549888
rect 224960 549296 225012 549302
rect 224960 549238 225012 549244
rect 226076 547262 226104 559830
rect 226064 547256 226116 547262
rect 226064 547198 226116 547204
rect 224224 542292 224276 542298
rect 224224 542234 224276 542240
rect 224038 541784 224094 541793
rect 224038 541719 224094 541728
rect 224236 541113 224264 542234
rect 224222 541104 224278 541113
rect 224222 541039 224278 541048
rect 225418 540696 225474 540705
rect 225418 540631 225474 540640
rect 222290 538928 222346 538937
rect 222290 538863 222346 538872
rect 222014 526688 222070 526697
rect 222014 526623 222070 526632
rect 222304 518106 222332 538863
rect 223854 525192 223910 525201
rect 223854 525127 223910 525136
rect 223868 518106 223896 525127
rect 225432 518106 225460 540631
rect 227088 538529 227116 559830
rect 228376 558521 228404 560102
rect 228362 558512 228418 558521
rect 228362 558447 228418 558456
rect 229388 552537 229416 560102
rect 229374 552528 229430 552537
rect 229374 552463 229430 552472
rect 229756 546825 229784 560487
rect 230078 559858 230106 560116
rect 231090 559858 231118 560116
rect 232102 559858 232130 560116
rect 233114 559858 233142 560116
rect 234126 559858 234154 560116
rect 235138 559858 235166 560116
rect 236150 559858 236178 560116
rect 237162 559858 237190 560116
rect 238174 559858 238202 560116
rect 239186 559858 239214 560116
rect 240198 559858 240226 560116
rect 241224 560102 241376 560130
rect 230078 559830 230152 559858
rect 231090 559830 231164 559858
rect 232102 559830 232176 559858
rect 233114 559830 233188 559858
rect 234126 559830 234200 559858
rect 235138 559830 235212 559858
rect 236150 559830 236224 559858
rect 237162 559830 237236 559858
rect 238174 559830 238248 559858
rect 239186 559830 239260 559858
rect 240198 559830 240272 559858
rect 229742 546816 229798 546825
rect 229742 546751 229798 546760
rect 228546 545592 228602 545601
rect 228546 545527 228602 545536
rect 227074 538520 227130 538529
rect 227074 538455 227130 538464
rect 226982 525056 227038 525065
rect 226982 524991 227038 525000
rect 226996 518106 227024 524991
rect 228560 518106 228588 545527
rect 230124 543266 230152 559830
rect 230386 547632 230442 547641
rect 230386 547567 230442 547576
rect 230400 546582 230428 547567
rect 230388 546576 230440 546582
rect 230388 546518 230440 546524
rect 230124 543238 230520 543266
rect 230386 543144 230442 543153
rect 230492 543130 230520 543238
rect 230662 543144 230718 543153
rect 230492 543102 230662 543130
rect 230386 543079 230442 543088
rect 230662 543079 230718 543088
rect 230400 542502 230428 543079
rect 230388 542496 230440 542502
rect 230388 542438 230440 542444
rect 230110 537840 230166 537849
rect 230110 537775 230166 537784
rect 230124 518106 230152 537775
rect 231136 525201 231164 559830
rect 231674 548720 231730 548729
rect 231674 548655 231730 548664
rect 231214 543280 231270 543289
rect 231214 543215 231270 543224
rect 231122 525192 231178 525201
rect 231122 525127 231178 525136
rect 231228 521257 231256 543215
rect 231214 521248 231270 521257
rect 231214 521183 231270 521192
rect 231688 518106 231716 548655
rect 232148 541929 232176 559830
rect 233160 557534 233188 559830
rect 233068 557506 233188 557534
rect 233068 550225 233096 557506
rect 233148 550316 233200 550322
rect 233148 550258 233200 550264
rect 233054 550216 233110 550225
rect 233054 550151 233110 550160
rect 233160 549409 233188 550258
rect 233146 549400 233202 549409
rect 233146 549335 233202 549344
rect 233882 546952 233938 546961
rect 233882 546887 233938 546896
rect 232134 541920 232190 541929
rect 232134 541855 232190 541864
rect 233146 541376 233202 541385
rect 233146 541311 233202 541320
rect 233160 541006 233188 541311
rect 233148 541000 233200 541006
rect 233148 540942 233200 540948
rect 233896 521257 233924 546887
rect 234172 525065 234200 559830
rect 235184 526833 235212 559830
rect 236196 537849 236224 559830
rect 237208 543289 237236 559830
rect 238220 548729 238248 559830
rect 238206 548720 238262 548729
rect 238206 548655 238262 548664
rect 237930 544640 237986 544649
rect 237930 544575 237986 544584
rect 237194 543280 237250 543289
rect 237194 543215 237250 543224
rect 236182 537840 236238 537849
rect 236182 537775 236238 537784
rect 236366 529680 236422 529689
rect 236366 529615 236422 529624
rect 235170 526824 235226 526833
rect 235170 526759 235226 526768
rect 234158 525056 234214 525065
rect 234158 524991 234214 525000
rect 233146 521248 233202 521257
rect 233146 521183 233202 521192
rect 233882 521248 233938 521257
rect 233882 521183 233938 521192
rect 234710 521248 234766 521257
rect 234710 521183 234766 521192
rect 215956 518078 216000 518106
rect 217520 518078 217564 518106
rect 219084 518078 219128 518106
rect 211280 517956 211308 518078
rect 212844 517956 212872 518078
rect 214408 517956 214436 518078
rect 215972 517956 216000 518078
rect 217536 517956 217564 518078
rect 219100 517956 219128 518078
rect 220664 518078 220768 518106
rect 222228 518078 222332 518106
rect 223792 518078 223896 518106
rect 225356 518078 225460 518106
rect 226920 518078 227024 518106
rect 228484 518078 228588 518106
rect 230048 518078 230152 518106
rect 231612 518078 231716 518106
rect 233160 518106 233188 521183
rect 234724 518106 234752 521183
rect 236380 518106 236408 529615
rect 237944 518106 237972 544575
rect 239232 540705 239260 559830
rect 239218 540696 239274 540705
rect 239218 540631 239274 540640
rect 240244 538937 240272 559830
rect 241348 551698 241376 560102
rect 242222 559858 242250 560116
rect 243234 559858 243262 560116
rect 244246 559858 244274 560116
rect 245258 559858 245286 560116
rect 246270 559858 246298 560116
rect 247296 560102 247448 560130
rect 242222 559830 242296 559858
rect 243234 559830 243308 559858
rect 244246 559830 244320 559858
rect 245258 559830 245332 559858
rect 246270 559830 246344 559858
rect 241348 551670 241560 551698
rect 241426 551576 241482 551585
rect 241532 551562 241560 551670
rect 241610 551576 241666 551585
rect 241532 551534 241610 551562
rect 241426 551511 241482 551520
rect 241610 551511 241666 551520
rect 241440 550730 241468 551511
rect 241428 550724 241480 550730
rect 241428 550666 241480 550672
rect 240782 539064 240838 539073
rect 240782 538999 240838 539008
rect 240230 538928 240286 538937
rect 240230 538863 240286 538872
rect 239494 536344 239550 536353
rect 239494 536279 239550 536288
rect 238758 521384 238814 521393
rect 238758 521319 238814 521328
rect 238772 520849 238800 521319
rect 238758 520840 238814 520849
rect 238758 520775 238814 520784
rect 239508 518106 239536 536279
rect 240796 521529 240824 538999
rect 242268 529689 242296 559830
rect 243280 535401 243308 559830
rect 243266 535392 243322 535401
rect 243266 535327 243322 535336
rect 243542 534440 243598 534449
rect 243542 534375 243598 534384
rect 243556 534342 243584 534375
rect 243544 534336 243596 534342
rect 243544 534278 243596 534284
rect 242254 529680 242310 529689
rect 242254 529615 242310 529624
rect 244292 525337 244320 559830
rect 245304 533769 245332 559830
rect 244370 533760 244426 533769
rect 244370 533695 244426 533704
rect 245290 533760 245346 533769
rect 245290 533695 245346 533704
rect 244384 532846 244412 533695
rect 244372 532840 244424 532846
rect 244372 532782 244424 532788
rect 246316 526969 246344 559830
rect 247316 553512 247368 553518
rect 247316 553454 247368 553460
rect 246394 547224 246450 547233
rect 246394 547159 246450 547168
rect 246302 526960 246358 526969
rect 246302 526895 246358 526904
rect 244278 525328 244334 525337
rect 244278 525263 244334 525272
rect 241058 523968 241114 523977
rect 241058 523903 241114 523912
rect 240782 521520 240838 521529
rect 240782 521455 240838 521464
rect 241072 518106 241100 523903
rect 246408 521529 246436 547159
rect 242530 521520 242586 521529
rect 242530 521455 242586 521464
rect 246394 521520 246450 521529
rect 246394 521455 246450 521464
rect 233160 518078 233204 518106
rect 234724 518078 234768 518106
rect 220664 517956 220692 518078
rect 222228 517956 222256 518078
rect 223792 517956 223820 518078
rect 225356 517956 225384 518078
rect 226920 517956 226948 518078
rect 228484 517956 228512 518078
rect 230048 517956 230076 518078
rect 231612 517956 231640 518078
rect 233176 517956 233204 518078
rect 234740 517956 234768 518078
rect 236304 518078 236408 518106
rect 237868 518078 237972 518106
rect 239432 518078 239536 518106
rect 240996 518078 241100 518106
rect 242544 518106 242572 521455
rect 245658 521248 245714 521257
rect 245658 521183 245714 521192
rect 244094 520840 244150 520849
rect 244094 520775 244150 520784
rect 244108 518106 244136 520775
rect 245672 518106 245700 521183
rect 247328 518106 247356 553454
rect 247420 547233 247448 560102
rect 248294 559858 248322 560116
rect 249306 559858 249334 560116
rect 250318 559858 250346 560116
rect 251330 559858 251358 560116
rect 252356 560102 252508 560130
rect 248294 559830 248368 559858
rect 249306 559830 249380 559858
rect 250318 559830 250392 559858
rect 251330 559830 251404 559858
rect 247406 547224 247462 547233
rect 247406 547159 247462 547168
rect 248340 532273 248368 559830
rect 248878 547496 248934 547505
rect 248878 547431 248934 547440
rect 248326 532264 248382 532273
rect 248326 532199 248382 532208
rect 248892 518106 248920 547431
rect 249352 544649 249380 559830
rect 249338 544640 249394 544649
rect 249338 544575 249394 544584
rect 250364 530369 250392 559830
rect 250442 557152 250498 557161
rect 250442 557087 250498 557096
rect 250350 530360 250406 530369
rect 250350 530295 250406 530304
rect 250456 518106 250484 557087
rect 251376 537985 251404 559830
rect 252480 554169 252508 560102
rect 253202 560008 253258 560017
rect 253202 559943 253258 559952
rect 252466 554160 252522 554169
rect 252466 554095 252522 554104
rect 252006 552664 252062 552673
rect 252006 552599 252062 552608
rect 251362 537976 251418 537985
rect 251362 537911 251418 537920
rect 251086 531312 251142 531321
rect 251086 531247 251142 531256
rect 251100 529990 251128 531247
rect 251088 529984 251140 529990
rect 251088 529926 251140 529932
rect 252020 518106 252048 552599
rect 252468 537872 252520 537878
rect 252468 537814 252520 537820
rect 252480 537033 252508 537814
rect 252466 537024 252522 537033
rect 252466 536959 252522 536968
rect 253216 520849 253244 559943
rect 253354 559858 253382 560116
rect 253354 559830 253428 559858
rect 253296 557660 253348 557666
rect 253296 557602 253348 557608
rect 253308 521286 253336 557602
rect 253400 536353 253428 559830
rect 254584 558952 254636 558958
rect 254584 558894 254636 558900
rect 253570 541512 253626 541521
rect 253570 541447 253626 541456
rect 253386 536344 253442 536353
rect 253386 536279 253442 536288
rect 253296 521280 253348 521286
rect 253296 521222 253348 521228
rect 253202 520840 253258 520849
rect 253202 520775 253258 520784
rect 253584 518106 253612 541447
rect 254596 521218 254624 558894
rect 255134 533216 255190 533225
rect 255134 533151 255190 533160
rect 254584 521212 254636 521218
rect 254584 521154 254636 521160
rect 255148 518106 255176 533151
rect 255412 526516 255464 526522
rect 255412 526458 255464 526464
rect 255320 525088 255372 525094
rect 255320 525030 255372 525036
rect 255332 521014 255360 525030
rect 255424 521082 255452 526458
rect 255976 521257 256004 635151
rect 256160 521393 256188 635831
rect 257986 594824 258042 594833
rect 257986 594759 258042 594768
rect 257894 574152 257950 574161
rect 257894 574087 257950 574096
rect 257908 539073 257936 574087
rect 257894 539064 257950 539073
rect 257894 538999 257950 539008
rect 256698 538520 256754 538529
rect 256698 538455 256754 538464
rect 256712 538354 256740 538455
rect 256700 538348 256752 538354
rect 256700 538290 256752 538296
rect 258000 523977 258028 594759
rect 258722 559872 258778 559881
rect 258722 559807 258778 559816
rect 258264 553444 258316 553450
rect 258264 553386 258316 553392
rect 257986 523968 258042 523977
rect 257986 523903 258042 523912
rect 256146 521384 256202 521393
rect 256146 521319 256202 521328
rect 256608 521280 256660 521286
rect 255962 521248 256018 521257
rect 256608 521222 256660 521228
rect 255962 521183 256018 521192
rect 255412 521076 255464 521082
rect 255412 521018 255464 521024
rect 255320 521008 255372 521014
rect 255320 520950 255372 520956
rect 242544 518078 242588 518106
rect 244108 518078 244152 518106
rect 245672 518078 245716 518106
rect 236304 517956 236332 518078
rect 237868 517956 237896 518078
rect 239432 517956 239460 518078
rect 240996 517956 241024 518078
rect 242560 517956 242588 518078
rect 244124 517956 244152 518078
rect 245688 517956 245716 518078
rect 247252 518078 247356 518106
rect 248816 518078 248920 518106
rect 250380 518078 250484 518106
rect 251944 518078 252048 518106
rect 253508 518078 253612 518106
rect 255072 518078 255176 518106
rect 256620 518106 256648 521222
rect 258276 518106 258304 553386
rect 258736 521665 258764 559807
rect 259828 557592 259880 557598
rect 259828 557534 259880 557540
rect 258446 521656 258502 521665
rect 258446 521591 258502 521600
rect 258722 521656 258778 521665
rect 258722 521591 258778 521600
rect 258460 520334 258488 521591
rect 258448 520328 258500 520334
rect 258448 520270 258500 520276
rect 259840 518106 259868 557534
rect 260794 549296 260846 549302
rect 260932 549296 260984 549302
rect 260846 549244 260932 549250
rect 260794 549238 260984 549244
rect 260806 549222 260972 549238
rect 260840 549160 260892 549166
rect 262876 549137 262904 636239
rect 264244 635520 264296 635526
rect 264244 635462 264296 635468
rect 262956 554804 263008 554810
rect 262956 554746 263008 554752
rect 261390 549128 261446 549137
rect 260892 549108 260972 549114
rect 260840 549102 260972 549108
rect 260852 549086 260972 549102
rect 260944 549030 260972 549086
rect 261390 549063 261446 549072
rect 262862 549128 262918 549137
rect 262862 549063 262918 549072
rect 260932 549024 260984 549030
rect 260932 548966 260984 548972
rect 261404 518106 261432 549063
rect 262968 518106 262996 554746
rect 264256 521014 264284 635462
rect 265624 634840 265676 634846
rect 265624 634782 265676 634788
rect 265636 556918 265664 634782
rect 268396 559638 268424 636822
rect 271236 636812 271288 636818
rect 271236 636754 271288 636760
rect 271144 635588 271196 635594
rect 271144 635530 271196 635536
rect 268384 559632 268436 559638
rect 268384 559574 268436 559580
rect 265624 556912 265676 556918
rect 265624 556854 265676 556860
rect 270774 551848 270830 551857
rect 270774 551783 270830 551792
rect 269118 551168 269174 551177
rect 269118 551103 269174 551112
rect 269132 550798 269160 551103
rect 269120 550792 269172 550798
rect 269120 550734 269172 550740
rect 269762 543688 269818 543697
rect 269762 543623 269818 543632
rect 264334 539472 264390 539481
rect 264334 539407 264390 539416
rect 264348 538214 264376 539407
rect 264348 538186 264652 538214
rect 264624 521529 264652 538186
rect 267646 531856 267702 531865
rect 267646 531791 267702 531800
rect 265990 521656 266046 521665
rect 265990 521591 266046 521600
rect 264426 521520 264482 521529
rect 264426 521455 264482 521464
rect 264610 521520 264666 521529
rect 264610 521455 264666 521464
rect 264244 521008 264296 521014
rect 264244 520950 264296 520956
rect 256620 518078 256664 518106
rect 247252 517956 247280 518078
rect 248816 517956 248844 518078
rect 250380 517956 250408 518078
rect 251944 517956 251972 518078
rect 253508 517956 253536 518078
rect 255072 517956 255100 518078
rect 256636 517956 256664 518078
rect 258200 518078 258304 518106
rect 259764 518078 259868 518106
rect 261328 518078 261432 518106
rect 262892 518078 262996 518106
rect 264440 518106 264468 521455
rect 266004 518106 266032 521591
rect 267660 518106 267688 531791
rect 269210 520840 269266 520849
rect 269210 520775 269266 520784
rect 269026 518800 269082 518809
rect 269026 518735 269028 518744
rect 269080 518735 269082 518744
rect 269028 518706 269080 518712
rect 269224 518106 269252 520775
rect 269776 520713 269804 543623
rect 269762 520704 269818 520713
rect 269762 520639 269818 520648
rect 270408 519920 270460 519926
rect 270408 519862 270460 519868
rect 270420 519353 270448 519862
rect 270406 519344 270462 519353
rect 270406 519279 270462 519288
rect 270788 518106 270816 551783
rect 271156 519994 271184 635530
rect 271248 558278 271276 636754
rect 273904 635452 273956 635458
rect 273904 635394 273956 635400
rect 271236 558272 271288 558278
rect 271236 558214 271288 558220
rect 273916 550118 273944 635394
rect 273904 550112 273956 550118
rect 273904 550054 273956 550060
rect 273902 544776 273958 544785
rect 273902 544711 273958 544720
rect 272524 540728 272576 540734
rect 272524 540670 272576 540676
rect 272536 539617 272564 540670
rect 272522 539608 272578 539617
rect 272522 539543 272578 539552
rect 272338 539200 272394 539209
rect 272338 539135 272394 539144
rect 271144 519988 271196 519994
rect 271144 519930 271196 519936
rect 272352 518106 272380 539135
rect 273916 518106 273944 544711
rect 274008 519858 274036 636890
rect 274088 635452 274140 635458
rect 274088 635394 274140 635400
rect 274100 525502 274128 635394
rect 274180 634500 274232 634506
rect 274180 634442 274232 634448
rect 274088 525496 274140 525502
rect 274088 525438 274140 525444
rect 274192 525434 274220 634442
rect 275296 528554 275324 647663
rect 278318 645416 278374 645425
rect 278318 645351 278374 645360
rect 275466 645280 275522 645289
rect 275466 645215 275522 645224
rect 275376 636812 275428 636818
rect 275376 636754 275428 636760
rect 275204 528526 275324 528554
rect 274180 525428 274232 525434
rect 274180 525370 274232 525376
rect 274640 524000 274692 524006
rect 274640 523942 274692 523948
rect 274652 523161 274680 523942
rect 275204 523569 275232 528526
rect 275190 523560 275246 523569
rect 275190 523495 275246 523504
rect 274638 523152 274694 523161
rect 274638 523087 274694 523096
rect 275388 520062 275416 636754
rect 275480 553625 275508 645215
rect 276662 644056 276718 644065
rect 276662 643991 276718 644000
rect 275926 555248 275982 555257
rect 275926 555183 275982 555192
rect 275940 554810 275968 555183
rect 275928 554804 275980 554810
rect 275928 554746 275980 554752
rect 275466 553616 275522 553625
rect 275466 553551 275522 553560
rect 275558 550488 275614 550497
rect 275558 550423 275614 550432
rect 275466 538112 275522 538121
rect 275466 538047 275522 538056
rect 275376 520056 275428 520062
rect 275376 519998 275428 520004
rect 273996 519852 274048 519858
rect 273996 519794 274048 519800
rect 275480 518106 275508 538047
rect 275572 520849 275600 550423
rect 276676 539209 276704 643991
rect 278226 642560 278282 642569
rect 278226 642495 278282 642504
rect 276754 641200 276810 641209
rect 276754 641135 276810 641144
rect 276768 544785 276796 641135
rect 278136 638308 278188 638314
rect 278136 638250 278188 638256
rect 278042 638072 278098 638081
rect 278042 638007 278098 638016
rect 276848 635520 276900 635526
rect 276848 635462 276900 635468
rect 276754 544776 276810 544785
rect 276754 544711 276810 544720
rect 276860 540802 276888 635462
rect 277306 571296 277362 571305
rect 277306 571231 277362 571240
rect 277320 560425 277348 571231
rect 277306 560416 277362 560425
rect 277306 560351 277362 560360
rect 276848 540796 276900 540802
rect 276848 540738 276900 540744
rect 276662 539200 276718 539209
rect 276662 539135 276718 539144
rect 278056 521529 278084 638007
rect 278148 531078 278176 638250
rect 278240 548457 278268 642495
rect 278332 552265 278360 645351
rect 279514 642424 279570 642433
rect 279514 642359 279570 642368
rect 279422 638208 279478 638217
rect 279422 638143 279478 638152
rect 278686 552528 278742 552537
rect 278686 552463 278742 552472
rect 278318 552256 278374 552265
rect 278700 552226 278728 552463
rect 278318 552191 278374 552200
rect 278688 552220 278740 552226
rect 278688 552162 278740 552168
rect 278686 549128 278742 549137
rect 278686 549063 278742 549072
rect 278226 548448 278282 548457
rect 278226 548383 278282 548392
rect 278700 547942 278728 549063
rect 278688 547936 278740 547942
rect 278688 547878 278740 547884
rect 278136 531072 278188 531078
rect 278136 531014 278188 531020
rect 279436 527513 279464 638143
rect 279528 535265 279556 642359
rect 279606 638344 279662 638353
rect 279606 638279 279662 638288
rect 279620 548321 279648 638279
rect 279700 636880 279752 636886
rect 279700 636822 279752 636828
rect 279712 549030 279740 636822
rect 279790 633992 279846 634001
rect 279790 633927 279846 633936
rect 279804 558482 279832 633927
rect 279882 582176 279938 582185
rect 279882 582111 279938 582120
rect 279792 558476 279844 558482
rect 279792 558418 279844 558424
rect 279896 550633 279924 582111
rect 280158 558104 280214 558113
rect 280158 558039 280214 558048
rect 280172 557666 280200 558039
rect 280160 557660 280212 557666
rect 280160 557602 280212 557608
rect 279882 550624 279938 550633
rect 279882 550559 279938 550568
rect 280068 549160 280120 549166
rect 280068 549102 280120 549108
rect 279700 549024 279752 549030
rect 279700 548966 279752 548972
rect 279606 548312 279662 548321
rect 279606 548247 279662 548256
rect 280080 547913 280108 549102
rect 280066 547904 280122 547913
rect 280066 547839 280122 547848
rect 280816 537305 280844 648071
rect 286322 648000 286378 648009
rect 286322 647935 286378 647944
rect 282182 645144 282238 645153
rect 282182 645079 282238 645088
rect 280896 638172 280948 638178
rect 280896 638114 280948 638120
rect 280802 537296 280858 537305
rect 280802 537231 280858 537240
rect 279514 535256 279570 535265
rect 279514 535191 279570 535200
rect 280908 533934 280936 638114
rect 281446 615904 281502 615913
rect 281446 615839 281502 615848
rect 281460 558113 281488 615839
rect 281446 558104 281502 558113
rect 281446 558039 281502 558048
rect 282196 553761 282224 645079
rect 283748 638444 283800 638450
rect 283748 638386 283800 638392
rect 283564 638104 283616 638110
rect 283564 638046 283616 638052
rect 282550 581088 282606 581097
rect 282550 581023 282606 581032
rect 282458 580000 282514 580009
rect 282458 579935 282514 579944
rect 282274 578912 282330 578921
rect 282274 578847 282330 578856
rect 282182 553752 282238 553761
rect 282182 553687 282238 553696
rect 282288 549273 282316 578847
rect 282366 576736 282422 576745
rect 282366 576671 282422 576680
rect 282274 549264 282330 549273
rect 282274 549199 282330 549208
rect 282380 546825 282408 576671
rect 282472 553081 282500 579935
rect 282564 555801 282592 581023
rect 282734 577824 282790 577833
rect 282734 577759 282790 577768
rect 282642 575648 282698 575657
rect 282642 575583 282698 575592
rect 282550 555792 282606 555801
rect 282550 555727 282606 555736
rect 282458 553072 282514 553081
rect 282458 553007 282514 553016
rect 282656 551993 282684 575583
rect 282748 554441 282776 577759
rect 282734 554432 282790 554441
rect 282734 554367 282790 554376
rect 282642 551984 282698 551993
rect 282642 551919 282698 551928
rect 282366 546816 282422 546825
rect 282366 546751 282422 546760
rect 280896 533928 280948 533934
rect 280896 533870 280948 533876
rect 280066 530496 280122 530505
rect 280066 530431 280122 530440
rect 279976 528352 280028 528358
rect 279976 528294 280028 528300
rect 279422 527504 279478 527513
rect 279422 527439 279478 527448
rect 279988 527241 280016 528294
rect 279974 527232 280030 527241
rect 279974 527167 280030 527176
rect 278042 521520 278098 521529
rect 278042 521455 278098 521464
rect 276940 521212 276992 521218
rect 276940 521154 276992 521160
rect 275558 520840 275614 520849
rect 275558 520775 275614 520784
rect 264440 518078 264484 518106
rect 266004 518078 266048 518106
rect 258200 517956 258228 518078
rect 259764 517956 259792 518078
rect 261328 517956 261356 518078
rect 262892 517956 262920 518078
rect 264456 517956 264484 518078
rect 266020 517956 266048 518078
rect 267584 518078 267688 518106
rect 269148 518078 269252 518106
rect 270712 518078 270816 518106
rect 272276 518078 272380 518106
rect 273840 518078 273944 518106
rect 275404 518078 275508 518106
rect 276952 518106 276980 521154
rect 278502 520704 278558 520713
rect 278502 520639 278558 520648
rect 278516 518106 278544 520639
rect 280080 518106 280108 530431
rect 283194 521656 283250 521665
rect 283194 521591 283250 521600
rect 281540 521144 281592 521150
rect 281540 521086 281592 521092
rect 281552 518894 281580 521086
rect 282920 520124 282972 520130
rect 282920 520066 282972 520072
rect 282932 519217 282960 520066
rect 282918 519208 282974 519217
rect 282918 519143 282974 519152
rect 281552 518866 281672 518894
rect 281644 518106 281672 518866
rect 283208 518106 283236 521591
rect 283576 520062 283604 638046
rect 283656 614168 283708 614174
rect 283656 614110 283708 614116
rect 283668 526930 283696 614110
rect 283760 550050 283788 638386
rect 284944 634568 284996 634574
rect 284944 634510 284996 634516
rect 283840 610020 283892 610026
rect 283840 609962 283892 609968
rect 283852 550322 283880 609962
rect 284206 558920 284262 558929
rect 284206 558855 284262 558864
rect 284220 557598 284248 558855
rect 284208 557592 284260 557598
rect 284208 557534 284260 557540
rect 283840 550316 283892 550322
rect 283840 550258 283892 550264
rect 283748 550044 283800 550050
rect 283748 549986 283800 549992
rect 284956 546174 284984 634510
rect 285312 594856 285364 594862
rect 285312 594798 285364 594804
rect 285218 594144 285274 594153
rect 285218 594079 285274 594088
rect 285126 593056 285182 593065
rect 285126 592991 285182 593000
rect 285036 567248 285088 567254
rect 285036 567190 285088 567196
rect 284944 546168 284996 546174
rect 284944 546110 284996 546116
rect 283748 543176 283800 543182
rect 283748 543118 283800 543124
rect 283656 526924 283708 526930
rect 283656 526866 283708 526872
rect 283760 526522 283788 543118
rect 284850 542328 284906 542337
rect 284850 542263 284906 542272
rect 283748 526516 283800 526522
rect 283748 526458 283800 526464
rect 283564 520056 283616 520062
rect 283564 519998 283616 520004
rect 284864 518106 284892 542263
rect 285048 532506 285076 567190
rect 285140 558793 285168 592991
rect 285232 559473 285260 594079
rect 285324 560590 285352 594798
rect 285402 591968 285458 591977
rect 285402 591903 285458 591912
rect 285312 560584 285364 560590
rect 285312 560526 285364 560532
rect 285416 560153 285444 591903
rect 285494 589792 285550 589801
rect 285494 589727 285550 589736
rect 285402 560144 285458 560153
rect 285402 560079 285458 560088
rect 285218 559464 285274 559473
rect 285218 559399 285274 559408
rect 285126 558784 285182 558793
rect 285126 558719 285182 558728
rect 285508 558657 285536 589727
rect 285586 574560 285642 574569
rect 285586 574495 285642 574504
rect 285494 558648 285550 558657
rect 285494 558583 285550 558592
rect 285600 549817 285628 574495
rect 286336 551857 286364 647935
rect 289266 647864 289322 647873
rect 289266 647799 289322 647808
rect 287794 643920 287850 643929
rect 287794 643855 287850 643864
rect 287702 639704 287758 639713
rect 287702 639639 287758 639648
rect 286416 634636 286468 634642
rect 286416 634578 286468 634584
rect 286428 553314 286456 634578
rect 286966 583808 287022 583817
rect 286966 583743 287022 583752
rect 286416 553308 286468 553314
rect 286416 553250 286468 553256
rect 286322 551848 286378 551857
rect 286322 551783 286378 551792
rect 285586 549808 285642 549817
rect 285586 549743 285642 549752
rect 286414 532536 286470 532545
rect 285036 532500 285088 532506
rect 286414 532471 286470 532480
rect 285036 532442 285088 532448
rect 286322 527640 286378 527649
rect 286322 527575 286378 527584
rect 286336 527270 286364 527575
rect 286324 527264 286376 527270
rect 286324 527206 286376 527212
rect 286428 518106 286456 532471
rect 286980 528554 287008 583743
rect 286888 528526 287008 528554
rect 286888 527105 286916 528526
rect 286874 527096 286930 527105
rect 286874 527031 286930 527040
rect 287716 521121 287744 639639
rect 287808 541521 287836 643855
rect 289084 638376 289136 638382
rect 289084 638318 289136 638324
rect 288164 590708 288216 590714
rect 288164 590650 288216 590656
rect 287978 588704 288034 588713
rect 287978 588639 288034 588648
rect 287886 586392 287942 586401
rect 287886 586327 287942 586336
rect 287900 554577 287928 586327
rect 287992 556617 288020 588639
rect 288070 587616 288126 587625
rect 288070 587551 288126 587560
rect 287978 556608 288034 556617
rect 287978 556543 288034 556552
rect 288084 556073 288112 587551
rect 288176 560658 288204 590650
rect 288254 585440 288310 585449
rect 288254 585375 288310 585384
rect 288164 560652 288216 560658
rect 288164 560594 288216 560600
rect 288268 559201 288296 585375
rect 288346 573472 288402 573481
rect 288346 573407 288402 573416
rect 288254 559192 288310 559201
rect 288254 559127 288310 559136
rect 288070 556064 288126 556073
rect 288070 555999 288126 556008
rect 287886 554568 287942 554577
rect 287886 554503 287942 554512
rect 288360 552809 288388 573407
rect 288346 552800 288402 552809
rect 288346 552735 288402 552744
rect 287978 543416 288034 543425
rect 287978 543351 288034 543360
rect 287794 541512 287850 541521
rect 287794 541447 287850 541456
rect 287702 521112 287758 521121
rect 287702 521047 287758 521056
rect 287992 518106 288020 543351
rect 289096 521082 289124 638318
rect 289176 635180 289228 635186
rect 289176 635122 289228 635128
rect 289084 521076 289136 521082
rect 289084 521018 289136 521024
rect 289188 520198 289216 635122
rect 289280 544105 289308 647799
rect 298006 644600 298062 644609
rect 298006 644535 298062 644544
rect 291842 643784 291898 643793
rect 291842 643719 291898 643728
rect 290464 635384 290516 635390
rect 290464 635326 290516 635332
rect 289360 611380 289412 611386
rect 289360 611322 289412 611328
rect 289372 558754 289400 611322
rect 289360 558748 289412 558754
rect 289360 558690 289412 558696
rect 289266 544096 289322 544105
rect 289266 544031 289322 544040
rect 290476 532234 290504 635326
rect 290554 584352 290610 584361
rect 290554 584287 290610 584296
rect 290568 557705 290596 584287
rect 290646 583264 290702 583273
rect 290646 583199 290702 583208
rect 290554 557696 290610 557705
rect 290554 557631 290610 557640
rect 290660 557433 290688 583199
rect 291014 578232 291070 578241
rect 291014 578167 291070 578176
rect 290738 572384 290794 572393
rect 290738 572319 290794 572328
rect 290646 557424 290702 557433
rect 290646 557359 290702 557368
rect 290752 555937 290780 572319
rect 290738 555928 290794 555937
rect 290738 555863 290794 555872
rect 290464 532228 290516 532234
rect 290464 532170 290516 532176
rect 289726 530496 289782 530505
rect 289726 530431 289782 530440
rect 289740 530058 289768 530431
rect 289728 530052 289780 530058
rect 289728 529994 289780 530000
rect 289726 529408 289782 529417
rect 289726 529343 289782 529352
rect 289740 528698 289768 529343
rect 289728 528692 289780 528698
rect 289728 528634 289780 528640
rect 291028 528554 291056 578167
rect 291750 553208 291806 553217
rect 291750 553143 291806 553152
rect 291764 552294 291792 553143
rect 291752 552288 291804 552294
rect 291752 552230 291804 552236
rect 291856 538214 291884 643719
rect 297454 643512 297510 643521
rect 297454 643447 297510 643456
rect 297362 641064 297418 641073
rect 297362 640999 297418 641008
rect 295984 638036 296036 638042
rect 295984 637978 296036 637984
rect 294602 637936 294658 637945
rect 294602 637871 294658 637880
rect 291934 635624 291990 635633
rect 291934 635559 291990 635568
rect 291948 600681 291976 635559
rect 293866 617808 293922 617817
rect 293866 617743 293922 617752
rect 293774 612776 293830 612785
rect 293774 612711 293830 612720
rect 291934 600672 291990 600681
rect 291934 600607 291990 600616
rect 292394 579592 292450 579601
rect 292394 579527 292450 579536
rect 292302 572928 292358 572937
rect 292302 572863 292358 572872
rect 292210 572792 292266 572801
rect 292210 572727 292266 572736
rect 291936 560924 291988 560930
rect 291936 560866 291988 560872
rect 291764 538186 291884 538214
rect 291106 536480 291162 536489
rect 291106 536415 291162 536424
rect 290936 528526 291056 528554
rect 289726 527096 289782 527105
rect 289726 527031 289782 527040
rect 289740 525910 289768 527031
rect 289728 525904 289780 525910
rect 289728 525846 289780 525852
rect 289450 520840 289506 520849
rect 289450 520775 289506 520784
rect 289176 520192 289228 520198
rect 289176 520134 289228 520140
rect 276952 518078 276996 518106
rect 278516 518078 278560 518106
rect 280080 518078 280124 518106
rect 281644 518078 281688 518106
rect 283208 518078 283252 518106
rect 267584 517956 267612 518078
rect 269148 517956 269176 518078
rect 270712 517956 270740 518078
rect 272276 517956 272304 518078
rect 273840 517956 273868 518078
rect 275404 517956 275432 518078
rect 276968 517956 276996 518078
rect 278532 517956 278560 518078
rect 280096 517956 280124 518078
rect 281660 517956 281688 518078
rect 283224 517956 283252 518078
rect 284788 518078 284892 518106
rect 286352 518078 286456 518106
rect 287916 518078 288020 518106
rect 289464 518106 289492 520775
rect 290936 520169 290964 528526
rect 291016 520192 291068 520198
rect 290922 520160 290978 520169
rect 291016 520134 291068 520140
rect 290922 520095 290978 520104
rect 291028 519081 291056 520134
rect 291014 519072 291070 519081
rect 291014 519007 291070 519016
rect 291120 518106 291148 536415
rect 291764 535922 291792 538186
rect 291844 537940 291896 537946
rect 291844 537882 291896 537888
rect 291856 536897 291884 537882
rect 291842 536888 291898 536897
rect 291842 536823 291898 536832
rect 291842 535936 291898 535945
rect 291764 535894 291842 535922
rect 291842 535871 291898 535880
rect 291948 519897 291976 560866
rect 292224 558793 292252 572727
rect 292210 558784 292266 558793
rect 292210 558719 292266 558728
rect 292316 540569 292344 572863
rect 292302 540560 292358 540569
rect 292302 540495 292358 540504
rect 292408 538121 292436 579527
rect 292486 578232 292542 578241
rect 292486 578167 292542 578176
rect 292394 538112 292450 538121
rect 292394 538047 292450 538056
rect 292500 523433 292528 578167
rect 293682 574152 293738 574161
rect 293682 574087 293738 574096
rect 293696 542337 293724 574087
rect 293682 542328 293738 542337
rect 293682 542263 293738 542272
rect 292580 536580 292632 536586
rect 292580 536522 292632 536528
rect 292592 535537 292620 536522
rect 293788 536489 293816 612711
rect 293774 536480 293830 536489
rect 293774 536415 293830 536424
rect 292578 535528 292634 535537
rect 292578 535463 292634 535472
rect 292670 529816 292726 529825
rect 292670 529751 292726 529760
rect 292578 523560 292634 523569
rect 292578 523495 292634 523504
rect 292486 523424 292542 523433
rect 292486 523359 292542 523368
rect 292592 523054 292620 523495
rect 292580 523048 292632 523054
rect 292580 522990 292632 522996
rect 291934 519888 291990 519897
rect 291934 519823 291990 519832
rect 291844 518968 291896 518974
rect 291842 518936 291844 518945
rect 291896 518936 291898 518945
rect 291842 518871 291898 518880
rect 292684 518106 292712 529751
rect 293880 523705 293908 617743
rect 293958 554704 294014 554713
rect 293958 554639 294014 554648
rect 293972 553450 294000 554639
rect 293960 553444 294012 553450
rect 293960 553386 294012 553392
rect 293958 544232 294014 544241
rect 293958 544167 294014 544176
rect 293972 543862 294000 544167
rect 293960 543856 294012 543862
rect 293960 543798 294012 543804
rect 293866 523696 293922 523705
rect 293866 523631 293922 523640
rect 293958 522200 294014 522209
rect 293958 522135 294014 522144
rect 293972 521694 294000 522135
rect 293960 521688 294012 521694
rect 294616 521665 294644 637871
rect 295062 636848 295118 636857
rect 295062 636783 295118 636792
rect 294694 635488 294750 635497
rect 294694 635423 294750 635432
rect 294708 597417 294736 635423
rect 294878 635352 294934 635361
rect 294878 635287 294934 635296
rect 294786 634536 294842 634545
rect 294786 634471 294842 634480
rect 294800 598505 294828 634471
rect 294786 598496 294842 598505
rect 294786 598431 294842 598440
rect 294694 597408 294750 597417
rect 294694 597343 294750 597352
rect 294892 596329 294920 635287
rect 294970 633584 295026 633593
rect 294970 633519 295026 633528
rect 294984 599593 295012 633519
rect 295076 601769 295104 636783
rect 295062 601760 295118 601769
rect 295062 601695 295118 601704
rect 294970 599584 295026 599593
rect 294970 599519 295026 599528
rect 295062 597544 295118 597553
rect 295062 597479 295118 597488
rect 294878 596320 294934 596329
rect 294878 596255 294934 596264
rect 295076 550497 295104 597479
rect 295246 592104 295302 592113
rect 295246 592039 295302 592048
rect 295154 571432 295210 571441
rect 295154 571367 295210 571376
rect 295062 550488 295118 550497
rect 295062 550423 295118 550432
rect 295168 522345 295196 571367
rect 295154 522336 295210 522345
rect 295154 522271 295210 522280
rect 295260 522209 295288 592039
rect 295340 552356 295392 552362
rect 295340 552298 295392 552304
rect 295352 552265 295380 552298
rect 295338 552256 295394 552265
rect 295338 552191 295394 552200
rect 295798 533896 295854 533905
rect 295798 533831 295854 533840
rect 295338 531312 295394 531321
rect 295338 531247 295394 531256
rect 295352 530126 295380 531247
rect 295340 530120 295392 530126
rect 295340 530062 295392 530068
rect 295246 522200 295302 522209
rect 295246 522135 295302 522144
rect 293960 521630 294012 521636
rect 294602 521656 294658 521665
rect 294602 521591 294658 521600
rect 294144 520940 294196 520946
rect 294144 520882 294196 520888
rect 289464 518078 289508 518106
rect 284788 517956 284816 518078
rect 286352 517956 286380 518078
rect 287916 517956 287944 518078
rect 289480 517956 289508 518078
rect 291044 518078 291148 518106
rect 292608 518078 292712 518106
rect 294156 518106 294184 520882
rect 295812 518106 295840 533831
rect 295996 521150 296024 637978
rect 296720 635724 296772 635730
rect 296720 635666 296772 635672
rect 296732 628969 296760 635666
rect 297180 634432 297232 634438
rect 297180 634374 297232 634380
rect 296718 628960 296774 628969
rect 296718 628895 296774 628904
rect 297192 626793 297220 634374
rect 297376 627881 297404 640999
rect 297468 633321 297496 643447
rect 297638 642152 297694 642161
rect 297638 642087 297694 642096
rect 297548 635316 297600 635322
rect 297548 635258 297600 635264
rect 297454 633312 297510 633321
rect 297454 633247 297510 633256
rect 297362 627872 297418 627881
rect 297362 627807 297418 627816
rect 297178 626784 297234 626793
rect 297178 626719 297234 626728
rect 297560 625705 297588 635258
rect 297652 632233 297680 642087
rect 297730 639432 297786 639441
rect 297730 639367 297786 639376
rect 297638 632224 297694 632233
rect 297638 632159 297694 632168
rect 297744 631145 297772 639367
rect 297914 634808 297970 634817
rect 297914 634743 297970 634752
rect 297730 631136 297786 631145
rect 297730 631071 297786 631080
rect 297546 625696 297602 625705
rect 297546 625631 297602 625640
rect 297546 624608 297602 624617
rect 297546 624543 297602 624552
rect 297454 620256 297510 620265
rect 297454 620191 297510 620200
rect 297362 618080 297418 618089
rect 297362 618015 297418 618024
rect 296626 590608 296682 590617
rect 296626 590543 296682 590552
rect 296534 585168 296590 585177
rect 296534 585103 296590 585112
rect 296350 575512 296406 575521
rect 296350 575447 296406 575456
rect 296364 555937 296392 575447
rect 296442 568712 296498 568721
rect 296442 568647 296498 568656
rect 296350 555928 296406 555937
rect 296350 555863 296406 555872
rect 296456 535129 296484 568647
rect 296442 535120 296498 535129
rect 296442 535055 296498 535064
rect 296548 533905 296576 585103
rect 296534 533896 296590 533905
rect 296534 533831 296590 533840
rect 296640 530505 296668 590543
rect 296718 568032 296774 568041
rect 296718 567967 296774 567976
rect 296732 567254 296760 567967
rect 296720 567248 296772 567254
rect 296720 567190 296772 567196
rect 296626 530496 296682 530505
rect 296626 530431 296682 530440
rect 297376 524006 297404 618015
rect 297468 554606 297496 620191
rect 297560 558414 297588 624543
rect 297928 622441 297956 634743
rect 298020 630057 298048 644535
rect 298006 630048 298062 630057
rect 298006 629983 298062 629992
rect 297914 622432 297970 622441
rect 297914 622367 297970 622376
rect 297638 619168 297694 619177
rect 297638 619103 297694 619112
rect 297652 560114 297680 619103
rect 298006 614816 298062 614825
rect 298006 614751 298062 614760
rect 298020 614174 298048 614751
rect 298008 614168 298060 614174
rect 298008 614110 298060 614116
rect 298006 612640 298062 612649
rect 298006 612575 298062 612584
rect 298020 611386 298048 612575
rect 298008 611380 298060 611386
rect 298008 611322 298060 611328
rect 298006 610464 298062 610473
rect 298006 610399 298062 610408
rect 298020 610026 298048 610399
rect 298008 610020 298060 610026
rect 298008 609962 298060 609968
rect 297822 608288 297878 608297
rect 297822 608223 297878 608232
rect 297730 606112 297786 606121
rect 297730 606047 297786 606056
rect 297640 560108 297692 560114
rect 297640 560050 297692 560056
rect 297548 558408 297600 558414
rect 297548 558350 297600 558356
rect 297456 554600 297508 554606
rect 297456 554542 297508 554548
rect 297744 553178 297772 606047
rect 297836 560182 297864 608223
rect 298006 595232 298062 595241
rect 298006 595167 298062 595176
rect 298020 594862 298048 595167
rect 298008 594856 298060 594862
rect 298008 594798 298060 594804
rect 298006 590880 298062 590889
rect 298006 590815 298062 590824
rect 298020 590714 298048 590815
rect 298008 590708 298060 590714
rect 298008 590650 298060 590656
rect 297914 569120 297970 569129
rect 297914 569055 297970 569064
rect 297824 560176 297876 560182
rect 297824 560118 297876 560124
rect 297928 557326 297956 569055
rect 298006 561368 298062 561377
rect 298006 561303 298062 561312
rect 298020 560930 298048 561303
rect 298008 560924 298060 560930
rect 298008 560866 298060 560872
rect 298756 558346 298784 657630
rect 300122 657591 300178 657600
rect 309796 650321 309824 657727
rect 364996 657694 365024 703520
rect 397472 700369 397500 703520
rect 413664 700505 413692 703520
rect 413650 700496 413706 700505
rect 413650 700431 413706 700440
rect 397458 700360 397514 700369
rect 365628 700324 365680 700330
rect 397458 700295 397514 700304
rect 365628 700266 365680 700272
rect 365640 695502 365668 700266
rect 365628 695496 365680 695502
rect 365628 695438 365680 695444
rect 371884 695496 371936 695502
rect 371884 695438 371936 695444
rect 366364 680332 366416 680338
rect 366364 680274 366416 680280
rect 366376 663066 366404 680274
rect 371896 664494 371924 695438
rect 371884 664488 371936 664494
rect 371884 664430 371936 664436
rect 377404 664488 377456 664494
rect 377404 664430 377456 664436
rect 366364 663060 366416 663066
rect 366364 663002 366416 663008
rect 364984 657688 365036 657694
rect 364984 657630 365036 657636
rect 309782 650312 309838 650321
rect 309782 650247 309838 650256
rect 312910 650312 312966 650321
rect 312910 650247 312966 650256
rect 312924 645153 312952 650247
rect 340050 650176 340106 650185
rect 340050 650111 340106 650120
rect 333610 646640 333666 646649
rect 333610 646575 333666 646584
rect 332322 646504 332378 646513
rect 332322 646439 332378 646448
rect 312910 645144 312966 645153
rect 312910 645079 312966 645088
rect 331862 645144 331918 645153
rect 331862 645079 331918 645088
rect 324596 644972 324648 644978
rect 324596 644914 324648 644920
rect 303986 643376 304042 643385
rect 303986 643311 304042 643320
rect 302700 636948 302752 636954
rect 302700 636890 302752 636896
rect 302712 634916 302740 636890
rect 304000 634916 304028 643311
rect 309138 642016 309194 642025
rect 309138 641951 309194 641960
rect 305274 640928 305330 640937
rect 305274 640863 305330 640872
rect 305288 634916 305316 640863
rect 306564 639464 306616 639470
rect 306564 639406 306616 639412
rect 306576 634916 306604 639406
rect 309152 634916 309180 641951
rect 315580 640892 315632 640898
rect 315580 640834 315632 640840
rect 310426 640520 310482 640529
rect 310426 640455 310482 640464
rect 310440 634916 310468 640455
rect 314292 636880 314344 636886
rect 314292 636822 314344 636828
rect 311716 636744 311768 636750
rect 311716 636686 311768 636692
rect 311728 634916 311756 636686
rect 314304 634916 314332 636822
rect 315592 634916 315620 640834
rect 320732 640824 320784 640830
rect 320732 640766 320784 640772
rect 318156 639396 318208 639402
rect 318156 639338 318208 639344
rect 318168 634916 318196 639338
rect 319444 639260 319496 639266
rect 319444 639202 319496 639208
rect 319456 634916 319484 639202
rect 320744 634916 320772 640766
rect 322020 639192 322072 639198
rect 322020 639134 322072 639140
rect 322032 634916 322060 639134
rect 323308 636472 323360 636478
rect 323308 636414 323360 636420
rect 323320 634916 323348 636414
rect 324608 634916 324636 644914
rect 328460 642252 328512 642258
rect 328460 642194 328512 642200
rect 327172 636812 327224 636818
rect 327172 636754 327224 636760
rect 325884 635588 325936 635594
rect 325884 635530 325936 635536
rect 325896 634916 325924 635530
rect 327184 634916 327212 636754
rect 328472 634916 328500 642194
rect 329748 640756 329800 640762
rect 329748 640698 329800 640704
rect 329760 634916 329788 640698
rect 331036 637968 331088 637974
rect 331036 637910 331088 637916
rect 331048 634916 331076 637910
rect 331876 636177 331904 645079
rect 331862 636168 331918 636177
rect 331862 636103 331918 636112
rect 332336 634916 332364 646439
rect 333624 634916 333652 646575
rect 336186 646368 336242 646377
rect 336186 646303 336242 646312
rect 334898 646232 334954 646241
rect 334898 646167 334954 646176
rect 334912 634916 334940 646167
rect 335174 636168 335230 636177
rect 335174 636103 335230 636112
rect 312648 634642 313030 634658
rect 312636 634636 313030 634642
rect 312688 634630 313030 634636
rect 312636 634578 312688 634584
rect 307668 634568 307720 634574
rect 335188 634545 335216 636103
rect 336200 634916 336228 646303
rect 338764 636404 338816 636410
rect 338764 636346 338816 636352
rect 337476 635520 337528 635526
rect 337476 635462 337528 635468
rect 337488 634916 337516 635462
rect 338776 634916 338804 636346
rect 340064 634916 340092 650111
rect 368386 650040 368442 650049
rect 368386 649975 368442 649984
rect 360658 648680 360714 648689
rect 360658 648615 360714 648624
rect 361948 648644 362000 648650
rect 358084 647488 358136 647494
rect 358084 647430 358136 647436
rect 345202 646096 345258 646105
rect 345202 646031 345258 646040
rect 354220 646060 354272 646066
rect 342628 642184 342680 642190
rect 342628 642126 342680 642132
rect 341340 635180 341392 635186
rect 341340 635122 341392 635128
rect 341352 634916 341380 635122
rect 342640 634916 342668 642126
rect 343916 638308 343968 638314
rect 343916 638250 343968 638256
rect 343928 634916 343956 638250
rect 345216 634916 345244 646031
rect 354220 646002 354272 646008
rect 351642 645960 351698 645969
rect 351642 645895 351698 645904
rect 349068 642116 349120 642122
rect 349068 642058 349120 642064
rect 346492 638172 346544 638178
rect 346492 638114 346544 638120
rect 346504 634916 346532 638114
rect 347780 638104 347832 638110
rect 347780 638046 347832 638052
rect 347792 634916 347820 638046
rect 349080 634916 349108 642058
rect 350356 637084 350408 637090
rect 350356 637026 350408 637032
rect 350368 634916 350396 637026
rect 351656 634916 351684 645895
rect 352932 644836 352984 644842
rect 352932 644778 352984 644784
rect 352944 634916 352972 644778
rect 354232 634916 354260 646002
rect 355508 644700 355560 644706
rect 355508 644642 355560 644648
rect 355520 634916 355548 644642
rect 356796 643612 356848 643618
rect 356796 643554 356848 643560
rect 356808 634916 356836 643554
rect 358096 634916 358124 647430
rect 359372 647420 359424 647426
rect 359372 647362 359424 647368
rect 358726 639840 358782 639849
rect 358726 639775 358782 639784
rect 358740 636857 358768 639775
rect 358726 636848 358782 636857
rect 358726 636783 358782 636792
rect 359384 634916 359412 647362
rect 360672 634916 360700 648615
rect 361948 648586 362000 648592
rect 361960 634916 361988 648586
rect 364524 643408 364576 643414
rect 364524 643350 364576 643356
rect 363236 640348 363288 640354
rect 363236 640290 363288 640296
rect 363248 634916 363276 640290
rect 364536 634916 364564 643350
rect 365812 643340 365864 643346
rect 365812 643282 365864 643288
rect 365824 634916 365852 643282
rect 367100 643272 367152 643278
rect 367100 643214 367152 643220
rect 367112 634916 367140 643214
rect 368400 634916 368428 649975
rect 375472 644904 375524 644910
rect 375472 644846 375524 644852
rect 369676 641776 369728 641782
rect 369676 641718 369728 641724
rect 369688 636274 369716 641718
rect 370962 636848 371018 636857
rect 370962 636783 371018 636792
rect 369676 636268 369728 636274
rect 369676 636210 369728 636216
rect 369688 634916 369716 636210
rect 370976 634916 371004 636783
rect 374552 636268 374604 636274
rect 374552 636210 374604 636216
rect 372252 635452 372304 635458
rect 372252 635394 372304 635400
rect 372264 634916 372292 635394
rect 335174 634536 335230 634545
rect 307720 634516 307878 634522
rect 307668 634510 307878 634516
rect 307680 634494 307878 634510
rect 316512 634506 316894 634522
rect 316500 634500 316894 634506
rect 316552 634494 316894 634500
rect 335174 634471 335230 634480
rect 316500 634442 316552 634448
rect 374564 632738 374592 636210
rect 374552 632732 374604 632738
rect 374552 632674 374604 632680
rect 375378 619440 375434 619449
rect 375378 619375 375434 619384
rect 374550 616720 374606 616729
rect 374550 616655 374606 616664
rect 299294 608560 299350 608569
rect 299294 608495 299350 608504
rect 299202 591424 299258 591433
rect 299202 591359 299258 591368
rect 299110 570072 299166 570081
rect 299110 570007 299166 570016
rect 298744 558340 298796 558346
rect 298744 558282 298796 558288
rect 297916 557320 297968 557326
rect 297916 557262 297968 557268
rect 297732 553172 297784 553178
rect 297732 553114 297784 553120
rect 299124 546417 299152 570007
rect 299216 554577 299244 591359
rect 299202 554568 299258 554577
rect 299202 554503 299258 554512
rect 299308 554418 299336 608495
rect 299386 604480 299442 604489
rect 299386 604415 299442 604424
rect 299216 554390 299336 554418
rect 299216 553194 299244 554390
rect 299294 553888 299350 553897
rect 299294 553823 299350 553832
rect 299308 553518 299336 553823
rect 299296 553512 299348 553518
rect 299296 553454 299348 553460
rect 299294 553344 299350 553353
rect 299294 553279 299296 553288
rect 299348 553279 299350 553288
rect 299296 553250 299348 553256
rect 299294 553208 299350 553217
rect 299216 553166 299294 553194
rect 299294 553143 299350 553152
rect 298926 546408 298982 546417
rect 298926 546343 298982 546352
rect 299110 546408 299166 546417
rect 299110 546343 299166 546352
rect 298744 539368 298796 539374
rect 298744 539310 298796 539316
rect 298756 525094 298784 539310
rect 298744 525088 298796 525094
rect 298744 525030 298796 525036
rect 297364 524000 297416 524006
rect 297364 523942 297416 523948
rect 297362 522608 297418 522617
rect 297362 522543 297418 522552
rect 295984 521144 296036 521150
rect 295984 521086 296036 521092
rect 297376 518106 297404 522543
rect 298940 518106 298968 546343
rect 299400 528554 299428 604415
rect 299846 570072 299902 570081
rect 299846 570007 299902 570016
rect 299754 561640 299810 561649
rect 299754 561575 299810 561584
rect 299768 560318 299796 561575
rect 299756 560312 299808 560318
rect 299756 560254 299808 560260
rect 299308 528526 299428 528554
rect 299308 523569 299336 528526
rect 299388 525496 299440 525502
rect 299388 525438 299440 525444
rect 299400 524521 299428 525438
rect 299386 524512 299442 524521
rect 299386 524447 299442 524456
rect 299388 523796 299440 523802
rect 299388 523738 299440 523744
rect 299294 523560 299350 523569
rect 299294 523495 299350 523504
rect 299400 523433 299428 523738
rect 299386 523424 299442 523433
rect 299386 523359 299442 523368
rect 299860 520985 299888 570007
rect 309784 560312 309836 560318
rect 309784 560254 309836 560260
rect 300490 540832 300546 540841
rect 300490 540767 300546 540776
rect 299846 520976 299902 520985
rect 299846 520911 299902 520920
rect 300504 518106 300532 540767
rect 300766 526144 300822 526153
rect 300766 526079 300822 526088
rect 300780 525978 300808 526079
rect 300768 525972 300820 525978
rect 300768 525914 300820 525920
rect 301516 521354 301544 560116
rect 302528 544882 302556 560116
rect 303264 560102 303554 560130
rect 303264 551449 303292 560102
rect 303528 553308 303580 553314
rect 303528 553250 303580 553256
rect 303250 551440 303306 551449
rect 303250 551375 303306 551384
rect 302516 544876 302568 544882
rect 302516 544818 302568 544824
rect 302054 542056 302110 542065
rect 302054 541991 302110 542000
rect 301504 521348 301556 521354
rect 301504 521290 301556 521296
rect 302068 518106 302096 541991
rect 294156 518078 294200 518106
rect 291044 517956 291072 518078
rect 292608 517956 292636 518078
rect 294172 517956 294200 518078
rect 295736 518078 295840 518106
rect 297300 518078 297404 518106
rect 298864 518078 298968 518106
rect 300428 518078 300532 518106
rect 301992 518078 302096 518106
rect 303540 518106 303568 553250
rect 304264 552696 304316 552702
rect 304264 552638 304316 552644
rect 304276 539374 304304 552638
rect 304552 540433 304580 560116
rect 305564 553246 305592 560116
rect 305552 553240 305604 553246
rect 305552 553182 305604 553188
rect 306576 547670 306604 560116
rect 306564 547664 306616 547670
rect 306564 547606 306616 547612
rect 305184 546576 305236 546582
rect 305184 546518 305236 546524
rect 304538 540424 304594 540433
rect 304538 540359 304594 540368
rect 304264 539368 304316 539374
rect 304264 539310 304316 539316
rect 305196 518106 305224 546518
rect 307588 543590 307616 560116
rect 308310 552392 308366 552401
rect 308310 552327 308366 552336
rect 307576 543584 307628 543590
rect 307576 543526 307628 543532
rect 306746 534984 306802 534993
rect 306746 534919 306802 534928
rect 306760 518106 306788 534919
rect 308324 518106 308352 552327
rect 308600 544950 308628 560116
rect 309612 546009 309640 560116
rect 309598 546000 309654 546009
rect 309598 545935 309654 545944
rect 308588 544944 308640 544950
rect 308588 544886 308640 544892
rect 303540 518078 303584 518106
rect 295736 517956 295764 518078
rect 297300 517956 297328 518078
rect 298864 517956 298892 518078
rect 300428 517956 300456 518078
rect 301992 517956 302020 518078
rect 303556 517956 303584 518078
rect 305120 518078 305224 518106
rect 306684 518078 306788 518106
rect 308248 518078 308352 518106
rect 309796 518106 309824 560254
rect 310624 554674 310652 560116
rect 310612 554668 310664 554674
rect 310612 554610 310664 554616
rect 311438 538656 311494 538665
rect 311438 538591 311494 538600
rect 311452 518106 311480 538591
rect 311636 536586 311664 560116
rect 311624 536580 311676 536586
rect 311624 536522 311676 536528
rect 312648 526998 312676 560116
rect 313660 549166 313688 560116
rect 313648 549160 313700 549166
rect 313648 549102 313700 549108
rect 314672 542230 314700 560116
rect 314660 542224 314712 542230
rect 314660 542166 314712 542172
rect 315684 537878 315712 560116
rect 316696 539442 316724 560116
rect 317708 540734 317736 560116
rect 318720 543658 318748 560116
rect 318708 543652 318760 543658
rect 318708 543594 318760 543600
rect 317696 540728 317748 540734
rect 317696 540670 317748 540676
rect 316684 539436 316736 539442
rect 316684 539378 316736 539384
rect 315672 537872 315724 537878
rect 315672 537814 315724 537820
rect 319732 531049 319760 560116
rect 320744 547738 320772 560116
rect 320824 554056 320876 554062
rect 320824 553998 320876 554004
rect 320732 547732 320784 547738
rect 320732 547674 320784 547680
rect 319718 531040 319774 531049
rect 319718 530975 319774 530984
rect 312636 526992 312688 526998
rect 312636 526934 312688 526940
rect 313004 523048 313056 523054
rect 313004 522990 313056 522996
rect 313016 518106 313044 522990
rect 314474 521656 314530 521665
rect 314474 521591 314530 521600
rect 309796 518078 309840 518106
rect 305120 517956 305148 518078
rect 306684 517956 306712 518078
rect 308248 517956 308276 518078
rect 309812 517956 309840 518078
rect 311376 518078 311480 518106
rect 312940 518078 313044 518106
rect 314488 518106 314516 521591
rect 317602 521520 317658 521529
rect 317602 521455 317658 521464
rect 316038 521112 316094 521121
rect 316038 521047 316094 521056
rect 316052 518106 316080 521047
rect 317616 518106 317644 521455
rect 319166 521384 319222 521393
rect 319166 521319 319222 521328
rect 319180 518106 319208 521319
rect 320836 518106 320864 553998
rect 321756 535362 321784 560116
rect 322768 549098 322796 560116
rect 322756 549092 322808 549098
rect 322756 549034 322808 549040
rect 323780 546242 323808 560116
rect 323768 546236 323820 546242
rect 323768 546178 323820 546184
rect 323950 545048 324006 545057
rect 323950 544983 324006 544992
rect 321744 535356 321796 535362
rect 321744 535298 321796 535304
rect 322294 521248 322350 521257
rect 322294 521183 322350 521192
rect 314488 518078 314532 518106
rect 316052 518078 316096 518106
rect 317616 518078 317660 518106
rect 319180 518078 319224 518106
rect 311376 517956 311404 518078
rect 312940 517956 312968 518078
rect 314504 517956 314532 518078
rect 316068 517956 316096 518078
rect 317632 517956 317660 518078
rect 319196 517956 319224 518078
rect 320760 518078 320864 518106
rect 322308 518106 322336 521183
rect 323964 518106 323992 544983
rect 324792 533497 324820 560116
rect 324778 533488 324834 533497
rect 324778 533423 324834 533432
rect 325514 529000 325570 529009
rect 325514 528935 325570 528944
rect 324318 524376 324374 524385
rect 324318 524311 324374 524320
rect 324332 521121 324360 524311
rect 324318 521112 324374 521121
rect 324318 521047 324374 521056
rect 325528 518106 325556 528935
rect 325804 525570 325832 560116
rect 326816 550390 326844 560116
rect 326804 550384 326856 550390
rect 326804 550326 326856 550332
rect 327828 533798 327856 560116
rect 328840 551818 328868 560116
rect 328828 551812 328880 551818
rect 328828 551754 328880 551760
rect 328644 549976 328696 549982
rect 328644 549918 328696 549924
rect 327816 533792 327868 533798
rect 327816 533734 327868 533740
rect 326986 527640 327042 527649
rect 326986 527575 327042 527584
rect 325792 525564 325844 525570
rect 325792 525506 325844 525512
rect 322308 518078 322352 518106
rect 320760 517956 320788 518078
rect 322324 517956 322352 518078
rect 323888 518078 323992 518106
rect 325452 518078 325556 518106
rect 327000 518106 327028 527575
rect 328656 518106 328684 549918
rect 329852 532574 329880 560116
rect 330864 536654 330892 560116
rect 331876 538014 331904 560116
rect 332600 555620 332652 555626
rect 332600 555562 332652 555568
rect 332612 552702 332640 555562
rect 332600 552696 332652 552702
rect 332600 552638 332652 552644
rect 332888 539510 332916 560116
rect 332876 539504 332928 539510
rect 332876 539446 332928 539452
rect 331864 538008 331916 538014
rect 331864 537950 331916 537956
rect 330852 536648 330904 536654
rect 330852 536590 330904 536596
rect 331770 535936 331826 535945
rect 331770 535871 331826 535880
rect 329840 532568 329892 532574
rect 329840 532510 329892 532516
rect 330208 532228 330260 532234
rect 330208 532170 330260 532176
rect 330220 518106 330248 532170
rect 331784 518106 331812 535871
rect 333334 534576 333390 534585
rect 333334 534511 333390 534520
rect 333348 518106 333376 534511
rect 333900 527066 333928 560116
rect 334912 529553 334940 560116
rect 335924 531146 335952 560116
rect 336936 538801 336964 560116
rect 336922 538792 336978 538801
rect 336922 538727 336978 538736
rect 336462 535256 336518 535265
rect 336462 535191 336518 535200
rect 335912 531140 335964 531146
rect 335912 531082 335964 531088
rect 334898 529544 334954 529553
rect 334898 529479 334954 529488
rect 334898 528456 334954 528465
rect 334898 528391 334954 528400
rect 333888 527060 333940 527066
rect 333888 527002 333940 527008
rect 334912 518106 334940 528391
rect 336476 518106 336504 535191
rect 337948 531010 337976 560116
rect 338026 539200 338082 539209
rect 338026 539135 338082 539144
rect 337936 531004 337988 531010
rect 337936 530946 337988 530952
rect 338040 518106 338068 539135
rect 338960 533866 338988 560116
rect 339972 556102 340000 560116
rect 339960 556096 340012 556102
rect 339960 556038 340012 556044
rect 339590 542872 339646 542881
rect 339590 542807 339646 542816
rect 338948 533860 339000 533866
rect 338948 533802 339000 533808
rect 339604 518106 339632 542807
rect 340984 532642 341012 560116
rect 341154 541512 341210 541521
rect 341154 541447 341210 541456
rect 340972 532636 341024 532642
rect 340972 532578 341024 532584
rect 341168 518106 341196 541447
rect 341996 536722 342024 560116
rect 343008 549234 343036 560116
rect 342996 549228 343048 549234
rect 342996 549170 343048 549176
rect 342718 548312 342774 548321
rect 342718 548247 342774 548256
rect 341984 536716 342036 536722
rect 341984 536658 342036 536664
rect 342732 518106 342760 548247
rect 344020 536790 344048 560116
rect 344282 544096 344338 544105
rect 344282 544031 344338 544040
rect 344008 536784 344060 536790
rect 344008 536726 344060 536732
rect 344296 518106 344324 544031
rect 345032 543726 345060 560116
rect 346044 547806 346072 560116
rect 347056 553382 347084 560116
rect 347044 553376 347096 553382
rect 347044 553318 347096 553324
rect 348068 551954 348096 560116
rect 348056 551948 348108 551954
rect 348056 551890 348108 551896
rect 347410 548448 347466 548457
rect 347410 548383 347466 548392
rect 346032 547800 346084 547806
rect 346032 547742 346084 547748
rect 345846 544776 345902 544785
rect 345846 544711 345902 544720
rect 345020 543720 345072 543726
rect 345020 543662 345072 543668
rect 345860 518106 345888 544711
rect 347424 518106 347452 548383
rect 348976 543856 349028 543862
rect 348976 543798 349028 543804
rect 348988 518106 349016 543798
rect 349080 540870 349108 560116
rect 350092 554742 350120 560116
rect 350080 554736 350132 554742
rect 350080 554678 350132 554684
rect 350446 551848 350502 551857
rect 350446 551783 350502 551792
rect 349068 540864 349120 540870
rect 349068 540806 349120 540812
rect 327000 518078 327044 518106
rect 323888 517956 323916 518078
rect 325452 517956 325480 518078
rect 327016 517956 327044 518078
rect 328580 518078 328684 518106
rect 330144 518078 330248 518106
rect 331708 518078 331812 518106
rect 333272 518078 333376 518106
rect 334836 518078 334940 518106
rect 336400 518078 336504 518106
rect 337964 518078 338068 518106
rect 339528 518078 339632 518106
rect 341092 518078 341196 518106
rect 342656 518078 342760 518106
rect 344220 518078 344324 518106
rect 345784 518078 345888 518106
rect 347348 518078 347452 518106
rect 348912 518078 349016 518106
rect 350460 518106 350488 551783
rect 351104 525706 351132 560116
rect 352024 560102 352130 560130
rect 352024 540938 352052 560102
rect 353128 550526 353156 560116
rect 353666 553616 353722 553625
rect 353666 553551 353722 553560
rect 353116 550520 353168 550526
rect 353116 550462 353168 550468
rect 352104 550112 352156 550118
rect 352104 550054 352156 550060
rect 352012 540932 352064 540938
rect 352012 540874 352064 540880
rect 351092 525700 351144 525706
rect 351092 525642 351144 525648
rect 352116 518106 352144 550054
rect 353680 518106 353708 553551
rect 354140 534002 354168 560116
rect 354128 533996 354180 534002
rect 354128 533938 354180 533944
rect 355152 531214 355180 560116
rect 356164 552022 356192 560116
rect 356152 552016 356204 552022
rect 356152 551958 356204 551964
rect 356796 547324 356848 547330
rect 356796 547266 356848 547272
rect 355232 541884 355284 541890
rect 355232 541826 355284 541832
rect 355140 531208 355192 531214
rect 355140 531150 355192 531156
rect 355244 518106 355272 541826
rect 356808 518106 356836 547266
rect 357176 543182 357204 560116
rect 357164 543176 357216 543182
rect 357164 543118 357216 543124
rect 358188 535430 358216 560116
rect 358360 552356 358412 552362
rect 358360 552298 358412 552304
rect 358176 535424 358228 535430
rect 358176 535366 358228 535372
rect 358372 518106 358400 552298
rect 359200 551342 359228 560116
rect 360212 558210 360240 560116
rect 361224 558822 361252 560116
rect 361212 558816 361264 558822
rect 361212 558758 361264 558764
rect 360200 558204 360252 558210
rect 360200 558146 360252 558152
rect 360844 555552 360896 555558
rect 360844 555494 360896 555500
rect 359188 551336 359240 551342
rect 359188 551278 359240 551284
rect 359922 537296 359978 537305
rect 359922 537231 359978 537240
rect 359936 518106 359964 537231
rect 360856 520946 360884 555494
rect 361486 553752 361542 553761
rect 361486 553687 361542 553696
rect 360844 520940 360896 520946
rect 360844 520882 360896 520888
rect 361500 518106 361528 553687
rect 362236 546310 362264 560116
rect 363052 548684 363104 548690
rect 363052 548626 363104 548632
rect 362224 546304 362276 546310
rect 362224 546246 362276 546252
rect 363064 518106 363092 548626
rect 363248 529854 363276 560116
rect 364260 542366 364288 560116
rect 365272 550594 365300 560116
rect 365260 550588 365312 550594
rect 365260 550530 365312 550536
rect 364616 550044 364668 550050
rect 364616 549986 364668 549992
rect 364248 542360 364300 542366
rect 364248 542302 364300 542308
rect 363236 529848 363288 529854
rect 363236 529790 363288 529796
rect 364628 518106 364656 549986
rect 366284 531282 366312 560116
rect 367296 538082 367324 560116
rect 367284 538076 367336 538082
rect 367284 538018 367336 538024
rect 368308 532710 368336 560116
rect 369216 543108 369268 543114
rect 369216 543050 369268 543056
rect 368296 532704 368348 532710
rect 368296 532646 368348 532652
rect 366272 531276 366324 531282
rect 366272 531218 366324 531224
rect 367006 523832 367062 523841
rect 367006 523767 367062 523776
rect 367020 521257 367048 523767
rect 367006 521248 367062 521257
rect 367006 521183 367062 521192
rect 367560 521144 367612 521150
rect 367560 521086 367612 521092
rect 366088 521076 366140 521082
rect 366088 521018 366140 521024
rect 350460 518078 350504 518106
rect 328580 517956 328608 518078
rect 330144 517956 330172 518078
rect 331708 517956 331736 518078
rect 333272 517956 333300 518078
rect 334836 517956 334864 518078
rect 336400 517956 336428 518078
rect 337964 517956 337992 518078
rect 339528 517956 339556 518078
rect 341092 517956 341120 518078
rect 342656 517956 342684 518078
rect 344220 517956 344248 518078
rect 345784 517956 345812 518078
rect 347348 517956 347376 518078
rect 348912 517956 348940 518078
rect 350476 517956 350504 518078
rect 352040 518078 352144 518106
rect 353604 518078 353708 518106
rect 355168 518078 355272 518106
rect 356732 518078 356836 518106
rect 358296 518078 358400 518106
rect 359860 518078 359964 518106
rect 361424 518078 361528 518106
rect 362988 518078 363092 518106
rect 364552 518078 364656 518106
rect 366100 518106 366128 521018
rect 367572 518894 367600 521086
rect 367572 518866 367692 518894
rect 367664 518106 367692 518866
rect 369228 518106 369256 543050
rect 369320 534070 369348 560116
rect 370332 538150 370360 560116
rect 371344 545018 371372 560116
rect 372068 559904 372120 559910
rect 372068 559846 372120 559852
rect 371884 559836 371936 559842
rect 371884 559778 371936 559784
rect 371332 545012 371384 545018
rect 371332 544954 371384 544960
rect 370320 538144 370372 538150
rect 370320 538086 370372 538092
rect 369308 534064 369360 534070
rect 369308 534006 369360 534012
rect 370780 521008 370832 521014
rect 370780 520950 370832 520956
rect 370792 518106 370820 520950
rect 371896 520130 371924 559778
rect 371976 559768 372028 559774
rect 371976 559710 372028 559716
rect 371988 522714 372016 559710
rect 372080 525502 372108 559846
rect 372160 559700 372212 559706
rect 372160 559642 372212 559648
rect 372172 527134 372200 559642
rect 372250 546680 372306 546689
rect 372250 546615 372306 546624
rect 372160 527128 372212 527134
rect 372160 527070 372212 527076
rect 372068 525496 372120 525502
rect 372068 525438 372120 525444
rect 371976 522708 372028 522714
rect 371976 522650 372028 522656
rect 372264 521393 372292 546615
rect 372356 546446 372384 560116
rect 372620 558204 372672 558210
rect 372620 558146 372672 558152
rect 372632 555626 372660 558146
rect 372620 555620 372672 555626
rect 372620 555562 372672 555568
rect 372344 546440 372396 546446
rect 372344 546382 372396 546388
rect 373368 539578 373396 560116
rect 373356 539572 373408 539578
rect 373356 539514 373408 539520
rect 372436 539028 372488 539034
rect 372436 538970 372488 538976
rect 372250 521384 372306 521393
rect 372250 521319 372306 521328
rect 371884 520124 371936 520130
rect 371884 520066 371936 520072
rect 372448 518106 372476 538970
rect 374564 529650 374592 616655
rect 374734 614816 374790 614825
rect 374734 614751 374790 614760
rect 374642 599176 374698 599185
rect 374642 599111 374698 599120
rect 374552 529644 374604 529650
rect 374552 529586 374604 529592
rect 373908 521008 373960 521014
rect 373908 520950 373960 520956
rect 366100 518078 366144 518106
rect 367664 518078 367708 518106
rect 369228 518078 369272 518106
rect 370792 518078 370836 518106
rect 352040 517956 352068 518078
rect 353604 517956 353632 518078
rect 355168 517956 355196 518078
rect 356732 517956 356760 518078
rect 358296 517956 358324 518078
rect 359860 517956 359888 518078
rect 361424 517956 361452 518078
rect 362988 517956 363016 518078
rect 364552 517956 364580 518078
rect 366116 517956 366144 518078
rect 367680 517956 367708 518078
rect 369244 517956 369272 518078
rect 370808 517956 370836 518078
rect 372372 518078 372476 518106
rect 373920 518106 373948 520950
rect 374656 518226 374684 599111
rect 374748 528494 374776 614751
rect 375392 529786 375420 619375
rect 375484 610473 375512 644846
rect 377416 643754 377444 664430
rect 382280 663060 382332 663066
rect 382280 663002 382332 663008
rect 382292 660346 382320 663002
rect 382280 660340 382332 660346
rect 382280 660282 382332 660288
rect 388444 660340 388496 660346
rect 388444 660282 388496 660288
rect 388456 658238 388484 660282
rect 388444 658232 388496 658238
rect 388444 658174 388496 658180
rect 393964 658232 394016 658238
rect 393964 658174 394016 658180
rect 393976 648582 394004 658174
rect 429856 657762 429884 703520
rect 429844 657756 429896 657762
rect 429844 657698 429896 657704
rect 393964 648576 394016 648582
rect 393964 648518 394016 648524
rect 397368 648576 397420 648582
rect 397368 648518 397420 648524
rect 397380 644706 397408 648518
rect 461674 647592 461730 647601
rect 461674 647527 461730 647536
rect 461582 644872 461638 644881
rect 461582 644807 461638 644816
rect 397368 644700 397420 644706
rect 397368 644642 397420 644648
rect 404360 644700 404412 644706
rect 404360 644642 404412 644648
rect 377404 643748 377456 643754
rect 377404 643690 377456 643696
rect 397460 643748 397512 643754
rect 397460 643690 397512 643696
rect 376758 642696 376814 642705
rect 376758 642631 376814 642640
rect 375564 637628 375616 637634
rect 375564 637570 375616 637576
rect 375470 610464 375526 610473
rect 375470 610399 375526 610408
rect 375576 609657 375604 637570
rect 376022 634536 376078 634545
rect 376022 634471 376078 634480
rect 376036 622985 376064 634471
rect 376022 622976 376078 622985
rect 376022 622911 376078 622920
rect 375654 618624 375710 618633
rect 375654 618559 375710 618568
rect 375562 609648 375618 609657
rect 375562 609583 375618 609592
rect 375470 600672 375526 600681
rect 375470 600607 375526 600616
rect 375380 529780 375432 529786
rect 375380 529722 375432 529728
rect 374736 528488 374788 528494
rect 374736 528430 374788 528436
rect 375484 524278 375512 600607
rect 375562 597408 375618 597417
rect 375562 597343 375618 597352
rect 375472 524272 375524 524278
rect 375472 524214 375524 524220
rect 375576 522850 375604 597343
rect 375668 547874 375696 618559
rect 375930 614544 375986 614553
rect 375930 614479 375986 614488
rect 375838 596592 375894 596601
rect 375838 596527 375894 596536
rect 375746 594144 375802 594153
rect 375746 594079 375802 594088
rect 375656 547868 375708 547874
rect 375656 547810 375708 547816
rect 375760 524210 375788 594079
rect 375852 528358 375880 596527
rect 375944 555490 375972 614479
rect 376772 608025 376800 642631
rect 376942 641336 376998 641345
rect 376942 641271 376998 641280
rect 376852 639124 376904 639130
rect 376852 639066 376904 639072
rect 376758 608016 376814 608025
rect 376758 607951 376814 607960
rect 376864 607209 376892 639066
rect 376956 611289 376984 641271
rect 397472 640286 397500 643690
rect 404372 640354 404400 644642
rect 404360 640348 404412 640354
rect 404360 640290 404412 640296
rect 410524 640348 410576 640354
rect 410524 640290 410576 640296
rect 397460 640280 397512 640286
rect 397460 640222 397512 640228
rect 400864 640280 400916 640286
rect 400864 640222 400916 640228
rect 381544 637696 381596 637702
rect 381544 637638 381596 637644
rect 377036 635656 377088 635662
rect 377036 635598 377088 635604
rect 377048 621897 377076 635598
rect 377220 634976 377272 634982
rect 377220 634918 377272 634924
rect 377128 634908 377180 634914
rect 377128 634850 377180 634856
rect 377140 625161 377168 634850
rect 377126 625152 377182 625161
rect 377126 625087 377182 625096
rect 377232 622713 377260 634918
rect 377678 625968 377734 625977
rect 377678 625903 377734 625912
rect 377692 625598 377720 625903
rect 377680 625592 377732 625598
rect 377680 625534 377732 625540
rect 380992 625592 381044 625598
rect 380992 625534 381044 625540
rect 377678 624336 377734 624345
rect 377678 624271 377734 624280
rect 377692 623830 377720 624271
rect 377680 623824 377732 623830
rect 377680 623766 377732 623772
rect 377770 623520 377826 623529
rect 377770 623455 377826 623464
rect 377218 622704 377274 622713
rect 377218 622639 377274 622648
rect 377784 622470 377812 623455
rect 377772 622464 377824 622470
rect 377772 622406 377824 622412
rect 377034 621888 377090 621897
rect 377034 621823 377090 621832
rect 377034 621072 377090 621081
rect 377034 621007 377036 621016
rect 377088 621007 377090 621016
rect 379520 621036 379572 621042
rect 377036 620978 377088 620984
rect 379520 620978 379572 620984
rect 378046 619712 378102 619721
rect 378102 619670 378272 619698
rect 378046 619647 378102 619656
rect 378046 616176 378102 616185
rect 378046 616111 378102 616120
rect 378060 615494 378088 616111
rect 378060 615466 378180 615494
rect 377126 612096 377182 612105
rect 377126 612031 377182 612040
rect 376942 611280 376998 611289
rect 376942 611215 376998 611224
rect 376850 607200 376906 607209
rect 376850 607135 376906 607144
rect 376758 601488 376814 601497
rect 376758 601423 376814 601432
rect 376114 575376 376170 575385
rect 376114 575311 376170 575320
rect 376022 573744 376078 573753
rect 376022 573679 376078 573688
rect 376036 557394 376064 573679
rect 376128 560250 376156 575311
rect 376116 560244 376168 560250
rect 376116 560186 376168 560192
rect 376024 557388 376076 557394
rect 376024 557330 376076 557336
rect 375932 555484 375984 555490
rect 375932 555426 375984 555432
rect 376772 530777 376800 601423
rect 376850 598224 376906 598233
rect 376850 598159 376906 598168
rect 376758 530768 376814 530777
rect 376758 530703 376814 530712
rect 376864 529281 376892 598159
rect 377034 588432 377090 588441
rect 377034 588367 377090 588376
rect 377048 587926 377076 588367
rect 377036 587920 377088 587926
rect 377036 587862 377088 587868
rect 377034 585984 377090 585993
rect 377034 585919 377090 585928
rect 377048 585206 377076 585919
rect 377036 585200 377088 585206
rect 377036 585142 377088 585148
rect 377034 579456 377090 579465
rect 377034 579391 377090 579400
rect 377048 578270 377076 579391
rect 377036 578264 377088 578270
rect 377036 578206 377088 578212
rect 377034 576192 377090 576201
rect 377034 576127 377090 576136
rect 377048 557462 377076 576127
rect 377140 558210 377168 612031
rect 378046 606384 378102 606393
rect 378046 606319 378102 606328
rect 378060 605878 378088 606319
rect 378048 605872 378100 605878
rect 378048 605814 378100 605820
rect 377954 605568 378010 605577
rect 377954 605503 378010 605512
rect 377968 604518 377996 605503
rect 378046 604752 378102 604761
rect 378046 604687 378102 604696
rect 378060 604586 378088 604687
rect 378048 604580 378100 604586
rect 378048 604522 378100 604528
rect 377956 604512 378008 604518
rect 377956 604454 378008 604460
rect 378046 603936 378102 603945
rect 378046 603871 378102 603880
rect 378060 603294 378088 603871
rect 378048 603288 378100 603294
rect 378048 603230 378100 603236
rect 378048 603152 378100 603158
rect 378046 603120 378048 603129
rect 378100 603120 378102 603129
rect 378046 603055 378102 603064
rect 378046 594960 378102 594969
rect 378046 594895 378102 594904
rect 378060 594862 378088 594895
rect 378048 594856 378100 594862
rect 378048 594798 378100 594804
rect 377954 593328 378010 593337
rect 377954 593263 378010 593272
rect 377968 592074 377996 593263
rect 378046 592512 378102 592521
rect 378046 592447 378102 592456
rect 378060 592142 378088 592447
rect 378048 592136 378100 592142
rect 378048 592078 378100 592084
rect 377956 592068 378008 592074
rect 377956 592010 378008 592016
rect 378046 590880 378102 590889
rect 378046 590815 378102 590824
rect 378060 590714 378088 590815
rect 378048 590708 378100 590714
rect 378048 590650 378100 590656
rect 378046 590064 378102 590073
rect 378046 589999 378102 590008
rect 378060 589694 378088 589999
rect 378048 589688 378100 589694
rect 378048 589630 378100 589636
rect 378046 589248 378102 589257
rect 378046 589183 378102 589192
rect 378060 587994 378088 589183
rect 378048 587988 378100 587994
rect 378048 587930 378100 587936
rect 377862 587616 377918 587625
rect 377862 587551 377918 587560
rect 377876 587110 377904 587551
rect 377864 587104 377916 587110
rect 377864 587046 377916 587052
rect 377862 586800 377918 586809
rect 377862 586735 377918 586744
rect 377876 586702 377904 586735
rect 377864 586696 377916 586702
rect 377864 586638 377916 586644
rect 377220 585268 377272 585274
rect 377220 585210 377272 585216
rect 377232 585177 377260 585210
rect 377218 585168 377274 585177
rect 377218 585103 377274 585112
rect 377770 584352 377826 584361
rect 377770 584287 377826 584296
rect 377784 583778 377812 584287
rect 377772 583772 377824 583778
rect 377772 583714 377824 583720
rect 378046 583536 378102 583545
rect 378046 583471 378102 583480
rect 378060 582826 378088 583471
rect 378048 582820 378100 582826
rect 378048 582762 378100 582768
rect 378046 582720 378102 582729
rect 378046 582655 378102 582664
rect 378060 582486 378088 582655
rect 378048 582480 378100 582486
rect 378048 582422 378100 582428
rect 378046 581088 378102 581097
rect 378046 581023 378048 581032
rect 378100 581023 378102 581032
rect 378048 580994 378100 581000
rect 378046 580272 378102 580281
rect 378046 580207 378102 580216
rect 378060 579698 378088 580207
rect 378048 579692 378100 579698
rect 378048 579634 378100 579640
rect 378046 578640 378102 578649
rect 378046 578575 378102 578584
rect 378060 578338 378088 578575
rect 378048 578332 378100 578338
rect 378048 578274 378100 578280
rect 378046 574560 378102 574569
rect 378046 574495 378102 574504
rect 378060 574122 378088 574495
rect 378048 574116 378100 574122
rect 378048 574058 378100 574064
rect 377586 572928 377642 572937
rect 377586 572863 377642 572872
rect 377600 572762 377628 572863
rect 377588 572756 377640 572762
rect 377588 572698 377640 572704
rect 377954 569664 378010 569673
rect 377954 569599 378010 569608
rect 377968 568614 377996 569599
rect 377956 568608 378008 568614
rect 377956 568550 378008 568556
rect 377128 558204 377180 558210
rect 377128 558146 377180 558152
rect 377036 557456 377088 557462
rect 377036 557398 377088 557404
rect 376850 529272 376906 529281
rect 376850 529207 376906 529216
rect 375840 528352 375892 528358
rect 375840 528294 375892 528300
rect 378152 524346 378180 615466
rect 378244 529922 378272 619670
rect 378322 617808 378378 617817
rect 378322 617743 378378 617752
rect 378232 529916 378284 529922
rect 378232 529858 378284 529864
rect 378336 529718 378364 617743
rect 378690 613728 378746 613737
rect 378690 613663 378746 613672
rect 378414 612912 378470 612921
rect 378414 612847 378470 612856
rect 378324 529712 378376 529718
rect 378324 529654 378376 529660
rect 378428 528562 378456 612847
rect 378598 599856 378654 599865
rect 378598 599791 378654 599800
rect 378506 595776 378562 595785
rect 378506 595711 378562 595720
rect 378416 528556 378468 528562
rect 378416 528498 378468 528504
rect 378140 524340 378192 524346
rect 378140 524282 378192 524288
rect 377126 524240 377182 524249
rect 375748 524204 375800 524210
rect 377126 524175 377182 524184
rect 375748 524146 375800 524152
rect 375564 522844 375616 522850
rect 375564 522786 375616 522792
rect 375470 519752 375526 519761
rect 375470 519687 375526 519696
rect 374644 518220 374696 518226
rect 374644 518162 374696 518168
rect 375484 518106 375512 519687
rect 377140 518106 377168 524175
rect 378520 522782 378548 595711
rect 378612 528426 378640 599791
rect 378704 556170 378732 613663
rect 378692 556164 378744 556170
rect 378692 556106 378744 556112
rect 378600 528420 378652 528426
rect 378600 528362 378652 528368
rect 379532 525774 379560 620978
rect 379796 587920 379848 587926
rect 379796 587862 379848 587868
rect 379704 585200 379756 585206
rect 379704 585142 379756 585148
rect 379610 577824 379666 577833
rect 379610 577759 379666 577768
rect 379624 534177 379652 577759
rect 379716 557530 379744 585142
rect 379808 559842 379836 587862
rect 379980 585268 380032 585274
rect 379980 585210 380032 585216
rect 379888 578264 379940 578270
rect 379888 578206 379940 578212
rect 379796 559836 379848 559842
rect 379796 559778 379848 559784
rect 379704 557524 379756 557530
rect 379704 557466 379756 557472
rect 379900 551886 379928 578206
rect 379992 559910 380020 585210
rect 380900 572756 380952 572762
rect 380900 572698 380952 572704
rect 379980 559904 380032 559910
rect 379980 559846 380032 559852
rect 379888 551880 379940 551886
rect 379888 551822 379940 551828
rect 380912 550458 380940 572698
rect 380900 550452 380952 550458
rect 380900 550394 380952 550400
rect 380254 544912 380310 544921
rect 380254 544847 380310 544856
rect 379610 534168 379666 534177
rect 379610 534103 379666 534112
rect 379520 525768 379572 525774
rect 379520 525710 379572 525716
rect 378508 522776 378560 522782
rect 378508 522718 378560 522724
rect 378598 521384 378654 521393
rect 378598 521319 378654 521328
rect 373920 518078 373964 518106
rect 375484 518078 375528 518106
rect 372372 517956 372400 518078
rect 373936 517956 373964 518078
rect 375500 517956 375528 518078
rect 377064 518078 377168 518106
rect 378612 518106 378640 521319
rect 380268 518106 380296 544847
rect 381004 524414 381032 625534
rect 381084 623824 381136 623830
rect 381084 623766 381136 623772
rect 381096 538218 381124 623766
rect 381176 622464 381228 622470
rect 381176 622406 381228 622412
rect 381188 545086 381216 622406
rect 381452 587104 381504 587110
rect 381452 587046 381504 587052
rect 381360 586696 381412 586702
rect 381360 586638 381412 586644
rect 381268 583772 381320 583778
rect 381268 583714 381320 583720
rect 381280 559774 381308 583714
rect 381268 559768 381320 559774
rect 381268 559710 381320 559716
rect 381372 558890 381400 586638
rect 381464 559706 381492 587046
rect 381452 559700 381504 559706
rect 381452 559642 381504 559648
rect 381360 558884 381412 558890
rect 381360 558826 381412 558832
rect 381176 545080 381228 545086
rect 381176 545022 381228 545028
rect 381084 538212 381136 538218
rect 381084 538154 381136 538160
rect 380992 524408 381044 524414
rect 380992 524350 381044 524356
rect 381556 521014 381584 637638
rect 384302 622976 384358 622985
rect 384302 622911 384358 622920
rect 384316 611425 384344 622911
rect 400876 617574 400904 640222
rect 410536 632058 410564 640290
rect 453304 632732 453356 632738
rect 453304 632674 453356 632680
rect 410524 632052 410576 632058
rect 410524 631994 410576 632000
rect 413284 632052 413336 632058
rect 413284 631994 413336 632000
rect 400864 617568 400916 617574
rect 400864 617510 400916 617516
rect 413296 612814 413324 631994
rect 426348 617568 426400 617574
rect 426348 617510 426400 617516
rect 413284 612808 413336 612814
rect 413284 612750 413336 612756
rect 416044 612808 416096 612814
rect 416044 612750 416096 612756
rect 384302 611416 384358 611425
rect 384302 611351 384358 611360
rect 391202 611416 391258 611425
rect 391202 611351 391258 611360
rect 385040 605872 385092 605878
rect 385040 605814 385092 605820
rect 383660 592136 383712 592142
rect 383660 592078 383712 592084
rect 382648 587988 382700 587994
rect 382648 587930 382700 587936
rect 382372 582820 382424 582826
rect 382372 582762 382424 582768
rect 382278 581904 382334 581913
rect 382278 581839 382334 581848
rect 381636 568608 381688 568614
rect 381636 568550 381688 568556
rect 381648 537946 381676 568550
rect 381818 557288 381874 557297
rect 381818 557223 381874 557232
rect 381636 537940 381688 537946
rect 381636 537882 381688 537888
rect 381544 521008 381596 521014
rect 381544 520950 381596 520956
rect 381832 518106 381860 557223
rect 382292 518129 382320 581839
rect 382384 524074 382412 582762
rect 382464 579692 382516 579698
rect 382464 579634 382516 579640
rect 382372 524068 382424 524074
rect 382372 524010 382424 524016
rect 382476 521422 382504 579634
rect 382556 578332 382608 578338
rect 382556 578274 382608 578280
rect 382568 522646 382596 578274
rect 382660 546106 382688 587930
rect 383382 557016 383438 557025
rect 383382 556951 383438 556960
rect 382648 546100 382700 546106
rect 382648 546042 382700 546048
rect 382556 522640 382608 522646
rect 382556 522582 382608 522588
rect 382464 521416 382516 521422
rect 382464 521358 382516 521364
rect 378612 518078 378656 518106
rect 377064 517956 377092 518078
rect 378628 517956 378656 518078
rect 380192 518078 380296 518106
rect 381756 518078 381860 518106
rect 382278 518120 382334 518129
rect 380192 517956 380220 518078
rect 381756 517956 381784 518078
rect 383396 518106 383424 556951
rect 383672 521558 383700 592078
rect 383842 591696 383898 591705
rect 383842 591631 383898 591640
rect 383752 581052 383804 581058
rect 383752 580994 383804 581000
rect 383660 521552 383712 521558
rect 383660 521494 383712 521500
rect 383764 520198 383792 580994
rect 383856 530641 383884 591631
rect 383936 582480 383988 582486
rect 383936 582422 383988 582428
rect 383842 530632 383898 530641
rect 383842 530567 383898 530576
rect 383948 524142 383976 582422
rect 383936 524136 383988 524142
rect 383936 524078 383988 524084
rect 384854 521112 384910 521121
rect 384854 521047 384910 521056
rect 383752 520192 383804 520198
rect 383752 520134 383804 520140
rect 382278 518055 382334 518064
rect 383320 518078 383424 518106
rect 384868 518106 384896 521047
rect 385052 519926 385080 605814
rect 386420 604580 386472 604586
rect 386420 604522 386472 604528
rect 385132 603288 385184 603294
rect 385132 603230 385184 603236
rect 385144 521626 385172 603230
rect 385224 594856 385276 594862
rect 385224 594798 385276 594804
rect 385132 521620 385184 521626
rect 385132 521562 385184 521568
rect 385040 519920 385092 519926
rect 385040 519862 385092 519868
rect 385236 518770 385264 594798
rect 385408 590708 385460 590714
rect 385408 590650 385460 590656
rect 385316 589688 385368 589694
rect 385316 589630 385368 589636
rect 385328 521490 385356 589630
rect 385420 522918 385448 590650
rect 385408 522912 385460 522918
rect 385408 522854 385460 522860
rect 385316 521484 385368 521490
rect 385316 521426 385368 521432
rect 386432 518838 386460 604522
rect 389180 604512 389232 604518
rect 389180 604454 389232 604460
rect 386604 603152 386656 603158
rect 386604 603094 386656 603100
rect 386510 556880 386566 556889
rect 386510 556815 386566 556824
rect 386420 518832 386472 518838
rect 386420 518774 386472 518780
rect 385224 518764 385276 518770
rect 385224 518706 385276 518712
rect 386524 518106 386552 556815
rect 386616 522986 386644 603094
rect 386696 592068 386748 592074
rect 386696 592010 386748 592016
rect 386708 525638 386736 592010
rect 386788 574116 386840 574122
rect 386788 574058 386840 574064
rect 386800 542298 386828 574058
rect 388074 556744 388130 556753
rect 388074 556679 388130 556688
rect 386788 542292 386840 542298
rect 386788 542234 386840 542240
rect 386696 525632 386748 525638
rect 386696 525574 386748 525580
rect 386604 522980 386656 522986
rect 386604 522922 386656 522928
rect 388088 518106 388116 556679
rect 389192 518906 389220 604454
rect 391216 599593 391244 611351
rect 391202 599584 391258 599593
rect 391202 599519 391258 599528
rect 403622 599584 403678 599593
rect 403622 599519 403678 599528
rect 403636 583001 403664 599519
rect 416056 584798 416084 612750
rect 426360 609278 426388 617510
rect 453316 613426 453344 632674
rect 453304 613420 453356 613426
rect 453304 613362 453356 613368
rect 426348 609272 426400 609278
rect 426348 609214 426400 609220
rect 442264 609272 442316 609278
rect 442264 609214 442316 609220
rect 442276 594862 442304 609214
rect 442264 594856 442316 594862
rect 442264 594798 442316 594804
rect 448520 594856 448572 594862
rect 448520 594798 448572 594804
rect 448532 591326 448560 594798
rect 448520 591320 448572 591326
rect 448520 591262 448572 591268
rect 454684 591320 454736 591326
rect 454684 591262 454736 591268
rect 416044 584792 416096 584798
rect 416044 584734 416096 584740
rect 423588 584792 423640 584798
rect 423588 584734 423640 584740
rect 403622 582992 403678 583001
rect 403622 582927 403678 582936
rect 423600 580310 423628 584734
rect 427082 582992 427138 583001
rect 427082 582927 427138 582936
rect 423588 580304 423640 580310
rect 423588 580246 423640 580252
rect 427096 578377 427124 582927
rect 432604 580304 432656 580310
rect 432604 580246 432656 580252
rect 427082 578368 427138 578377
rect 427082 578303 427138 578312
rect 431958 578368 432014 578377
rect 431958 578303 432014 578312
rect 431972 572801 432000 578303
rect 431958 572792 432014 572801
rect 431958 572727 432014 572736
rect 408406 559736 408462 559745
rect 408406 559671 408462 559680
rect 406842 551712 406898 551721
rect 406842 551647 406898 551656
rect 400586 543552 400642 543561
rect 400586 543487 400642 543496
rect 389638 539336 389694 539345
rect 389638 539271 389694 539280
rect 389180 518900 389232 518906
rect 389180 518842 389232 518848
rect 389652 518106 389680 539271
rect 397366 536752 397422 536761
rect 397366 536687 397422 536696
rect 395894 534032 395950 534041
rect 395894 533967 395950 533976
rect 394330 532672 394386 532681
rect 394330 532607 394386 532616
rect 392766 524104 392822 524113
rect 392766 524039 392822 524048
rect 391110 521248 391166 521257
rect 391110 521183 391166 521192
rect 384868 518078 384912 518106
rect 383320 517956 383348 518078
rect 384884 517956 384912 518078
rect 386448 518078 386552 518106
rect 388012 518078 388116 518106
rect 389576 518078 389680 518106
rect 391124 518106 391152 521183
rect 392780 518106 392808 524039
rect 394344 518106 394372 532607
rect 395908 518106 395936 533967
rect 391124 518078 391168 518106
rect 386448 517956 386476 518078
rect 388012 517956 388040 518078
rect 389576 517956 389604 518078
rect 391140 517956 391168 518078
rect 392704 518078 392808 518106
rect 394268 518078 394372 518106
rect 395832 518078 395936 518106
rect 397380 518106 397408 536687
rect 399022 536616 399078 536625
rect 399022 536551 399078 536560
rect 399036 518106 399064 536551
rect 400600 518106 400628 543487
rect 403716 532160 403768 532166
rect 403716 532102 403768 532108
rect 402150 525464 402206 525473
rect 402150 525399 402206 525408
rect 402164 518106 402192 525399
rect 403728 518106 403756 532102
rect 405278 522744 405334 522753
rect 405278 522679 405334 522688
rect 405292 518106 405320 522679
rect 406856 518106 406884 551647
rect 408420 518106 408448 559671
rect 420826 559600 420882 559609
rect 420826 559535 420882 559544
rect 416226 547360 416282 547369
rect 416226 547295 416282 547304
rect 414662 546272 414718 546281
rect 414662 546207 414718 546216
rect 413098 542192 413154 542201
rect 413098 542127 413154 542136
rect 409970 540968 410026 540977
rect 409970 540903 410026 540912
rect 409984 518106 410012 540903
rect 411534 528320 411590 528329
rect 411534 528255 411590 528264
rect 411548 518106 411576 528255
rect 413112 518106 413140 542127
rect 414676 518106 414704 546207
rect 416240 518106 416268 547295
rect 417790 544504 417846 544513
rect 417790 544439 417846 544448
rect 417804 518106 417832 544439
rect 419354 537704 419410 537713
rect 419354 537639 419410 537648
rect 419368 518106 419396 537639
rect 397380 518078 397424 518106
rect 392704 517956 392732 518078
rect 394268 517956 394296 518078
rect 395832 517956 395860 518078
rect 397396 517956 397424 518078
rect 398960 518078 399064 518106
rect 400524 518078 400628 518106
rect 402088 518078 402192 518106
rect 403652 518078 403756 518106
rect 405216 518078 405320 518106
rect 406780 518078 406884 518106
rect 408344 518078 408448 518106
rect 409908 518078 410012 518106
rect 411472 518078 411576 518106
rect 413036 518078 413140 518106
rect 414600 518078 414704 518106
rect 416164 518078 416268 518106
rect 417728 518078 417832 518106
rect 419292 518078 419396 518106
rect 420840 518106 420868 559535
rect 424048 556844 424100 556850
rect 424048 556786 424100 556792
rect 422484 556232 422536 556238
rect 422484 556174 422536 556180
rect 422496 518106 422524 556174
rect 424060 518106 424088 556786
rect 432616 548690 432644 580246
rect 454696 574802 454724 591262
rect 454684 574796 454736 574802
rect 454684 574738 454736 574744
rect 435362 572792 435418 572801
rect 435362 572727 435418 572736
rect 435376 560289 435404 572727
rect 435362 560280 435418 560289
rect 435362 560215 435418 560224
rect 437662 560280 437718 560289
rect 437662 560215 437718 560224
rect 437676 553353 437704 560215
rect 453762 555656 453818 555665
rect 453762 555591 453818 555600
rect 437662 553344 437718 553353
rect 437662 553279 437718 553288
rect 439688 552288 439740 552294
rect 439688 552230 439740 552236
rect 434994 550080 435050 550089
rect 434994 550015 435050 550024
rect 432604 548684 432656 548690
rect 432604 548626 432656 548632
rect 430302 548584 430358 548593
rect 430302 548519 430358 548528
rect 428738 541648 428794 541657
rect 428738 541583 428794 541592
rect 427084 534268 427136 534274
rect 427084 534210 427136 534216
rect 425610 528184 425666 528193
rect 425610 528119 425666 528128
rect 425624 518106 425652 528119
rect 427096 521014 427124 534210
rect 427174 533624 427230 533633
rect 427174 533559 427230 533568
rect 427084 521008 427136 521014
rect 427084 520950 427136 520956
rect 427188 518106 427216 533559
rect 428752 518106 428780 541583
rect 430316 518106 430344 548519
rect 433432 526448 433484 526454
rect 433432 526390 433484 526396
rect 431684 520328 431736 520334
rect 431684 520270 431736 520276
rect 431696 518894 431724 520270
rect 431696 518866 431816 518894
rect 420840 518078 420884 518106
rect 398960 517956 398988 518078
rect 400524 517956 400552 518078
rect 402088 517956 402116 518078
rect 403652 517956 403680 518078
rect 405216 517956 405244 518078
rect 406780 517956 406808 518078
rect 408344 517956 408372 518078
rect 409908 517956 409936 518078
rect 411472 517956 411500 518078
rect 413036 517956 413064 518078
rect 414600 517956 414628 518078
rect 416164 517956 416192 518078
rect 417728 517956 417756 518078
rect 419292 517956 419320 518078
rect 420856 517956 420884 518078
rect 422420 518078 422524 518106
rect 423984 518078 424088 518106
rect 425548 518078 425652 518106
rect 427112 518078 427216 518106
rect 428676 518078 428780 518106
rect 430240 518078 430344 518106
rect 431788 518106 431816 518866
rect 433444 518106 433472 526390
rect 435008 518106 435036 550015
rect 436560 543788 436612 543794
rect 436560 543730 436612 543736
rect 436572 518106 436600 543730
rect 438122 537568 438178 537577
rect 438122 537503 438178 537512
rect 438136 518106 438164 537503
rect 439700 518106 439728 552230
rect 443644 548684 443696 548690
rect 443644 548626 443696 548632
rect 443656 540530 443684 548626
rect 452198 545728 452254 545737
rect 452198 545663 452254 545672
rect 444286 543008 444342 543017
rect 444286 542943 444342 542952
rect 443644 540524 443696 540530
rect 443644 540466 443696 540472
rect 442814 540288 442870 540297
rect 442814 540223 442870 540232
rect 441250 528048 441306 528057
rect 441250 527983 441306 527992
rect 441264 518106 441292 527983
rect 442828 518106 442856 540223
rect 431788 518078 431832 518106
rect 422420 517956 422448 518078
rect 423984 517956 424012 518078
rect 425548 517956 425576 518078
rect 427112 517956 427140 518078
rect 428676 517956 428704 518078
rect 430240 517956 430268 518078
rect 431804 517956 431832 518078
rect 433368 518078 433472 518106
rect 434932 518078 435036 518106
rect 436496 518078 436600 518106
rect 438060 518078 438164 518106
rect 439624 518078 439728 518106
rect 441188 518078 441292 518106
rect 442752 518078 442856 518106
rect 444300 518106 444328 542943
rect 447508 538280 447560 538286
rect 447508 538222 447560 538228
rect 445942 537432 445998 537441
rect 445942 537367 445998 537376
rect 445956 518106 445984 537367
rect 447520 518106 447548 538222
rect 450636 532092 450688 532098
rect 450636 532034 450688 532040
rect 449070 531176 449126 531185
rect 449070 531111 449126 531120
rect 449084 518106 449112 531111
rect 450648 518106 450676 532034
rect 452212 518106 452240 545663
rect 453304 540524 453356 540530
rect 453304 540466 453356 540472
rect 453316 526454 453344 540466
rect 453304 526448 453356 526454
rect 453304 526390 453356 526396
rect 453776 518106 453804 555591
rect 456892 546508 456944 546514
rect 456892 546450 456944 546456
rect 455328 532024 455380 532030
rect 455328 531966 455380 531972
rect 455340 518106 455368 531966
rect 456904 518106 456932 546450
rect 461492 534812 461544 534818
rect 461492 534754 461544 534760
rect 460018 528728 460074 528737
rect 460018 528663 460074 528672
rect 458454 527776 458510 527785
rect 458454 527711 458510 527720
rect 458468 518106 458496 527711
rect 460032 518106 460060 528663
rect 444300 518078 444344 518106
rect 433368 517956 433396 518078
rect 434932 517956 434960 518078
rect 436496 517956 436524 518078
rect 438060 517956 438088 518078
rect 439624 517956 439652 518078
rect 441188 517956 441216 518078
rect 442752 517956 442780 518078
rect 444316 517956 444344 518078
rect 445880 518078 445984 518106
rect 447444 518078 447548 518106
rect 449008 518078 449112 518106
rect 450572 518078 450676 518106
rect 452136 518078 452240 518106
rect 453700 518078 453804 518106
rect 455264 518078 455368 518106
rect 456828 518078 456932 518106
rect 458392 518078 458496 518106
rect 459956 518078 460060 518106
rect 461504 518106 461532 534754
rect 461596 518401 461624 644807
rect 461688 521121 461716 647527
rect 461768 645992 461820 645998
rect 461768 645934 461820 645940
rect 461674 521112 461730 521121
rect 461780 521082 461808 645934
rect 461858 645008 461914 645017
rect 461858 644943 461914 644952
rect 461872 521257 461900 644943
rect 462332 599593 462360 703520
rect 473266 656024 473322 656033
rect 473266 655959 473322 655968
rect 467286 647456 467342 647465
rect 467286 647391 467342 647400
rect 467102 647320 467158 647329
rect 467102 647255 467158 647264
rect 464342 646776 464398 646785
rect 464342 646711 464398 646720
rect 462962 639568 463018 639577
rect 462962 639503 463018 639512
rect 462318 599584 462374 599593
rect 462318 599519 462374 599528
rect 462226 553344 462282 553353
rect 462226 553279 462282 553288
rect 462240 550089 462268 553279
rect 462226 550080 462282 550089
rect 462226 550015 462282 550024
rect 461858 521248 461914 521257
rect 461858 521183 461914 521192
rect 461674 521047 461730 521056
rect 461768 521076 461820 521082
rect 461768 521018 461820 521024
rect 462976 519761 463004 639503
rect 463148 535560 463200 535566
rect 463148 535502 463200 535508
rect 462962 519752 463018 519761
rect 462962 519687 463018 519696
rect 461582 518392 461638 518401
rect 461582 518327 461638 518336
rect 463160 518106 463188 535502
rect 463608 526448 463660 526454
rect 463608 526390 463660 526396
rect 463620 522986 463648 526390
rect 463608 522980 463660 522986
rect 463608 522922 463660 522928
rect 464356 522617 464384 646711
rect 464436 640484 464488 640490
rect 464436 640426 464488 640432
rect 464342 522608 464398 522617
rect 464342 522543 464398 522552
rect 464448 522374 464476 640426
rect 465816 636676 465868 636682
rect 465816 636618 465868 636624
rect 464618 636576 464674 636585
rect 464618 636511 464674 636520
rect 464526 634944 464582 634953
rect 464526 634879 464582 634888
rect 464436 522368 464488 522374
rect 464436 522310 464488 522316
rect 464540 521393 464568 634879
rect 464632 522753 464660 636511
rect 465724 635248 465776 635254
rect 465724 635190 465776 635196
rect 464712 534744 464764 534750
rect 464712 534686 464764 534692
rect 464618 522744 464674 522753
rect 464618 522679 464674 522688
rect 464526 521384 464582 521393
rect 464526 521319 464582 521328
rect 464724 518106 464752 534686
rect 465736 522442 465764 635190
rect 465828 525094 465856 636618
rect 466276 542428 466328 542434
rect 466276 542370 466328 542376
rect 465816 525088 465868 525094
rect 465816 525030 465868 525036
rect 465724 522436 465776 522442
rect 465724 522378 465776 522384
rect 466288 518106 466316 542370
rect 467116 519654 467144 647255
rect 467196 643476 467248 643482
rect 467196 643418 467248 643424
rect 467208 519722 467236 643418
rect 467300 519790 467328 647391
rect 471244 647352 471296 647358
rect 471244 647294 471296 647300
rect 468484 647284 468536 647290
rect 468484 647226 468536 647232
rect 467746 555520 467802 555529
rect 467746 555455 467802 555464
rect 467288 519784 467340 519790
rect 467288 519726 467340 519732
rect 467196 519716 467248 519722
rect 467196 519658 467248 519664
rect 467104 519648 467156 519654
rect 467104 519590 467156 519596
rect 461504 518078 461548 518106
rect 445880 517956 445908 518078
rect 447444 517956 447472 518078
rect 449008 517956 449036 518078
rect 450572 517956 450600 518078
rect 452136 517956 452164 518078
rect 453700 517956 453728 518078
rect 455264 517956 455292 518078
rect 456828 517956 456856 518078
rect 458392 517956 458420 518078
rect 459956 517956 459984 518078
rect 461520 517956 461548 518078
rect 463084 518078 463188 518106
rect 464648 518078 464752 518106
rect 466212 518078 466316 518106
rect 467760 518106 467788 555455
rect 467840 522980 467892 522986
rect 467840 522922 467892 522928
rect 467852 520062 467880 522922
rect 468496 521218 468524 647226
rect 468576 637016 468628 637022
rect 468576 636958 468628 636964
rect 468484 521212 468536 521218
rect 468484 521154 468536 521160
rect 467840 520056 467892 520062
rect 467840 519998 467892 520004
rect 468588 519586 468616 636958
rect 468668 636608 468720 636614
rect 468668 636550 468720 636556
rect 468680 521150 468708 636550
rect 468760 636540 468812 636546
rect 468760 636482 468812 636488
rect 468772 522306 468800 636482
rect 469404 550792 469456 550798
rect 469404 550734 469456 550740
rect 468760 522300 468812 522306
rect 468760 522242 468812 522248
rect 468668 521144 468720 521150
rect 468668 521086 468720 521092
rect 468576 519580 468628 519586
rect 468576 519522 468628 519528
rect 469416 518106 469444 550734
rect 470968 540388 471020 540394
rect 470968 540330 471020 540336
rect 470980 518106 471008 540330
rect 471256 519926 471284 647294
rect 471336 645924 471388 645930
rect 471336 645866 471388 645872
rect 471348 521286 471376 645866
rect 472622 643648 472678 643657
rect 472622 643583 472678 643592
rect 471518 637800 471574 637809
rect 471518 637735 471574 637744
rect 471426 635080 471482 635089
rect 471426 635015 471482 635024
rect 471336 521280 471388 521286
rect 471336 521222 471388 521228
rect 471244 519920 471296 519926
rect 471244 519862 471296 519868
rect 471440 519858 471468 635015
rect 471532 522073 471560 637735
rect 471610 550080 471666 550089
rect 471610 550015 471666 550024
rect 471624 524385 471652 550015
rect 472532 527196 472584 527202
rect 472532 527138 472584 527144
rect 471610 524376 471666 524385
rect 471610 524311 471666 524320
rect 471886 523016 471942 523025
rect 471886 522951 471942 522960
rect 471518 522064 471574 522073
rect 471518 521999 471574 522008
rect 471900 521762 471928 522951
rect 471888 521756 471940 521762
rect 471888 521698 471940 521704
rect 471428 519852 471480 519858
rect 471428 519794 471480 519800
rect 472544 518106 472572 527138
rect 472636 521529 472664 643583
rect 473280 521665 473308 655959
rect 476026 655888 476082 655897
rect 476026 655823 476082 655832
rect 475934 654664 475990 654673
rect 475934 654599 475990 654608
rect 474004 643136 474056 643142
rect 474004 643078 474056 643084
rect 473358 524376 473414 524385
rect 473358 524311 473414 524320
rect 473266 521656 473322 521665
rect 473266 521591 473322 521600
rect 472622 521520 472678 521529
rect 472622 521455 472678 521464
rect 473372 520849 473400 524311
rect 474016 523682 474044 643078
rect 474096 642048 474148 642054
rect 474096 641990 474148 641996
rect 474108 538214 474136 641990
rect 475384 574796 475436 574802
rect 475384 574738 475436 574744
rect 474108 538186 474320 538214
rect 474016 523654 474136 523682
rect 474004 520940 474056 520946
rect 474004 520882 474056 520888
rect 473358 520840 473414 520849
rect 473358 520775 473414 520784
rect 467760 518078 467804 518106
rect 463084 517956 463112 518078
rect 464648 517956 464676 518078
rect 466212 517956 466240 518078
rect 467776 517956 467804 518078
rect 469340 518078 469444 518106
rect 470904 518078 471008 518106
rect 472468 518078 472572 518106
rect 474016 518106 474044 520882
rect 474108 518226 474136 523654
rect 474292 522578 474320 538186
rect 474280 522572 474332 522578
rect 474280 522514 474332 522520
rect 475396 520266 475424 574738
rect 475948 522510 475976 654599
rect 475936 522504 475988 522510
rect 475936 522446 475988 522452
rect 475476 521008 475528 521014
rect 475476 520950 475528 520956
rect 475384 520260 475436 520266
rect 475384 520202 475436 520208
rect 475488 518894 475516 520950
rect 476040 519994 476068 655823
rect 477406 655752 477462 655761
rect 477406 655687 477462 655696
rect 476764 635044 476816 635050
rect 476764 634986 476816 634992
rect 476028 519988 476080 519994
rect 476028 519930 476080 519936
rect 475488 518866 475608 518894
rect 474096 518220 474148 518226
rect 474096 518162 474148 518168
rect 475580 518106 475608 518866
rect 476118 518392 476174 518401
rect 476118 518327 476174 518336
rect 476132 518158 476160 518327
rect 476776 518294 476804 634986
rect 476946 547088 477002 547097
rect 476946 547023 477002 547032
rect 476764 518288 476816 518294
rect 476960 518265 476988 547023
rect 477420 522646 477448 655687
rect 477500 613420 477552 613426
rect 477500 613362 477552 613368
rect 477512 612814 477540 613362
rect 477500 612808 477552 612814
rect 477500 612750 477552 612756
rect 478524 599729 478552 703520
rect 486974 657792 487030 657801
rect 478880 657756 478932 657762
rect 478880 657698 478932 657704
rect 485596 657756 485648 657762
rect 494808 657762 494836 703520
rect 508502 700360 508558 700369
rect 527192 700330 527220 703520
rect 508502 700295 508558 700304
rect 527180 700324 527232 700330
rect 507124 670744 507176 670750
rect 507124 670686 507176 670692
rect 501786 657792 501842 657801
rect 486974 657727 487030 657736
rect 494796 657756 494848 657762
rect 485596 657698 485648 657704
rect 478892 657150 478920 657698
rect 484030 657384 484086 657393
rect 484030 657319 484086 657328
rect 478880 657144 478932 657150
rect 478880 657086 478932 657092
rect 480168 657144 480220 657150
rect 480168 657086 480220 657092
rect 479432 641980 479484 641986
rect 479432 641922 479484 641928
rect 479340 639328 479392 639334
rect 479246 639296 479302 639305
rect 479340 639270 479392 639276
rect 479246 639231 479302 639240
rect 478788 612808 478840 612814
rect 478788 612750 478840 612756
rect 478510 599720 478566 599729
rect 478510 599655 478566 599664
rect 477408 522640 477460 522646
rect 477408 522582 477460 522588
rect 478800 518894 478828 612750
rect 478800 518866 479012 518894
rect 477406 518800 477462 518809
rect 477406 518735 477462 518744
rect 478786 518800 478842 518809
rect 478786 518735 478842 518744
rect 477420 518498 477448 518735
rect 478800 518566 478828 518735
rect 478788 518560 478840 518566
rect 478788 518502 478840 518508
rect 477408 518492 477460 518498
rect 477408 518434 477460 518440
rect 477316 518424 477368 518430
rect 477316 518366 477368 518372
rect 476764 518230 476816 518236
rect 476946 518256 477002 518265
rect 476946 518191 477002 518200
rect 476120 518152 476172 518158
rect 474016 518078 474060 518106
rect 475580 518078 475624 518106
rect 477328 518129 477356 518366
rect 478510 518256 478566 518265
rect 478510 518191 478566 518200
rect 476120 518094 476172 518100
rect 477314 518120 477370 518129
rect 469340 517956 469368 518078
rect 470904 517956 470932 518078
rect 472468 517956 472496 518078
rect 474032 517956 474060 518078
rect 475596 517956 475624 518078
rect 477314 518055 477370 518064
rect 61566 517919 61622 517928
rect 478524 517857 478552 518191
rect 478786 518120 478842 518129
rect 478786 518055 478788 518064
rect 478840 518055 478842 518064
rect 478788 518026 478840 518032
rect 478984 518022 479012 518866
rect 478972 518016 479024 518022
rect 478972 517958 479024 517964
rect 478510 517848 478566 517857
rect 478510 517783 478566 517792
rect 60924 517676 60976 517682
rect 60924 517618 60976 517624
rect 60832 517608 60884 517614
rect 60832 517550 60884 517556
rect 60740 517540 60792 517546
rect 60740 517482 60792 517488
rect 479260 478038 479288 639231
rect 479248 478032 479300 478038
rect 479248 477974 479300 477980
rect 479352 467401 479380 639270
rect 479338 467392 479394 467401
rect 479338 467327 479394 467336
rect 479444 453257 479472 641922
rect 479982 637664 480038 637673
rect 479982 637599 480038 637608
rect 479890 539064 479946 539073
rect 479890 538999 479946 539008
rect 479616 529984 479668 529990
rect 479616 529926 479668 529932
rect 479524 478032 479576 478038
rect 479524 477974 479576 477980
rect 479536 476105 479564 477974
rect 479522 476096 479578 476105
rect 479522 476031 479578 476040
rect 479430 453248 479486 453257
rect 479430 453183 479486 453192
rect 479522 449984 479578 449993
rect 479522 449919 479578 449928
rect 94134 390144 94190 390153
rect 60738 389056 60794 389065
rect 60738 388991 60794 389000
rect 60646 387696 60702 387705
rect 60646 387631 60702 387640
rect 60556 387524 60608 387530
rect 60556 387466 60608 387472
rect 60462 387424 60518 387433
rect 60462 387359 60518 387368
rect 59266 387223 59322 387232
rect 60280 387252 60332 387258
rect 60280 387194 60332 387200
rect 60752 383761 60780 388991
rect 62118 387424 62174 387433
rect 62118 387359 62174 387368
rect 62132 387190 62160 387359
rect 62120 387184 62172 387190
rect 62120 387126 62172 387132
rect 62578 387016 62634 387025
rect 62578 386951 62634 386960
rect 60922 386880 60978 386889
rect 60922 386815 60978 386824
rect 60738 383752 60794 383761
rect 60738 383687 60794 383696
rect 58624 341692 58676 341698
rect 58624 341634 58676 341640
rect 59266 298752 59322 298761
rect 59266 298687 59322 298696
rect 54668 263016 54720 263022
rect 50986 262984 51042 262993
rect 54668 262958 54720 262964
rect 50986 262919 51042 262928
rect 39948 261520 40000 261526
rect 39948 261462 40000 261468
rect 47582 261216 47638 261225
rect 47582 261151 47638 261160
rect 40682 261080 40738 261089
rect 40682 261015 40738 261024
rect 35162 260944 35218 260953
rect 11704 260908 11756 260914
rect 35162 260879 35218 260888
rect 11704 260850 11756 260856
rect 11716 215286 11744 260850
rect 11704 215280 11756 215286
rect 11704 215222 11756 215228
rect 15842 193896 15898 193905
rect 15842 193831 15898 193840
rect 14738 127664 14794 127673
rect 14738 127599 14794 127608
rect 11702 126304 11758 126313
rect 11702 126239 11758 126248
rect 8758 98696 8814 98705
rect 8758 98631 8814 98640
rect 4894 32872 4950 32881
rect 4894 32807 4950 32816
rect 4802 32464 4858 32473
rect 4802 32399 4858 32408
rect 4066 27024 4122 27033
rect 4066 26959 4122 26968
rect 4080 480 4108 26959
rect 4908 3505 4936 32807
rect 7654 4856 7710 4865
rect 7654 4791 7710 4800
rect 4894 3496 4950 3505
rect 4894 3431 4950 3440
rect 6458 3496 6514 3505
rect 6458 3431 6514 3440
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3431
rect 7668 480 7696 4791
rect 8772 480 8800 98631
rect 11716 3505 11744 126239
rect 13542 100056 13598 100065
rect 13542 99991 13598 100000
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 9954 3496 10010 3505
rect 9954 3431 10010 3440
rect 11702 3496 11758 3505
rect 11702 3431 11758 3440
rect 9968 480 9996 3431
rect 12360 480 12388 6151
rect 13556 480 13584 99991
rect 14752 480 14780 127599
rect 15856 3777 15884 193831
rect 31298 181384 31354 181393
rect 31298 181319 31354 181328
rect 23018 144120 23074 144129
rect 23018 144055 23074 144064
rect 17038 137728 17094 137737
rect 17038 137663 17094 137672
rect 15842 3768 15898 3777
rect 15842 3703 15898 3712
rect 17052 480 17080 137663
rect 21822 137592 21878 137601
rect 21822 137527 21878 137536
rect 18234 122224 18290 122233
rect 18234 122159 18290 122168
rect 18248 480 18276 122159
rect 19430 116512 19486 116521
rect 19430 116447 19486 116456
rect 19444 480 19472 116447
rect 21836 480 21864 137527
rect 23032 480 23060 144055
rect 26514 137864 26570 137873
rect 26514 137799 26570 137808
rect 24214 115152 24270 115161
rect 24214 115087 24270 115096
rect 24228 480 24256 115087
rect 26528 480 26556 137799
rect 30102 137184 30158 137193
rect 30102 137119 30158 137128
rect 28906 134464 28962 134473
rect 28906 134399 28962 134408
rect 27710 3496 27766 3505
rect 27710 3431 27766 3440
rect 27724 480 27752 3431
rect 28920 480 28948 134399
rect 30116 480 30144 137119
rect 31312 480 31340 181319
rect 33598 137048 33654 137057
rect 33598 136983 33654 136992
rect 32402 101416 32458 101425
rect 32402 101351 32458 101360
rect 32416 480 32444 101351
rect 33612 480 33640 136983
rect 34794 109712 34850 109721
rect 34794 109647 34850 109656
rect 34808 480 34836 109647
rect 35176 71641 35204 260879
rect 40696 162897 40724 261015
rect 40682 162888 40738 162897
rect 40682 162823 40738 162832
rect 44178 137728 44234 137737
rect 44178 137663 44234 137672
rect 44192 137630 44220 137663
rect 44180 137624 44232 137630
rect 44180 137566 44232 137572
rect 44270 137320 44326 137329
rect 44270 137255 44326 137264
rect 37186 136912 37242 136921
rect 37186 136847 37242 136856
rect 35990 120728 36046 120737
rect 35990 120663 36046 120672
rect 35254 112432 35310 112441
rect 35254 112367 35310 112376
rect 35162 71632 35218 71641
rect 35162 71567 35218 71576
rect 35268 3505 35296 112367
rect 35254 3496 35310 3505
rect 35254 3431 35310 3440
rect 36004 480 36032 120663
rect 37200 480 37228 136847
rect 40682 136776 40738 136785
rect 40682 136711 40738 136720
rect 38382 113792 38438 113801
rect 38382 113727 38438 113736
rect 38396 480 38424 113727
rect 39578 104136 39634 104145
rect 39578 104071 39634 104080
rect 39592 480 39620 104071
rect 40696 480 40724 136711
rect 43074 122088 43130 122097
rect 43074 122023 43130 122032
rect 41878 111072 41934 111081
rect 41878 111007 41934 111016
rect 41892 480 41920 111007
rect 43088 480 43116 122023
rect 44284 480 44312 137255
rect 45466 124944 45522 124953
rect 45466 124879 45522 124888
rect 45480 480 45508 124879
rect 47596 110673 47624 261151
rect 51000 260114 51028 262919
rect 52918 262848 52974 262857
rect 52918 262783 52974 262792
rect 50954 260086 51028 260114
rect 50954 259964 50982 260086
rect 52932 259978 52960 262783
rect 54680 259978 54708 262958
rect 56324 262948 56376 262954
rect 56324 262890 56376 262896
rect 56336 259978 56364 262890
rect 57888 262880 57940 262886
rect 57888 262822 57940 262828
rect 57900 259978 57928 262822
rect 59280 260250 59308 298687
rect 60936 260250 60964 386815
rect 62592 260250 62620 386951
rect 63498 383616 63554 383625
rect 63498 383551 63554 383560
rect 63512 375465 63540 383551
rect 63498 375456 63554 375465
rect 63498 375391 63554 375400
rect 65062 375456 65118 375465
rect 65062 375391 65118 375400
rect 65076 369753 65104 375391
rect 65062 369744 65118 369753
rect 65062 369679 65118 369688
rect 65444 338745 65472 390116
rect 67546 385656 67602 385665
rect 67546 385591 67602 385600
rect 65890 373280 65946 373289
rect 65890 373215 65946 373224
rect 65430 338736 65486 338745
rect 65430 338671 65486 338680
rect 65444 335354 65472 338671
rect 65444 335326 65564 335354
rect 64510 265568 64566 265577
rect 64510 265503 64566 265512
rect 52624 259950 52960 259978
rect 54280 259950 54708 259978
rect 55936 259950 56364 259978
rect 57592 259950 57928 259978
rect 59234 260222 59308 260250
rect 60890 260222 60964 260250
rect 62546 260222 62620 260250
rect 59234 259964 59262 260222
rect 60890 259964 60918 260222
rect 62546 259964 62574 260222
rect 64524 259978 64552 265503
rect 65536 262993 65564 335326
rect 65522 262984 65578 262993
rect 65522 262919 65578 262928
rect 65904 260250 65932 373215
rect 67560 260250 67588 385591
rect 69032 347041 69060 390116
rect 70306 369744 70362 369753
rect 70306 369679 70362 369688
rect 70320 368370 70348 369679
rect 70320 368342 70440 368370
rect 70412 366353 70440 368342
rect 70398 366344 70454 366353
rect 70398 366279 70454 366288
rect 72620 355366 72648 390116
rect 76208 364334 76236 390116
rect 77942 366344 77998 366353
rect 77942 366279 77998 366288
rect 76208 364306 76604 364334
rect 72608 355360 72660 355366
rect 72608 355302 72660 355308
rect 72620 354674 72648 355302
rect 72436 354646 72648 354674
rect 69018 347032 69074 347041
rect 69018 346967 69074 346976
rect 69032 345014 69060 346967
rect 69032 344986 69704 345014
rect 69204 271244 69256 271250
rect 69204 271186 69256 271192
rect 69216 260250 69244 271186
rect 69676 262857 69704 344986
rect 70860 279472 70912 279478
rect 70860 279414 70912 279420
rect 69662 262848 69718 262857
rect 69662 262783 69718 262792
rect 70872 260250 70900 279414
rect 72436 263022 72464 354646
rect 76576 344350 76604 364306
rect 77956 347721 77984 366279
rect 77942 347712 77998 347721
rect 77942 347647 77998 347656
rect 78862 347712 78918 347721
rect 78862 347647 78918 347656
rect 78876 344729 78904 347647
rect 78862 344720 78918 344729
rect 78862 344655 78918 344664
rect 76564 344344 76616 344350
rect 76564 344286 76616 344292
rect 75828 300144 75880 300150
rect 75828 300086 75880 300092
rect 74172 297424 74224 297430
rect 74172 297366 74224 297372
rect 72514 272640 72570 272649
rect 72514 272575 72570 272584
rect 72424 263016 72476 263022
rect 72424 262958 72476 262964
rect 72528 260250 72556 272575
rect 74184 260250 74212 297366
rect 75840 260250 75868 300086
rect 76576 262954 76604 344286
rect 79796 340202 79824 390116
rect 83384 383654 83412 390116
rect 86972 386889 87000 390116
rect 90560 388793 90588 390116
rect 94134 390079 94190 390088
rect 97276 390102 97750 390130
rect 90546 388784 90602 388793
rect 90546 388719 90602 388728
rect 90560 387025 90588 388719
rect 90546 387016 90602 387025
rect 90546 386951 90602 386960
rect 86958 386880 87014 386889
rect 86958 386815 87014 386824
rect 84108 384328 84160 384334
rect 84108 384270 84160 384276
rect 83384 383626 83504 383654
rect 83476 363633 83504 383626
rect 83462 363624 83518 363633
rect 83462 363559 83518 363568
rect 79324 340196 79376 340202
rect 79324 340138 79376 340144
rect 79784 340196 79836 340202
rect 79784 340138 79836 340144
rect 79138 301472 79194 301481
rect 79138 301407 79194 301416
rect 77484 282192 77536 282198
rect 77484 282134 77536 282140
rect 76564 262948 76616 262954
rect 76564 262890 76616 262896
rect 77496 260250 77524 282134
rect 79152 260250 79180 301407
rect 79336 262886 79364 340138
rect 82452 304292 82504 304298
rect 82452 304234 82504 304240
rect 80796 302932 80848 302938
rect 80796 302874 80848 302880
rect 79324 262880 79376 262886
rect 79324 262822 79376 262828
rect 80808 260250 80836 302874
rect 82464 260250 82492 304234
rect 83476 298761 83504 363559
rect 83462 298752 83518 298761
rect 83462 298687 83518 298696
rect 84120 260250 84148 384270
rect 86866 344720 86922 344729
rect 86866 344655 86922 344664
rect 86880 342009 86908 344655
rect 86866 342000 86922 342009
rect 86866 341935 86922 341944
rect 90362 342000 90418 342009
rect 90362 341935 90418 341944
rect 90376 332625 90404 341935
rect 90362 332616 90418 332625
rect 90362 332551 90418 332560
rect 91742 332616 91798 332625
rect 91742 332551 91798 332560
rect 91756 323649 91784 332551
rect 91742 323640 91798 323649
rect 91742 323575 91798 323584
rect 94044 312588 94096 312594
rect 94044 312530 94096 312536
rect 92388 311160 92440 311166
rect 92388 311102 92440 311108
rect 90732 309800 90784 309806
rect 90732 309742 90784 309748
rect 87420 308440 87472 308446
rect 87420 308382 87472 308388
rect 85764 307080 85816 307086
rect 85764 307022 85816 307028
rect 85776 260250 85804 307022
rect 87432 260250 87460 308382
rect 89076 271176 89128 271182
rect 89076 271118 89128 271124
rect 89088 260250 89116 271118
rect 90744 260250 90772 309742
rect 92400 260250 92428 311102
rect 94056 260250 94084 312530
rect 94148 265577 94176 390079
rect 97276 389065 97304 390102
rect 97262 389056 97318 389065
rect 97262 388991 97318 389000
rect 95700 388476 95752 388482
rect 95700 388418 95752 388424
rect 95712 386617 95740 388418
rect 95698 386608 95754 386617
rect 95698 386543 95754 386552
rect 94134 265568 94190 265577
rect 94134 265503 94190 265512
rect 95712 260250 95740 386543
rect 97276 373289 97304 388991
rect 101324 388929 101352 390116
rect 104926 390102 105676 390130
rect 101310 388920 101366 388929
rect 101310 388855 101366 388864
rect 101324 385665 101352 388855
rect 105648 386753 105676 390102
rect 108408 390102 108514 390130
rect 106188 387388 106240 387394
rect 106188 387330 106240 387336
rect 106200 387161 106228 387330
rect 108304 387320 108356 387326
rect 108304 387262 108356 387268
rect 106186 387152 106242 387161
rect 106186 387087 106242 387096
rect 105634 386744 105690 386753
rect 105634 386679 105690 386688
rect 105544 386436 105596 386442
rect 105544 386378 105596 386384
rect 101310 385656 101366 385665
rect 101310 385591 101366 385600
rect 97262 373280 97318 373289
rect 97262 373215 97318 373224
rect 97354 371920 97410 371929
rect 97354 371855 97410 371864
rect 95882 323640 95938 323649
rect 95882 323575 95938 323584
rect 95896 311953 95924 323575
rect 95882 311944 95938 311953
rect 95882 311879 95938 311888
rect 97368 260250 97396 371855
rect 99010 319288 99066 319297
rect 99010 319223 99066 319232
rect 99024 260250 99052 319223
rect 99378 311944 99434 311953
rect 99378 311879 99434 311888
rect 99392 307737 99420 311879
rect 99378 307728 99434 307737
rect 99378 307663 99434 307672
rect 102046 307728 102102 307737
rect 102046 307663 102102 307672
rect 102060 304609 102088 307663
rect 102046 304600 102102 304609
rect 102046 304535 102102 304544
rect 104806 304600 104862 304609
rect 104806 304535 104862 304544
rect 104820 300665 104848 304535
rect 104806 300656 104862 300665
rect 104806 300591 104862 300600
rect 100574 267200 100630 267209
rect 64216 259950 64552 259978
rect 65858 260222 65932 260250
rect 67514 260222 67588 260250
rect 69170 260222 69244 260250
rect 70826 260222 70900 260250
rect 72482 260222 72556 260250
rect 74138 260222 74212 260250
rect 75794 260222 75868 260250
rect 77450 260222 77524 260250
rect 79106 260222 79180 260250
rect 80762 260222 80836 260250
rect 82418 260222 82492 260250
rect 84074 260222 84148 260250
rect 85730 260222 85804 260250
rect 87386 260222 87460 260250
rect 89042 260222 89116 260250
rect 90698 260222 90772 260250
rect 92354 260222 92428 260250
rect 94010 260222 94084 260250
rect 95666 260222 95740 260250
rect 97322 260222 97396 260250
rect 98978 260222 99052 260250
rect 100496 267158 100574 267186
rect 65858 259964 65886 260222
rect 67514 259964 67542 260222
rect 69170 259964 69198 260222
rect 70826 259964 70854 260222
rect 72482 259964 72510 260222
rect 74138 259964 74166 260222
rect 75794 259964 75822 260222
rect 77450 259964 77478 260222
rect 79106 259964 79134 260222
rect 80762 259964 80790 260222
rect 82418 259964 82446 260222
rect 84074 259964 84102 260222
rect 85730 259964 85758 260222
rect 87386 259964 87414 260222
rect 89042 259964 89070 260222
rect 90698 259964 90726 260222
rect 92354 259964 92382 260222
rect 94010 259964 94038 260222
rect 95666 259964 95694 260222
rect 97322 259964 97350 260222
rect 98978 259964 99006 260222
rect 100496 259706 100524 267158
rect 100574 267135 100630 267144
rect 105556 263537 105584 386378
rect 105648 271250 105676 386679
rect 108316 386617 108344 387262
rect 108408 387025 108436 390102
rect 108394 387016 108450 387025
rect 108394 386951 108450 386960
rect 108302 386608 108358 386617
rect 108302 386543 108358 386552
rect 108408 373994 108436 386951
rect 112088 386345 112116 390116
rect 115308 390102 115690 390130
rect 119278 390102 119384 390130
rect 115308 387161 115336 390102
rect 118700 387796 118752 387802
rect 118700 387738 118752 387744
rect 115294 387152 115350 387161
rect 115294 387087 115350 387096
rect 115848 387116 115900 387122
rect 112074 386336 112130 386345
rect 112074 386271 112130 386280
rect 112442 386336 112498 386345
rect 112442 386271 112498 386280
rect 108316 373966 108436 373994
rect 108316 279478 108344 373966
rect 109682 300656 109738 300665
rect 109682 300591 109738 300600
rect 109696 295361 109724 300591
rect 109682 295352 109738 295361
rect 109682 295287 109738 295296
rect 108304 279472 108356 279478
rect 108304 279414 108356 279420
rect 112456 272649 112484 386271
rect 115308 373994 115336 387087
rect 115848 387058 115900 387064
rect 115860 386889 115888 387058
rect 115846 386880 115902 386889
rect 115846 386815 115902 386824
rect 118712 386753 118740 387738
rect 119356 387297 119384 390102
rect 122104 389904 122156 389910
rect 122104 389846 122156 389852
rect 119342 387288 119398 387297
rect 119342 387223 119398 387232
rect 118698 386744 118754 386753
rect 118698 386679 118754 386688
rect 115216 373966 115336 373994
rect 115216 297430 115244 373966
rect 119356 300150 119384 387223
rect 122116 382974 122144 389846
rect 122852 387705 122880 390116
rect 122838 387696 122894 387705
rect 122838 387631 122894 387640
rect 122104 382968 122156 382974
rect 122104 382910 122156 382916
rect 119344 300144 119396 300150
rect 119344 300086 119396 300092
rect 115204 297424 115256 297430
rect 115204 297366 115256 297372
rect 113822 295352 113878 295361
rect 113822 295287 113878 295296
rect 112442 272640 112498 272649
rect 112442 272575 112498 272584
rect 105636 271244 105688 271250
rect 105636 271186 105688 271192
rect 102138 263528 102194 263537
rect 102138 263463 102194 263472
rect 105542 263528 105598 263537
rect 105542 263463 105598 263472
rect 102152 260914 102180 263463
rect 108946 263256 109002 263265
rect 108946 263191 109002 263200
rect 105910 263120 105966 263129
rect 105910 263055 105966 263064
rect 104806 262848 104862 262857
rect 104806 262783 104862 262792
rect 104820 261089 104848 262783
rect 105924 261225 105952 263055
rect 107566 262984 107622 262993
rect 107566 262919 107622 262928
rect 105910 261216 105966 261225
rect 105910 261151 105966 261160
rect 103794 261080 103850 261089
rect 103794 261015 103850 261024
rect 104806 261080 104862 261089
rect 104806 261015 104862 261024
rect 102140 260908 102192 260914
rect 102140 260850 102192 260856
rect 102152 259978 102180 260850
rect 102152 259950 102304 259978
rect 103808 259706 103836 261015
rect 105924 259978 105952 261151
rect 107580 260953 107608 262919
rect 108960 262313 108988 263191
rect 108946 262304 109002 262313
rect 108946 262239 109002 262248
rect 107566 260944 107622 260953
rect 107566 260879 107622 260888
rect 107580 259978 107608 260879
rect 108960 260114 108988 262239
rect 105616 259950 105952 259978
rect 107272 259950 107608 259978
rect 108914 260086 108988 260114
rect 108914 259964 108942 260086
rect 100496 259678 100648 259706
rect 103808 259678 103960 259706
rect 113836 245721 113864 295287
rect 122852 282198 122880 387631
rect 126440 387569 126468 390116
rect 129752 390102 130042 390130
rect 125598 387560 125654 387569
rect 124128 387524 124180 387530
rect 125598 387495 125654 387504
rect 126426 387560 126482 387569
rect 126426 387495 126482 387504
rect 124128 387466 124180 387472
rect 124140 386889 124168 387466
rect 124126 386880 124182 386889
rect 124126 386815 124182 386824
rect 125612 301481 125640 387495
rect 129752 387433 129780 390102
rect 132500 387592 132552 387598
rect 132500 387534 132552 387540
rect 129738 387424 129794 387433
rect 129738 387359 129794 387368
rect 127624 382968 127676 382974
rect 127624 382910 127676 382916
rect 127636 378146 127664 382910
rect 127624 378140 127676 378146
rect 127624 378082 127676 378088
rect 129752 302938 129780 387359
rect 132512 384470 132540 387534
rect 133616 386481 133644 390116
rect 137204 387598 137232 390116
rect 137192 387592 137244 387598
rect 137192 387534 137244 387540
rect 140792 387258 140820 390116
rect 144380 387666 144408 390116
rect 147692 390102 147982 390130
rect 143540 387660 143592 387666
rect 143540 387602 143592 387608
rect 144368 387660 144420 387666
rect 144368 387602 144420 387608
rect 140780 387252 140832 387258
rect 140780 387194 140832 387200
rect 134522 386744 134578 386753
rect 134522 386679 134578 386688
rect 132590 386472 132646 386481
rect 132590 386407 132646 386416
rect 133602 386472 133658 386481
rect 133602 386407 133658 386416
rect 132500 384464 132552 384470
rect 132500 384406 132552 384412
rect 132604 373994 132632 386407
rect 133144 378140 133196 378146
rect 133144 378082 133196 378088
rect 132512 373966 132632 373994
rect 132512 304298 132540 373966
rect 133156 368490 133184 378082
rect 133144 368484 133196 368490
rect 133144 368426 133196 368432
rect 132500 304292 132552 304298
rect 132500 304234 132552 304240
rect 129740 302932 129792 302938
rect 129740 302874 129792 302880
rect 125598 301472 125654 301481
rect 125598 301407 125654 301416
rect 122840 282192 122892 282198
rect 122840 282134 122892 282140
rect 134536 262857 134564 386679
rect 135902 386608 135958 386617
rect 135902 386543 135958 386552
rect 135916 263129 135944 386543
rect 138664 386504 138716 386510
rect 137282 386472 137338 386481
rect 138664 386446 138716 386452
rect 137282 386407 137338 386416
rect 135902 263120 135958 263129
rect 135902 263055 135958 263064
rect 137296 262993 137324 386407
rect 138020 368484 138072 368490
rect 138020 368426 138072 368432
rect 138032 365702 138060 368426
rect 138020 365696 138072 365702
rect 138020 365638 138072 365644
rect 138676 263265 138704 386446
rect 140792 307086 140820 387194
rect 141424 365696 141476 365702
rect 141424 365638 141476 365644
rect 141436 354754 141464 365638
rect 141424 354748 141476 354754
rect 141424 354690 141476 354696
rect 143552 308446 143580 387602
rect 147692 387394 147720 390102
rect 150440 387728 150492 387734
rect 150440 387670 150492 387676
rect 150452 387433 150480 387670
rect 150438 387424 150494 387433
rect 147680 387388 147732 387394
rect 150438 387359 150494 387368
rect 147680 387330 147732 387336
rect 144184 354748 144236 354754
rect 144184 354690 144236 354696
rect 144196 343670 144224 354690
rect 144184 343664 144236 343670
rect 144184 343606 144236 343612
rect 147588 343664 147640 343670
rect 147588 343606 147640 343612
rect 147600 340882 147628 343606
rect 147588 340876 147640 340882
rect 147588 340818 147640 340824
rect 143540 308440 143592 308446
rect 143540 308382 143592 308388
rect 140780 307080 140832 307086
rect 140780 307022 140832 307028
rect 147692 271182 147720 387330
rect 151556 386889 151584 390116
rect 155144 387190 155172 390116
rect 158732 387433 158760 390116
rect 158718 387424 158774 387433
rect 158718 387359 158774 387368
rect 154580 387184 154632 387190
rect 154580 387126 154632 387132
rect 155132 387184 155184 387190
rect 155132 387126 155184 387132
rect 150438 386880 150494 386889
rect 150438 386815 150494 386824
rect 151542 386880 151598 386889
rect 151542 386815 151598 386824
rect 150452 309806 150480 386815
rect 154488 340876 154540 340882
rect 154488 340818 154540 340824
rect 154500 336734 154528 340818
rect 154488 336728 154540 336734
rect 154488 336670 154540 336676
rect 154592 311166 154620 387126
rect 158732 312594 158760 387359
rect 162320 387326 162348 390116
rect 165922 390102 166304 390130
rect 166276 388657 166304 390102
rect 169036 390102 169510 390130
rect 173098 390102 173204 390130
rect 176686 390102 177344 390130
rect 166262 388648 166318 388657
rect 166262 388583 166318 388592
rect 162308 387320 162360 387326
rect 162308 387262 162360 387268
rect 162768 387320 162820 387326
rect 162768 387262 162820 387268
rect 162780 385014 162808 387262
rect 162768 385008 162820 385014
rect 162768 384950 162820 384956
rect 166276 371929 166304 388583
rect 169036 383625 169064 390102
rect 173176 384985 173204 390102
rect 177316 386442 177344 390102
rect 180260 386753 180288 390116
rect 179418 386744 179474 386753
rect 179418 386679 179474 386688
rect 180246 386744 180302 386753
rect 180246 386679 180302 386688
rect 177304 386436 177356 386442
rect 177304 386378 177356 386384
rect 173162 384976 173218 384985
rect 173162 384911 173218 384920
rect 169022 383616 169078 383625
rect 169022 383551 169078 383560
rect 166262 371920 166318 371929
rect 166262 371855 166318 371864
rect 158812 336728 158864 336734
rect 158812 336670 158864 336676
rect 158824 332450 158852 336670
rect 158812 332444 158864 332450
rect 158812 332386 158864 332392
rect 162124 332444 162176 332450
rect 162124 332386 162176 332392
rect 162136 321638 162164 332386
rect 162124 321632 162176 321638
rect 162124 321574 162176 321580
rect 166264 321632 166316 321638
rect 166264 321574 166316 321580
rect 158720 312588 158772 312594
rect 158720 312530 158772 312536
rect 154580 311160 154632 311166
rect 154580 311102 154632 311108
rect 150440 309800 150492 309806
rect 150440 309742 150492 309748
rect 166276 292602 166304 321574
rect 169036 319433 169064 383551
rect 169022 319424 169078 319433
rect 169022 319359 169078 319368
rect 166264 292596 166316 292602
rect 166264 292538 166316 292544
rect 169024 292596 169076 292602
rect 169024 292538 169076 292544
rect 169036 279478 169064 292538
rect 169024 279472 169076 279478
rect 169024 279414 169076 279420
rect 147680 271176 147732 271182
rect 147680 271118 147732 271124
rect 173176 267073 173204 384911
rect 177316 383654 177344 386378
rect 179432 384849 179460 386679
rect 183848 386617 183876 390116
rect 186976 390102 187450 390130
rect 183834 386608 183890 386617
rect 183834 386543 183890 386552
rect 184846 386608 184902 386617
rect 184846 386543 184902 386552
rect 184860 386209 184888 386543
rect 186976 386481 187004 390102
rect 191024 386510 191052 390116
rect 191012 386504 191064 386510
rect 186962 386472 187018 386481
rect 191012 386446 191064 386452
rect 191748 386504 191800 386510
rect 191748 386446 191800 386452
rect 186962 386407 187018 386416
rect 184846 386200 184902 386209
rect 184846 386135 184902 386144
rect 179418 384840 179474 384849
rect 179418 384775 179474 384784
rect 177304 383648 177356 383654
rect 177304 383590 177356 383596
rect 186976 383489 187004 386407
rect 191760 384946 191788 386446
rect 191748 384940 191800 384946
rect 191748 384882 191800 384888
rect 186962 383480 187018 383489
rect 186962 383415 187018 383424
rect 182824 279472 182876 279478
rect 182824 279414 182876 279420
rect 173162 267064 173218 267073
rect 173162 266999 173218 267008
rect 138662 263256 138718 263265
rect 138662 263191 138718 263200
rect 137282 262984 137338 262993
rect 137282 262919 137338 262928
rect 134522 262848 134578 262857
rect 134522 262783 134578 262792
rect 117962 257952 118018 257961
rect 117962 257887 118018 257896
rect 116398 252512 116454 252521
rect 116398 252447 116454 252456
rect 113822 245712 113878 245721
rect 113822 245647 113878 245656
rect 114650 245712 114706 245721
rect 114650 245647 114706 245656
rect 114664 240145 114692 245647
rect 114650 240136 114706 240145
rect 114650 240071 114706 240080
rect 48226 215112 48282 215121
rect 48226 215047 48282 215056
rect 48240 200122 48268 215047
rect 111064 214600 111116 214606
rect 111064 214542 111116 214548
rect 48228 200116 48280 200122
rect 48228 200058 48280 200064
rect 50954 199866 50982 200124
rect 52624 200110 52960 200138
rect 54280 200110 54616 200138
rect 55936 200110 56272 200138
rect 57592 200110 57928 200138
rect 50954 199838 51028 199866
rect 51000 198529 51028 199838
rect 50986 198520 51042 198529
rect 50986 198455 51042 198464
rect 52932 197441 52960 200110
rect 54588 197713 54616 200110
rect 56244 197849 56272 200110
rect 57900 198257 57928 200110
rect 59234 199866 59262 200124
rect 60904 200110 61056 200138
rect 62560 200110 62712 200138
rect 64216 200110 64552 200138
rect 59234 199838 59308 199866
rect 57886 198248 57942 198257
rect 57886 198183 57942 198192
rect 56230 197840 56286 197849
rect 56230 197775 56286 197784
rect 54574 197704 54630 197713
rect 54574 197639 54630 197648
rect 52918 197432 52974 197441
rect 52918 197367 52974 197376
rect 59280 140321 59308 199838
rect 61028 180794 61056 200110
rect 62684 180794 62712 200110
rect 64524 198393 64552 200110
rect 65858 199866 65886 200124
rect 67514 199866 67542 200124
rect 69184 200110 69520 200138
rect 70840 200110 71176 200138
rect 72496 200110 72832 200138
rect 74152 200110 74488 200138
rect 75808 200110 75960 200138
rect 77464 200110 77800 200138
rect 79120 200110 79456 200138
rect 80776 200110 81112 200138
rect 82432 200110 82768 200138
rect 65858 199838 65932 199866
rect 67514 199838 67588 199866
rect 64510 198384 64566 198393
rect 64510 198319 64566 198328
rect 60936 180766 61056 180794
rect 62592 180766 62712 180794
rect 59266 140312 59322 140321
rect 59266 140247 59322 140256
rect 60936 138825 60964 180766
rect 62592 138961 62620 180766
rect 62578 138952 62634 138961
rect 62578 138887 62634 138896
rect 60922 138816 60978 138825
rect 60922 138751 60978 138760
rect 65904 138009 65932 199838
rect 67560 197305 67588 199838
rect 69492 197985 69520 200110
rect 70398 198520 70454 198529
rect 70398 198455 70454 198464
rect 69478 197976 69534 197985
rect 69478 197911 69534 197920
rect 70412 197538 70440 198455
rect 71148 197577 71176 200110
rect 72804 198121 72832 200110
rect 72790 198112 72846 198121
rect 72790 198047 72846 198056
rect 71778 197840 71834 197849
rect 71778 197775 71834 197784
rect 71134 197568 71190 197577
rect 70400 197532 70452 197538
rect 71134 197503 71190 197512
rect 70400 197474 70452 197480
rect 71792 197402 71820 197775
rect 74460 197713 74488 200110
rect 75932 200025 75960 200110
rect 75918 200016 75974 200025
rect 75918 199951 75974 199960
rect 77772 198665 77800 200110
rect 77758 198656 77814 198665
rect 77758 198591 77814 198600
rect 79322 198248 79378 198257
rect 79322 198183 79378 198192
rect 73158 197704 73214 197713
rect 73158 197639 73214 197648
rect 74446 197704 74502 197713
rect 74446 197639 74502 197648
rect 78588 197668 78640 197674
rect 73172 197470 73200 197639
rect 78588 197610 78640 197616
rect 73160 197464 73212 197470
rect 78600 197441 78628 197610
rect 79336 197606 79364 198183
rect 79324 197600 79376 197606
rect 79324 197542 79376 197548
rect 79428 197441 79456 200110
rect 81084 198937 81112 200110
rect 82740 199753 82768 200110
rect 84074 199866 84102 200124
rect 85744 200110 86080 200138
rect 87400 200110 87736 200138
rect 89056 200110 89392 200138
rect 90712 200110 91048 200138
rect 84074 199838 84148 199866
rect 82726 199744 82782 199753
rect 82726 199679 82782 199688
rect 84120 199345 84148 199838
rect 84106 199336 84162 199345
rect 84106 199271 84162 199280
rect 81070 198928 81126 198937
rect 81070 198863 81126 198872
rect 85578 198384 85634 198393
rect 85578 198319 85634 198328
rect 85592 197742 85620 198319
rect 86052 198257 86080 200110
rect 86960 198620 87012 198626
rect 86960 198562 87012 198568
rect 86038 198248 86094 198257
rect 86038 198183 86094 198192
rect 85580 197736 85632 197742
rect 85580 197678 85632 197684
rect 86972 197577 87000 198562
rect 87708 198529 87736 200110
rect 88340 198688 88392 198694
rect 88340 198630 88392 198636
rect 87694 198520 87750 198529
rect 87694 198455 87750 198464
rect 88352 197985 88380 198630
rect 89364 198393 89392 200110
rect 91020 198801 91048 200110
rect 92354 199866 92382 200124
rect 94024 200110 94360 200138
rect 95680 200110 96016 200138
rect 97336 200110 97672 200138
rect 98992 200110 99236 200138
rect 92354 199838 92428 199866
rect 92400 199481 92428 199838
rect 92386 199472 92442 199481
rect 92386 199407 92442 199416
rect 94332 199073 94360 200110
rect 95988 200025 96016 200110
rect 94502 200016 94558 200025
rect 94502 199951 94558 199960
rect 95974 200016 96030 200025
rect 95974 199951 96030 199960
rect 94516 199646 94544 199951
rect 95240 199844 95292 199850
rect 95240 199786 95292 199792
rect 94504 199640 94556 199646
rect 94504 199582 94556 199588
rect 95252 199345 95280 199786
rect 95238 199336 95294 199345
rect 95238 199271 95294 199280
rect 94318 199064 94374 199073
rect 94318 198999 94374 199008
rect 91006 198792 91062 198801
rect 91006 198727 91062 198736
rect 96620 198484 96672 198490
rect 96620 198426 96672 198432
rect 89350 198384 89406 198393
rect 89350 198319 89406 198328
rect 88338 197976 88394 197985
rect 88338 197911 88394 197920
rect 96632 197713 96660 198426
rect 96618 197704 96674 197713
rect 96618 197639 96674 197648
rect 97644 197577 97672 200110
rect 98000 198552 98052 198558
rect 98000 198494 98052 198500
rect 98012 198121 98040 198494
rect 97998 198112 98054 198121
rect 97998 198047 98054 198056
rect 99208 197985 99236 200110
rect 100634 199889 100662 200124
rect 102304 200110 102640 200138
rect 103960 200110 104296 200138
rect 105616 200110 105952 200138
rect 107272 200110 107608 200138
rect 100620 199880 100676 199889
rect 100620 199815 100676 199824
rect 100668 199776 100720 199782
rect 100666 199744 100668 199753
rect 102612 199753 102640 200110
rect 100720 199744 100722 199753
rect 100666 199679 100722 199688
rect 102598 199744 102654 199753
rect 102598 199679 102654 199688
rect 103428 199708 103480 199714
rect 103428 199650 103480 199656
rect 103440 198937 103468 199650
rect 103426 198928 103482 198937
rect 103426 198863 103482 198872
rect 104164 198416 104216 198422
rect 104164 198358 104216 198364
rect 99194 197976 99250 197985
rect 99194 197911 99250 197920
rect 86958 197568 87014 197577
rect 86958 197503 87014 197512
rect 97630 197568 97686 197577
rect 97630 197503 97686 197512
rect 104176 197441 104204 198358
rect 104268 197849 104296 200110
rect 104900 199980 104952 199986
rect 104900 199922 104952 199928
rect 104912 199481 104940 199922
rect 105924 199617 105952 200110
rect 106280 199912 106332 199918
rect 106280 199854 106332 199860
rect 105910 199608 105966 199617
rect 105910 199543 105966 199552
rect 104898 199472 104954 199481
rect 104898 199407 104954 199416
rect 106292 198801 106320 199854
rect 107580 199481 107608 200110
rect 107658 200016 107714 200025
rect 107658 199951 107714 199960
rect 107672 199578 107700 199951
rect 108914 199866 108942 200124
rect 111076 200122 111104 214542
rect 110420 200116 110472 200122
rect 110420 200058 110472 200064
rect 111064 200116 111116 200122
rect 111064 200058 111116 200064
rect 108914 199838 108988 199866
rect 107660 199572 107712 199578
rect 107660 199514 107712 199520
rect 107566 199472 107622 199481
rect 107566 199407 107622 199416
rect 108960 199345 108988 199838
rect 108946 199336 109002 199345
rect 108946 199271 109002 199280
rect 106278 198792 106334 198801
rect 106278 198727 106334 198736
rect 104254 197840 104310 197849
rect 104254 197775 104310 197784
rect 73160 197406 73212 197412
rect 78586 197432 78642 197441
rect 71780 197396 71832 197402
rect 78586 197367 78642 197376
rect 79414 197432 79470 197441
rect 79414 197367 79470 197376
rect 104162 197432 104218 197441
rect 104162 197367 104218 197376
rect 71780 197338 71832 197344
rect 67546 197296 67602 197305
rect 67546 197231 67602 197240
rect 95146 195256 95202 195265
rect 95146 195191 95202 195200
rect 65890 138000 65946 138009
rect 65890 137935 65946 137944
rect 66168 137896 66220 137902
rect 66168 137838 66220 137844
rect 66180 137601 66208 137838
rect 66166 137592 66222 137601
rect 66166 137527 66222 137536
rect 89166 130384 89222 130393
rect 89166 130319 89222 130328
rect 85670 129024 85726 129033
rect 85670 128959 85726 128968
rect 47582 110664 47638 110673
rect 47582 110599 47638 110608
rect 46662 97200 46718 97209
rect 46662 97135 46718 97144
rect 46676 480 46704 97135
rect 65614 87952 65670 87961
rect 65536 87910 65614 87938
rect 52918 87816 52974 87825
rect 52918 87751 52974 87760
rect 50986 85776 51042 85785
rect 50908 85734 50986 85762
rect 50908 84810 50936 85734
rect 50986 85711 51042 85720
rect 52932 84946 52960 87751
rect 60646 87680 60702 87689
rect 60646 87615 60702 87624
rect 57610 87408 57666 87417
rect 57610 87343 57666 87352
rect 54666 87136 54722 87145
rect 54588 87094 54666 87122
rect 54588 84946 54616 87094
rect 54666 87071 54722 87080
rect 56506 86184 56562 86193
rect 56152 86142 56506 86170
rect 56152 84946 56180 86142
rect 56506 86119 56562 86128
rect 57624 84946 57652 87343
rect 59266 87272 59322 87281
rect 59266 87207 59322 87216
rect 59280 84946 59308 87207
rect 60660 84946 60688 87615
rect 62026 87544 62082 87553
rect 62026 87479 62082 87488
rect 62040 85082 62068 87479
rect 63866 85640 63922 85649
rect 63866 85575 63922 85584
rect 52624 84918 52960 84946
rect 54188 84918 54616 84946
rect 55752 84918 56180 84946
rect 57316 84918 57652 84946
rect 58880 84918 59308 84946
rect 60444 84918 60688 84946
rect 61994 85054 62068 85082
rect 61994 84932 62022 85054
rect 63880 84946 63908 85575
rect 65536 84946 65564 87910
rect 65614 87887 65670 87896
rect 84842 87680 84898 87689
rect 84842 87615 84898 87624
rect 73068 87372 73120 87378
rect 73068 87314 73120 87320
rect 66996 87236 67048 87242
rect 66996 87178 67048 87184
rect 67008 84946 67036 87178
rect 70124 87168 70176 87174
rect 70124 87110 70176 87116
rect 68650 85912 68706 85921
rect 68650 85847 68706 85856
rect 68664 84946 68692 85847
rect 70136 84946 70164 87110
rect 73080 84946 73108 87314
rect 74448 87304 74500 87310
rect 74448 87246 74500 87252
rect 74460 85082 74488 87246
rect 76472 87100 76524 87106
rect 76472 87042 76524 87048
rect 63572 84918 63908 84946
rect 65136 84918 65564 84946
rect 66700 84918 67036 84946
rect 68264 84918 68692 84946
rect 69828 84918 70164 84946
rect 72956 84918 73108 84946
rect 74368 85054 74488 85082
rect 74368 84810 74396 85054
rect 76484 84946 76512 87042
rect 82728 87032 82780 87038
rect 82728 86974 82780 86980
rect 76084 84918 76512 84946
rect 80748 84960 80804 84969
rect 82740 84946 82768 86974
rect 82340 84918 82768 84946
rect 80748 84895 80804 84904
rect 77620 84824 77676 84833
rect 50908 84782 51060 84810
rect 74368 84782 74520 84810
rect 77620 84759 77676 84768
rect 71364 84688 71420 84697
rect 71364 84623 71420 84632
rect 79184 84552 79240 84561
rect 83904 84510 84240 84538
rect 79184 84487 79240 84496
rect 84212 82822 84240 84510
rect 84200 82816 84252 82822
rect 84200 82758 84252 82764
rect 48226 81696 48282 81705
rect 48226 81631 48282 81640
rect 47858 80336 47914 80345
rect 47858 80271 47914 80280
rect 47490 64016 47546 64025
rect 47490 63951 47546 63960
rect 47504 15881 47532 63951
rect 47582 61296 47638 61305
rect 47582 61231 47638 61240
rect 47596 21321 47624 61231
rect 47766 58576 47822 58585
rect 47766 58511 47822 58520
rect 47674 57216 47730 57225
rect 47674 57151 47730 57160
rect 47688 28257 47716 57151
rect 47674 28248 47730 28257
rect 47674 28183 47730 28192
rect 47780 26897 47808 58511
rect 47872 46345 47900 80271
rect 48134 65376 48190 65385
rect 48134 65311 48190 65320
rect 48042 62656 48098 62665
rect 48042 62591 48098 62600
rect 47950 59936 48006 59945
rect 47950 59871 48006 59880
rect 47858 46336 47914 46345
rect 47858 46271 47914 46280
rect 47766 26888 47822 26897
rect 47766 26823 47822 26832
rect 47964 25537 47992 59871
rect 47950 25528 48006 25537
rect 47950 25463 48006 25472
rect 48056 22681 48084 62591
rect 48148 43625 48176 65311
rect 48240 49065 48268 81631
rect 84856 79393 84884 87615
rect 85026 87408 85082 87417
rect 85026 87343 85082 87352
rect 84936 87236 84988 87242
rect 84936 87178 84988 87184
rect 84948 83502 84976 87178
rect 84936 83496 84988 83502
rect 84936 83438 84988 83444
rect 85040 80753 85068 87343
rect 85026 80744 85082 80753
rect 85026 80679 85082 80688
rect 84842 79384 84898 79393
rect 84842 79319 84898 79328
rect 49422 78976 49478 78985
rect 49422 78911 49478 78920
rect 49330 77616 49386 77625
rect 49330 77551 49386 77560
rect 49238 69456 49294 69465
rect 49238 69391 49294 69400
rect 49146 68096 49202 68105
rect 49146 68031 49202 68040
rect 49054 55856 49110 55865
rect 49054 55791 49110 55800
rect 48226 49056 48282 49065
rect 48226 48991 48282 49000
rect 48134 43616 48190 43625
rect 48134 43551 48190 43560
rect 48962 28520 49018 28529
rect 48962 28455 49018 28464
rect 48042 22672 48098 22681
rect 48042 22607 48098 22616
rect 47582 21312 47638 21321
rect 47582 21247 47638 21256
rect 47490 15872 47546 15881
rect 47490 15807 47546 15816
rect 47858 6352 47914 6361
rect 47858 6287 47914 6296
rect 47872 480 47900 6287
rect 48976 480 49004 28455
rect 49068 24177 49096 55791
rect 49160 39273 49188 68031
rect 49146 39264 49202 39273
rect 49146 39199 49202 39208
rect 49252 37913 49280 69391
rect 49344 48929 49372 77551
rect 49330 48920 49386 48929
rect 49330 48855 49386 48864
rect 49436 44849 49464 78911
rect 50434 75984 50490 75993
rect 50434 75919 50490 75928
rect 49606 74896 49662 74905
rect 49606 74831 49662 74840
rect 49514 72176 49570 72185
rect 49514 72111 49570 72120
rect 49422 44840 49478 44849
rect 49422 44775 49478 44784
rect 49238 37904 49294 37913
rect 49238 37839 49294 37848
rect 49528 36553 49556 72111
rect 49514 36544 49570 36553
rect 49514 36479 49570 36488
rect 49620 33833 49648 74831
rect 50158 70408 50214 70417
rect 50158 70343 50214 70352
rect 50066 52592 50122 52601
rect 50066 52527 50122 52536
rect 50080 42265 50108 52527
rect 50066 42256 50122 42265
rect 50066 42191 50122 42200
rect 49606 33824 49662 33833
rect 49606 33759 49662 33768
rect 49054 24168 49110 24177
rect 49054 24103 49110 24112
rect 50172 18601 50200 70343
rect 50250 66328 50306 66337
rect 50250 66263 50306 66272
rect 50158 18592 50214 18601
rect 50158 18527 50214 18536
rect 50264 17241 50292 66263
rect 50342 49192 50398 49201
rect 50342 49127 50398 49136
rect 50250 17232 50306 17241
rect 50250 17167 50306 17176
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 354 50242 480
rect 50356 354 50384 49127
rect 50448 30977 50476 75919
rect 50526 73264 50582 73273
rect 50526 73199 50582 73208
rect 50540 35193 50568 73199
rect 50618 53952 50674 53961
rect 50618 53887 50674 53896
rect 50526 35184 50582 35193
rect 50526 35119 50582 35128
rect 50434 30968 50490 30977
rect 50434 30903 50490 30912
rect 50632 29617 50660 53887
rect 84658 53272 84714 53281
rect 84658 53207 84714 53216
rect 67914 50280 67970 50289
rect 67914 50215 67970 50224
rect 50876 50102 51028 50130
rect 52256 50102 52408 50130
rect 53636 50102 53788 50130
rect 51000 47841 51028 50102
rect 50986 47832 51042 47841
rect 50986 47767 51042 47776
rect 52380 47705 52408 50102
rect 52366 47696 52422 47705
rect 52366 47631 52422 47640
rect 53760 47569 53788 50102
rect 55002 49858 55030 50116
rect 56396 50102 56548 50130
rect 55002 49830 55076 49858
rect 53746 47560 53802 47569
rect 53746 47495 53802 47504
rect 51354 38176 51410 38185
rect 51354 38111 51410 38120
rect 50618 29608 50674 29617
rect 50618 29543 50674 29552
rect 51368 480 51396 38111
rect 52550 29880 52606 29889
rect 52550 29815 52606 29824
rect 52564 480 52592 29815
rect 54942 21584 54998 21593
rect 54942 21519 54998 21528
rect 53746 2816 53802 2825
rect 53746 2751 53802 2760
rect 53760 480 53788 2751
rect 54956 480 54984 21519
rect 55048 9081 55076 49830
rect 56520 46209 56548 50102
rect 57762 49858 57790 50116
rect 59142 49858 59170 50116
rect 60536 50102 60688 50130
rect 57762 49830 57836 49858
rect 59142 49830 59216 49858
rect 56506 46200 56562 46209
rect 56506 46135 56562 46144
rect 56046 31240 56102 31249
rect 56046 31175 56102 31184
rect 55034 9072 55090 9081
rect 55034 9007 55090 9016
rect 56060 480 56088 31175
rect 57242 14784 57298 14793
rect 57242 14719 57298 14728
rect 57256 480 57284 14719
rect 57808 8945 57836 49830
rect 58438 25664 58494 25673
rect 58438 25599 58494 25608
rect 57794 8936 57850 8945
rect 57794 8871 57850 8880
rect 58452 480 58480 25599
rect 59188 10305 59216 49830
rect 60660 47977 60688 50102
rect 61902 49858 61930 50116
rect 63282 49858 63310 50116
rect 64676 50102 64828 50130
rect 61902 49830 61976 49858
rect 63282 49830 63356 49858
rect 60646 47968 60702 47977
rect 60646 47903 60702 47912
rect 60830 44976 60886 44985
rect 60830 44911 60886 44920
rect 59634 32736 59690 32745
rect 59634 32671 59690 32680
rect 59174 10296 59230 10305
rect 59174 10231 59230 10240
rect 59648 480 59676 32671
rect 60844 480 60872 44911
rect 61948 13025 61976 49830
rect 62762 47968 62818 47977
rect 62762 47903 62818 47912
rect 62026 22808 62082 22817
rect 62026 22743 62082 22752
rect 61934 13016 61990 13025
rect 61934 12951 61990 12960
rect 62040 480 62068 22743
rect 62776 11665 62804 47903
rect 63328 43489 63356 49830
rect 64800 47025 64828 50102
rect 66042 49858 66070 50116
rect 67422 49858 67450 50116
rect 66042 49830 66116 49858
rect 67422 49830 67496 49858
rect 64786 47016 64842 47025
rect 64786 46951 64842 46960
rect 65614 47016 65670 47025
rect 65614 46951 65670 46960
rect 63314 43480 63370 43489
rect 63314 43415 63370 43424
rect 65522 36680 65578 36689
rect 65522 36615 65578 36624
rect 63222 28384 63278 28393
rect 63222 28319 63278 28328
rect 62762 11656 62818 11665
rect 62762 11591 62818 11600
rect 63236 480 63264 28319
rect 64326 3496 64382 3505
rect 64326 3431 64382 3440
rect 64340 480 64368 3431
rect 65536 480 65564 36615
rect 65628 19961 65656 46951
rect 66088 42129 66116 49830
rect 66074 42120 66130 42129
rect 66074 42055 66130 42064
rect 65614 19952 65670 19961
rect 65614 19887 65670 19896
rect 67468 14521 67496 49830
rect 67454 14512 67510 14521
rect 67454 14447 67510 14456
rect 66718 10432 66774 10441
rect 66718 10367 66774 10376
rect 66732 480 66760 10367
rect 67928 480 67956 50215
rect 68802 49858 68830 50116
rect 70182 49858 70210 50116
rect 71576 50102 71728 50130
rect 68802 49830 68876 49858
rect 70182 49830 70256 49858
rect 68848 40633 68876 49830
rect 68834 40624 68890 40633
rect 68834 40559 68890 40568
rect 69110 33960 69166 33969
rect 69110 33895 69166 33904
rect 69124 480 69152 33895
rect 70228 32473 70256 49830
rect 71502 49328 71558 49337
rect 71502 49263 71558 49272
rect 70214 32464 70270 32473
rect 70214 32399 70270 32408
rect 70306 31104 70362 31113
rect 70306 31039 70362 31048
rect 70320 480 70348 31039
rect 71516 480 71544 49263
rect 71700 47818 71728 50102
rect 72942 49858 72970 50116
rect 74336 50102 74488 50130
rect 75716 50102 75868 50130
rect 77096 50102 77248 50130
rect 78476 50102 78628 50130
rect 79856 50102 80008 50130
rect 72942 49830 73016 49858
rect 71700 47790 72464 47818
rect 72436 11801 72464 47790
rect 72988 13161 73016 49830
rect 74460 47025 74488 50102
rect 75840 47818 75868 50102
rect 77220 48113 77248 50102
rect 77206 48104 77262 48113
rect 77206 48039 77262 48048
rect 78600 47977 78628 50102
rect 79322 48104 79378 48113
rect 79322 48039 79378 48048
rect 78586 47968 78642 47977
rect 78586 47903 78642 47912
rect 75840 47790 76604 47818
rect 74446 47016 74502 47025
rect 74446 46951 74502 46960
rect 75182 47016 75238 47025
rect 75182 46951 75238 46960
rect 74998 38040 75054 38049
rect 74998 37975 75054 37984
rect 72974 13152 73030 13161
rect 72974 13087 73030 13096
rect 72422 11792 72478 11801
rect 72422 11727 72478 11736
rect 73802 7848 73858 7857
rect 73802 7783 73858 7792
rect 72606 6488 72662 6497
rect 72606 6423 72662 6432
rect 72620 480 72648 6423
rect 73816 480 73844 7783
rect 75012 480 75040 37975
rect 75196 20097 75224 46951
rect 75182 20088 75238 20097
rect 75182 20023 75238 20032
rect 76576 14657 76604 47790
rect 78586 21448 78642 21457
rect 78586 21383 78642 21392
rect 76562 14648 76618 14657
rect 76562 14583 76618 14592
rect 76194 6624 76250 6633
rect 76194 6559 76250 6568
rect 76208 480 76236 6559
rect 77390 5128 77446 5137
rect 77390 5063 77446 5072
rect 77404 480 77432 5063
rect 78600 480 78628 21383
rect 79336 16017 79364 48039
rect 79506 47968 79562 47977
rect 79506 47903 79562 47912
rect 79520 24313 79548 47903
rect 79980 47818 80008 50102
rect 81222 49858 81250 50116
rect 82616 50102 82768 50130
rect 83996 50102 84148 50130
rect 81222 49830 81296 49858
rect 79980 47790 80744 47818
rect 79506 24304 79562 24313
rect 79506 24239 79562 24248
rect 80716 17377 80744 47790
rect 81268 40769 81296 49830
rect 82740 47818 82768 50102
rect 84120 47977 84148 50102
rect 84106 47968 84162 47977
rect 84106 47903 84162 47912
rect 82740 47790 83044 47818
rect 81254 40760 81310 40769
rect 81254 40695 81310 40704
rect 83016 39409 83044 47790
rect 83002 39400 83058 39409
rect 83002 39335 83058 39344
rect 83278 35320 83334 35329
rect 83278 35255 83334 35264
rect 82082 32600 82138 32609
rect 82082 32535 82138 32544
rect 80886 29744 80942 29753
rect 80886 29679 80942 29688
rect 80702 17368 80758 17377
rect 80702 17303 80758 17312
rect 79322 16008 79378 16017
rect 79322 15943 79378 15952
rect 79690 6760 79746 6769
rect 79690 6695 79746 6704
rect 79704 480 79732 6695
rect 80900 480 80928 29679
rect 82096 480 82124 32535
rect 83292 480 83320 35255
rect 84672 6914 84700 53207
rect 84488 6886 84700 6914
rect 84488 480 84516 6886
rect 85684 480 85712 128959
rect 86866 93120 86922 93129
rect 86866 93055 86922 93064
rect 86222 87816 86278 87825
rect 86222 87751 86278 87760
rect 86236 51921 86264 87751
rect 86316 87304 86368 87310
rect 86316 87246 86368 87252
rect 86328 69698 86356 87246
rect 86316 69692 86368 69698
rect 86316 69634 86368 69640
rect 86222 51912 86278 51921
rect 86222 51847 86278 51856
rect 86880 480 86908 93055
rect 87694 90536 87750 90545
rect 87694 90471 87750 90480
rect 87602 87136 87658 87145
rect 87602 87071 87658 87080
rect 87050 52592 87106 52601
rect 87050 52527 87106 52536
rect 86958 51776 87014 51785
rect 86958 51711 87014 51720
rect 86972 40730 87000 51711
rect 86960 40724 87012 40730
rect 86960 40666 87012 40672
rect 87064 32881 87092 52527
rect 87050 32872 87106 32881
rect 87050 32807 87106 32816
rect 87616 5001 87644 87071
rect 87708 52601 87736 90471
rect 87786 87544 87842 87553
rect 87786 87479 87842 87488
rect 87800 54641 87828 87479
rect 87786 54632 87842 54641
rect 87786 54567 87842 54576
rect 87694 52592 87750 52601
rect 87694 52527 87750 52536
rect 88246 51776 88302 51785
rect 88246 51711 88248 51720
rect 88300 51711 88302 51720
rect 88248 51682 88300 51688
rect 87694 47968 87750 47977
rect 87694 47903 87750 47912
rect 87708 18737 87736 47903
rect 87694 18728 87750 18737
rect 87694 18663 87750 18672
rect 87970 9208 88026 9217
rect 87970 9143 88026 9152
rect 87602 4992 87658 5001
rect 87602 4927 87658 4936
rect 87984 480 88012 9143
rect 89180 480 89208 130319
rect 92754 124808 92810 124817
rect 92754 124743 92810 124752
rect 91558 123584 91614 123593
rect 91558 123519 91614 123528
rect 90362 108352 90418 108361
rect 90362 108287 90418 108296
rect 90376 480 90404 108287
rect 90456 87032 90508 87038
rect 90456 86974 90508 86980
rect 90468 50386 90496 86974
rect 90456 50380 90508 50386
rect 90456 50322 90508 50328
rect 91572 480 91600 123519
rect 91742 87952 91798 87961
rect 91742 87887 91798 87896
rect 91756 7585 91784 87887
rect 91926 87272 91982 87281
rect 91926 87207 91982 87216
rect 91940 53145 91968 87207
rect 91926 53136 91982 53145
rect 91926 53071 91982 53080
rect 91742 7576 91798 7585
rect 91742 7511 91798 7520
rect 92768 480 92796 124743
rect 93950 118008 94006 118017
rect 93950 117943 94006 117952
rect 93964 480 93992 117943
rect 95160 480 95188 195191
rect 105726 141400 105782 141409
rect 105726 141335 105782 141344
rect 101402 133240 101458 133249
rect 101402 133175 101458 133184
rect 98642 120864 98698 120873
rect 98642 120799 98698 120808
rect 96250 119368 96306 119377
rect 96250 119303 96306 119312
rect 96264 480 96292 119303
rect 97446 106856 97502 106865
rect 97446 106791 97502 106800
rect 97460 480 97488 106791
rect 98656 480 98684 120799
rect 99838 102776 99894 102785
rect 99838 102711 99894 102720
rect 98736 87168 98788 87174
rect 98736 87110 98788 87116
rect 98748 10334 98776 87110
rect 98736 10328 98788 10334
rect 98736 10270 98788 10276
rect 99852 480 99880 102711
rect 101034 94480 101090 94489
rect 101034 94415 101090 94424
rect 101048 480 101076 94415
rect 101416 3505 101444 133175
rect 103334 131744 103390 131753
rect 103334 131679 103390 131688
rect 102230 101552 102286 101561
rect 102230 101487 102286 101496
rect 101402 3496 101458 3505
rect 101402 3431 101458 3440
rect 102244 480 102272 101487
rect 103348 480 103376 131679
rect 104530 105496 104586 105505
rect 104530 105431 104586 105440
rect 104544 480 104572 105431
rect 105542 80336 105598 80345
rect 105542 80271 105598 80280
rect 105556 51785 105584 80271
rect 105542 51776 105598 51785
rect 105542 51711 105598 51720
rect 105740 480 105768 141335
rect 106922 98832 106978 98841
rect 106922 98767 106978 98776
rect 106936 480 106964 98767
rect 108118 95840 108174 95849
rect 108118 95775 108174 95784
rect 108132 480 108160 95775
rect 110432 51746 110460 200058
rect 112810 192536 112866 192545
rect 112810 192471 112866 192480
rect 110510 108488 110566 108497
rect 110510 108423 110566 108432
rect 110420 51740 110472 51746
rect 110420 51682 110472 51688
rect 109314 3496 109370 3505
rect 109314 3431 109370 3440
rect 109328 480 109356 3431
rect 110524 480 110552 108423
rect 111614 97336 111670 97345
rect 111614 97271 111670 97280
rect 111628 480 111656 97271
rect 112824 480 112852 192471
rect 115846 137864 115902 137873
rect 115846 137799 115848 137808
rect 115900 137799 115902 137808
rect 115848 137770 115900 137776
rect 115202 137456 115258 137465
rect 115202 137391 115258 137400
rect 114006 123448 114062 123457
rect 114006 123383 114062 123392
rect 114020 480 114048 123383
rect 115216 480 115244 137391
rect 116412 480 116440 252447
rect 116582 240136 116638 240145
rect 116582 240071 116638 240080
rect 116596 224233 116624 240071
rect 116582 224224 116638 224233
rect 116582 224159 116638 224168
rect 117976 3369 118004 257887
rect 178682 256864 178738 256873
rect 178682 256799 178738 256808
rect 123482 254688 123538 254697
rect 123482 254623 123538 254632
rect 120722 224224 120778 224233
rect 120722 224159 120778 224168
rect 120736 213874 120764 224159
rect 120736 213846 121500 213874
rect 121472 211177 121500 213846
rect 121458 211168 121514 211177
rect 121458 211103 121514 211112
rect 118700 137760 118752 137766
rect 118700 137702 118752 137708
rect 118712 137193 118740 137702
rect 118790 137592 118846 137601
rect 118790 137527 118846 137536
rect 118698 137184 118754 137193
rect 118698 137119 118754 137128
rect 117962 3360 118018 3369
rect 117962 3295 118018 3304
rect 117594 2952 117650 2961
rect 117594 2887 117650 2896
rect 117608 480 117636 2887
rect 118804 480 118832 137527
rect 122286 104272 122342 104281
rect 122286 104207 122342 104216
rect 119894 102912 119950 102921
rect 119894 102847 119950 102856
rect 119908 480 119936 102847
rect 121090 90400 121146 90409
rect 121090 90335 121146 90344
rect 121104 480 121132 90335
rect 122300 480 122328 104207
rect 123496 480 123524 254623
rect 163502 250336 163558 250345
rect 163502 250271 163558 250280
rect 126242 243808 126298 243817
rect 126242 243743 126298 243752
rect 123574 211168 123630 211177
rect 123574 211103 123630 211112
rect 123588 200705 123616 211103
rect 123574 200696 123630 200705
rect 123574 200631 123630 200640
rect 124678 100192 124734 100201
rect 124678 100127 124734 100136
rect 124692 480 124720 100127
rect 126256 9217 126284 243743
rect 142802 240544 142858 240553
rect 142802 240479 142858 240488
rect 140042 237280 140098 237289
rect 140042 237215 140098 237224
rect 138662 231840 138718 231849
rect 138662 231775 138718 231784
rect 126978 134600 127034 134609
rect 126978 134535 127034 134544
rect 126242 9208 126298 9217
rect 126242 9143 126298 9152
rect 126992 480 127020 134535
rect 130566 127800 130622 127809
rect 130566 127735 130622 127744
rect 130580 480 130608 127735
rect 134154 119504 134210 119513
rect 134154 119439 134210 119448
rect 134168 480 134196 119439
rect 137650 118144 137706 118153
rect 137650 118079 137706 118088
rect 137664 480 137692 118079
rect 138676 28529 138704 231775
rect 138662 28520 138718 28529
rect 138662 28455 138718 28464
rect 140056 10441 140084 237215
rect 141238 130520 141294 130529
rect 141238 130455 141294 130464
rect 140042 10432 140098 10441
rect 140042 10367 140098 10376
rect 141252 480 141280 130455
rect 142816 5137 142844 240479
rect 151082 239456 151138 239465
rect 151082 239391 151138 239400
rect 146942 234016 146998 234025
rect 146942 233951 146998 233960
rect 144182 228576 144238 228585
rect 144182 228511 144238 228520
rect 144196 113801 144224 228511
rect 144734 138272 144790 138281
rect 144734 138207 144790 138216
rect 144182 113792 144238 113801
rect 144182 113727 144238 113736
rect 142802 5128 142858 5137
rect 142802 5063 142858 5072
rect 144748 480 144776 138207
rect 146956 31249 146984 233951
rect 148322 116648 148378 116657
rect 148322 116583 148378 116592
rect 146942 31240 146998 31249
rect 146942 31175 146998 31184
rect 148336 480 148364 116583
rect 151096 7857 151124 239391
rect 152462 229664 152518 229673
rect 152462 229599 152518 229608
rect 151818 129160 151874 129169
rect 151818 129095 151874 129104
rect 151082 7848 151138 7857
rect 151082 7783 151138 7792
rect 151832 480 151860 129095
rect 152476 111081 152504 229599
rect 155222 227488 155278 227497
rect 155222 227423 155278 227432
rect 152462 111072 152518 111081
rect 152462 111007 152518 111016
rect 155236 109721 155264 227423
rect 158718 218784 158774 218793
rect 158718 218719 158774 218728
rect 158732 214606 158760 218719
rect 158720 214600 158772 214606
rect 158720 214542 158772 214548
rect 162490 136096 162546 136105
rect 162490 136031 162546 136040
rect 155406 111072 155462 111081
rect 155406 111007 155462 111016
rect 155222 109712 155278 109721
rect 155222 109647 155278 109656
rect 155420 480 155448 111007
rect 158902 109712 158958 109721
rect 158902 109647 158958 109656
rect 158916 480 158944 109647
rect 162504 480 162532 136031
rect 163516 3505 163544 250271
rect 174542 232928 174598 232937
rect 174542 232863 174598 232872
rect 166078 136232 166134 136241
rect 166078 136167 166134 136176
rect 163502 3496 163558 3505
rect 163502 3431 163558 3440
rect 166092 480 166120 136167
rect 174556 29889 174584 232863
rect 176658 138408 176714 138417
rect 176658 138343 176714 138352
rect 174542 29880 174598 29889
rect 174542 29815 174598 29824
rect 173162 3496 173218 3505
rect 173162 3431 173218 3440
rect 169574 3360 169630 3369
rect 169574 3295 169630 3304
rect 169588 480 169616 3295
rect 173176 480 173204 3431
rect 176672 480 176700 138343
rect 178696 27033 178724 256799
rect 182836 249762 182864 279414
rect 194612 260273 194640 390116
rect 198200 261225 198228 390116
rect 201788 262177 201816 390116
rect 205376 263401 205404 390116
rect 208964 264489 208992 390116
rect 212552 265577 212580 390116
rect 214654 382936 214710 382945
rect 214654 382871 214710 382880
rect 212538 265568 212594 265577
rect 212538 265503 212594 265512
rect 208950 264480 209006 264489
rect 208950 264415 209006 264424
rect 205362 263392 205418 263401
rect 205362 263327 205418 263336
rect 201774 262168 201830 262177
rect 201774 262103 201830 262112
rect 198186 261216 198242 261225
rect 198186 261151 198242 261160
rect 194598 260264 194654 260273
rect 194598 260199 194654 260208
rect 198002 253600 198058 253609
rect 198002 253535 198058 253544
rect 182824 249756 182876 249762
rect 182824 249698 182876 249704
rect 189724 249756 189776 249762
rect 189724 249698 189776 249704
rect 188342 242720 188398 242729
rect 188342 242655 188398 242664
rect 187330 139088 187386 139097
rect 187330 139023 187386 139032
rect 183742 138680 183798 138689
rect 183742 138615 183798 138624
rect 178682 27024 178738 27033
rect 178682 26959 178738 26968
rect 180246 3632 180302 3641
rect 180246 3567 180302 3576
rect 180260 480 180288 3567
rect 183756 480 183784 138615
rect 187344 480 187372 139023
rect 188356 53281 188384 242655
rect 189736 235278 189764 249698
rect 189724 235272 189776 235278
rect 189724 235214 189776 235220
rect 191102 230752 191158 230761
rect 191102 230687 191158 230696
rect 190826 129296 190882 129305
rect 190826 129231 190882 129240
rect 188342 53272 188398 53281
rect 188342 53207 188398 53216
rect 190840 480 190868 129231
rect 191116 124953 191144 230687
rect 195242 220824 195298 220833
rect 195242 220759 195298 220768
rect 194414 134736 194470 134745
rect 194414 134671 194470 134680
rect 191102 124944 191158 124953
rect 191102 124879 191158 124888
rect 194428 480 194456 134671
rect 195256 98705 195284 220759
rect 197910 131880 197966 131889
rect 197910 131815 197966 131824
rect 195242 98696 195298 98705
rect 195242 98631 195298 98640
rect 197924 480 197952 131815
rect 198016 102921 198044 253535
rect 202142 249248 202198 249257
rect 202142 249183 202198 249192
rect 199382 235104 199438 235113
rect 199382 235039 199438 235048
rect 198002 102912 198058 102921
rect 198002 102847 198058 102856
rect 199396 32745 199424 235039
rect 202156 141409 202184 249183
rect 209042 248160 209098 248169
rect 209042 248095 209098 248104
rect 207664 235272 207716 235278
rect 207664 235214 207716 235220
rect 206282 224224 206338 224233
rect 206282 224159 206338 224168
rect 203522 222048 203578 222057
rect 203522 221983 203578 221992
rect 202142 141400 202198 141409
rect 202142 141335 202198 141344
rect 201498 140040 201554 140049
rect 201498 139975 201554 139984
rect 199382 32736 199438 32745
rect 199382 32671 199438 32680
rect 201512 480 201540 139975
rect 203536 100065 203564 221983
rect 206296 144129 206324 224159
rect 207676 211818 207704 235214
rect 207664 211812 207716 211818
rect 207664 211754 207716 211760
rect 206282 144120 206338 144129
rect 206282 144055 206338 144064
rect 206282 139360 206338 139369
rect 206282 139295 206338 139304
rect 205640 139256 205692 139262
rect 205640 139198 205692 139204
rect 205652 138281 205680 139198
rect 205638 138272 205694 138281
rect 205638 138207 205694 138216
rect 203522 100056 203578 100065
rect 203522 99991 203578 100000
rect 206296 3777 206324 139295
rect 208582 132016 208638 132025
rect 208582 131951 208638 131960
rect 205086 3768 205142 3777
rect 205086 3703 205142 3712
rect 206282 3768 206338 3777
rect 206282 3703 206338 3712
rect 205100 480 205128 3703
rect 208596 480 208624 131951
rect 209056 101561 209084 248095
rect 211802 244896 211858 244905
rect 211802 244831 211858 244840
rect 210422 241496 210478 241505
rect 210422 241431 210478 241440
rect 209042 101552 209098 101561
rect 209042 101487 209098 101496
rect 210436 29753 210464 241431
rect 211816 123593 211844 244831
rect 214562 238368 214618 238377
rect 214562 238303 214618 238312
rect 213182 219872 213238 219881
rect 213182 219807 213238 219816
rect 212170 126440 212226 126449
rect 212170 126375 212226 126384
rect 211802 123584 211858 123593
rect 211802 123519 211858 123528
rect 210422 29744 210478 29753
rect 210422 29679 210478 29688
rect 212184 480 212212 126375
rect 213196 90545 213224 219807
rect 213182 90536 213238 90545
rect 213182 90471 213238 90480
rect 214576 31113 214604 238303
rect 214668 205601 214696 382871
rect 216140 266665 216168 390116
rect 219728 267753 219756 390116
rect 220176 343732 220228 343738
rect 220176 343674 220228 343680
rect 220084 343664 220136 343670
rect 220084 343606 220136 343612
rect 219714 267744 219770 267753
rect 219714 267679 219770 267688
rect 216126 266656 216182 266665
rect 216126 266591 216182 266600
rect 216034 245984 216090 245993
rect 216034 245919 216090 245928
rect 215942 223136 215998 223145
rect 215942 223071 215998 223080
rect 214654 205592 214710 205601
rect 214654 205527 214710 205536
rect 215300 139188 215352 139194
rect 215300 139130 215352 139136
rect 215312 138417 215340 139130
rect 215666 138544 215722 138553
rect 215666 138479 215722 138488
rect 215298 138408 215354 138417
rect 215298 138343 215354 138352
rect 214562 31104 214618 31113
rect 214562 31039 214618 31048
rect 215680 480 215708 138479
rect 215956 122233 215984 223071
rect 216048 195265 216076 245919
rect 218704 211812 218756 211818
rect 218704 211754 218756 211760
rect 218716 200054 218744 211754
rect 219438 200696 219494 200705
rect 219438 200631 219494 200640
rect 218704 200048 218756 200054
rect 218704 199990 218756 199996
rect 219452 199209 219480 200631
rect 220096 199850 220124 343606
rect 220084 199844 220136 199850
rect 220084 199786 220136 199792
rect 220188 199782 220216 343674
rect 223028 342440 223080 342446
rect 222934 342408 222990 342417
rect 223028 342382 223080 342388
rect 222934 342343 222990 342352
rect 220268 342304 220320 342310
rect 220268 342246 220320 342252
rect 220176 199776 220228 199782
rect 220176 199718 220228 199724
rect 220280 199714 220308 342246
rect 222842 259040 222898 259049
rect 222842 258975 222898 258984
rect 220268 199708 220320 199714
rect 220268 199650 220320 199656
rect 219438 199200 219494 199209
rect 219438 199135 219494 199144
rect 216034 195256 216090 195265
rect 216034 195191 216090 195200
rect 218060 139120 218112 139126
rect 218060 139062 218112 139068
rect 218072 138689 218100 139062
rect 218058 138680 218114 138689
rect 218058 138615 218114 138624
rect 219254 138680 219310 138689
rect 219254 138615 219310 138624
rect 215942 122224 215998 122233
rect 215942 122159 215998 122168
rect 219268 480 219296 138615
rect 222750 124944 222806 124953
rect 222750 124879 222806 124888
rect 222764 480 222792 124879
rect 222856 91769 222884 258975
rect 222948 198257 222976 342343
rect 223040 199646 223068 342382
rect 223120 341216 223172 341222
rect 223120 341158 223172 341164
rect 223028 199640 223080 199646
rect 223028 199582 223080 199588
rect 223132 198490 223160 341158
rect 223210 340912 223266 340921
rect 223210 340847 223266 340856
rect 223224 198665 223252 340847
rect 223316 268841 223344 390116
rect 226340 342508 226392 342514
rect 226340 342450 226392 342456
rect 226352 342417 226380 342450
rect 226338 342408 226394 342417
rect 226338 342343 226394 342352
rect 226616 342372 226668 342378
rect 226616 342314 226668 342320
rect 226628 342281 226656 342314
rect 226614 342272 226670 342281
rect 226614 342207 226670 342216
rect 225050 341864 225106 341873
rect 225050 341799 225106 341808
rect 224958 341592 225014 341601
rect 224958 341527 225014 341536
rect 224972 341154 225000 341527
rect 224960 341148 225012 341154
rect 224960 341090 225012 341096
rect 225064 341086 225092 341799
rect 225142 341728 225198 341737
rect 225142 341663 225198 341672
rect 225052 341080 225104 341086
rect 225052 341022 225104 341028
rect 225156 340950 225184 341663
rect 225786 341456 225842 341465
rect 225786 341391 225842 341400
rect 225696 341284 225748 341290
rect 225696 341226 225748 341232
rect 225144 340944 225196 340950
rect 225144 340886 225196 340892
rect 225602 340096 225658 340105
rect 225602 340031 225658 340040
rect 225418 339824 225474 339833
rect 225418 339759 225474 339768
rect 223488 339652 223540 339658
rect 223488 339594 223540 339600
rect 223396 339584 223448 339590
rect 223396 339526 223448 339532
rect 223302 268832 223358 268841
rect 223302 268767 223358 268776
rect 223302 226264 223358 226273
rect 223302 226199 223358 226208
rect 223210 198656 223266 198665
rect 223210 198591 223266 198600
rect 223120 198484 223172 198490
rect 223120 198426 223172 198432
rect 222934 198248 222990 198257
rect 222934 198183 222990 198192
rect 223316 181393 223344 226199
rect 223408 198422 223436 339526
rect 223500 198626 223528 339594
rect 225432 199617 225460 339759
rect 225418 199608 225474 199617
rect 225418 199543 225474 199552
rect 223488 198620 223540 198626
rect 223488 198562 223540 198568
rect 223396 198416 223448 198422
rect 223396 198358 223448 198364
rect 225616 197305 225644 340031
rect 225708 198558 225736 341226
rect 225696 198552 225748 198558
rect 225696 198494 225748 198500
rect 225800 197849 225828 341391
rect 225970 341184 226026 341193
rect 225970 341119 226026 341128
rect 225880 339720 225932 339726
rect 225880 339662 225932 339668
rect 225892 198694 225920 339662
rect 225984 199481 226012 341119
rect 226154 340776 226210 340785
rect 226154 340711 226210 340720
rect 225970 199472 226026 199481
rect 225970 199407 226026 199416
rect 226168 199345 226196 340711
rect 226904 269929 226932 390116
rect 228914 380760 228970 380769
rect 228914 380695 228970 380704
rect 228730 380352 228786 380361
rect 228730 380287 228786 380296
rect 228638 377360 228694 377369
rect 228638 377295 228694 377304
rect 227626 342272 227682 342281
rect 227626 342207 227682 342216
rect 227534 338464 227590 338473
rect 227534 338399 227590 338408
rect 226890 269920 226946 269929
rect 226890 269855 226946 269864
rect 227548 256737 227576 338399
rect 227640 257825 227668 342207
rect 227718 342136 227774 342145
rect 227718 342071 227774 342080
rect 227732 341018 227760 342071
rect 227812 341352 227864 341358
rect 227812 341294 227864 341300
rect 227720 341012 227772 341018
rect 227720 340954 227772 340960
rect 227824 340921 227852 341294
rect 228362 341048 228418 341057
rect 228362 340983 228418 340992
rect 227810 340912 227866 340921
rect 227810 340847 227866 340856
rect 228178 340912 228234 340921
rect 228178 340847 228234 340856
rect 227626 257816 227682 257825
rect 227626 257751 227682 257760
rect 227534 256728 227590 256737
rect 227534 256663 227590 256672
rect 226982 246936 227038 246945
rect 226982 246871 227038 246880
rect 226154 199336 226210 199345
rect 226154 199271 226210 199280
rect 226338 199200 226394 199209
rect 226338 199135 226394 199144
rect 225880 198688 225932 198694
rect 225880 198630 225932 198636
rect 226352 198121 226380 199135
rect 226338 198112 226394 198121
rect 226338 198047 226394 198056
rect 225786 197840 225842 197849
rect 225786 197775 225842 197784
rect 225602 197296 225658 197305
rect 225602 197231 225658 197240
rect 223302 181384 223358 181393
rect 223302 181319 223358 181328
rect 226338 123584 226394 123593
rect 226338 123519 226394 123528
rect 222842 91760 222898 91769
rect 222842 91695 222898 91704
rect 226352 480 226380 123519
rect 226996 120873 227024 246871
rect 228192 199753 228220 340847
rect 228270 339688 228326 339697
rect 228270 339623 228326 339632
rect 228284 199889 228312 339623
rect 228270 199880 228326 199889
rect 228270 199815 228326 199824
rect 228178 199744 228234 199753
rect 228178 199679 228234 199688
rect 228376 197985 228404 340983
rect 228546 340368 228602 340377
rect 228546 340303 228602 340312
rect 228456 339788 228508 339794
rect 228456 339730 228508 339736
rect 228468 199578 228496 339730
rect 228456 199572 228508 199578
rect 228456 199514 228508 199520
rect 228362 197976 228418 197985
rect 228362 197911 228418 197920
rect 228560 197577 228588 340303
rect 228652 327593 228680 377295
rect 228638 327584 228694 327593
rect 228638 327519 228694 327528
rect 228744 317801 228772 380287
rect 228822 380216 228878 380225
rect 228822 380151 228878 380160
rect 228836 322153 228864 380151
rect 228822 322144 228878 322153
rect 228822 322079 228878 322088
rect 228730 317792 228786 317801
rect 228730 317727 228786 317736
rect 228928 316713 228956 380695
rect 230386 380624 230442 380633
rect 230386 380559 230442 380568
rect 230202 378720 230258 378729
rect 230202 378655 230258 378664
rect 229006 374640 229062 374649
rect 229006 374575 229062 374584
rect 228730 316704 228786 316713
rect 228730 316639 228786 316648
rect 228914 316704 228970 316713
rect 228914 316639 228970 316648
rect 228744 202473 228772 316639
rect 229020 309097 229048 374575
rect 230216 328681 230244 378655
rect 230294 377496 230350 377505
rect 230294 377431 230350 377440
rect 230202 328672 230258 328681
rect 230202 328607 230258 328616
rect 230308 323241 230336 377431
rect 230294 323232 230350 323241
rect 230294 323167 230350 323176
rect 230400 318753 230428 380559
rect 230386 318744 230442 318753
rect 230386 318679 230442 318688
rect 229006 309088 229062 309097
rect 229006 309023 229062 309032
rect 230492 271017 230520 390116
rect 231766 387832 231822 387841
rect 231766 387767 231822 387776
rect 231582 382936 231638 382945
rect 231582 382871 231638 382880
rect 231490 376816 231546 376825
rect 231490 376751 231546 376760
rect 231216 342644 231268 342650
rect 231216 342586 231268 342592
rect 231030 338872 231086 338881
rect 231030 338807 231086 338816
rect 230938 338600 230994 338609
rect 230938 338535 230994 338544
rect 230478 271008 230534 271017
rect 230478 270943 230534 270952
rect 228914 251424 228970 251433
rect 228914 251359 228970 251368
rect 228730 202464 228786 202473
rect 228730 202399 228786 202408
rect 228546 197568 228602 197577
rect 228546 197503 228602 197512
rect 228928 192545 228956 251359
rect 230952 199073 230980 338535
rect 231044 199986 231072 338807
rect 231122 236192 231178 236201
rect 231122 236127 231178 236136
rect 231032 199980 231084 199986
rect 231032 199922 231084 199928
rect 230938 199064 230994 199073
rect 230938 198999 230994 199008
rect 228914 192536 228970 192545
rect 228914 192471 228970 192480
rect 226982 120864 227038 120873
rect 226982 120799 227038 120808
rect 231136 28393 231164 236127
rect 231228 198529 231256 342586
rect 231400 342576 231452 342582
rect 231400 342518 231452 342524
rect 231308 339448 231360 339454
rect 231308 339390 231360 339396
rect 231320 199918 231348 339390
rect 231308 199912 231360 199918
rect 231308 199854 231360 199860
rect 231214 198520 231270 198529
rect 231214 198455 231270 198464
rect 231412 198393 231440 342518
rect 231504 329633 231532 376751
rect 231490 329624 231546 329633
rect 231490 329559 231546 329568
rect 231596 313449 231624 382871
rect 231674 380488 231730 380497
rect 231674 380423 231730 380432
rect 231688 319977 231716 380423
rect 231674 319968 231730 319977
rect 231674 319903 231730 319912
rect 231582 313440 231638 313449
rect 231582 313375 231638 313384
rect 231398 198384 231454 198393
rect 231398 198319 231454 198328
rect 231780 193769 231808 387767
rect 233146 383344 233202 383353
rect 233146 383279 233202 383288
rect 233054 383072 233110 383081
rect 233054 383007 233110 383016
rect 232962 380896 233018 380905
rect 232962 380831 233018 380840
rect 232870 377768 232926 377777
rect 232870 377703 232926 377712
rect 232884 324329 232912 377703
rect 232870 324320 232926 324329
rect 232870 324255 232926 324264
rect 232976 314537 233004 380831
rect 232962 314528 233018 314537
rect 232962 314463 233018 314472
rect 233068 311273 233096 383007
rect 233054 311264 233110 311273
rect 233054 311199 233110 311208
rect 232594 222728 232650 222737
rect 232594 222663 232650 222672
rect 232502 221096 232558 221105
rect 232502 221031 232558 221040
rect 231766 193760 231822 193769
rect 231766 193695 231822 193704
rect 232516 138281 232544 221031
rect 232608 141953 232636 222663
rect 232686 219464 232742 219473
rect 232686 219399 232742 219408
rect 232700 142050 232728 219399
rect 232778 216200 232834 216209
rect 232778 216135 232834 216144
rect 232688 142044 232740 142050
rect 232688 141986 232740 141992
rect 232594 141944 232650 141953
rect 232594 141879 232650 141888
rect 232792 139777 232820 216135
rect 232962 214568 233018 214577
rect 232962 214503 233018 214512
rect 232976 140185 233004 214503
rect 233160 194857 233188 383279
rect 233698 377632 233754 377641
rect 233698 377567 233754 377576
rect 233712 325417 233740 377567
rect 233882 364984 233938 364993
rect 233882 364919 233938 364928
rect 233790 351384 233846 351393
rect 233790 351319 233846 351328
rect 233698 325408 233754 325417
rect 233698 325343 233754 325352
rect 233804 297129 233832 351319
rect 233896 308009 233924 364919
rect 233974 352608 234030 352617
rect 233974 352543 234030 352552
rect 233882 308000 233938 308009
rect 233882 307935 233938 307944
rect 233790 297120 233846 297129
rect 233790 297055 233846 297064
rect 233988 296041 234016 352543
rect 233974 296032 234030 296041
rect 233974 295967 234030 295976
rect 234080 274553 234108 390116
rect 234526 388512 234582 388521
rect 234526 388447 234582 388456
rect 234434 380080 234490 380089
rect 234434 380015 234490 380024
rect 234250 362536 234306 362545
rect 234250 362471 234306 362480
rect 234158 356960 234214 356969
rect 234158 356895 234214 356904
rect 234172 294953 234200 356895
rect 234158 294944 234214 294953
rect 234158 294879 234214 294888
rect 234264 290601 234292 362471
rect 234342 361040 234398 361049
rect 234342 360975 234398 360984
rect 234250 290592 234306 290601
rect 234250 290527 234306 290536
rect 234356 287337 234384 360975
rect 234448 306921 234476 380015
rect 234434 306912 234490 306921
rect 234434 306847 234490 306856
rect 234342 287328 234398 287337
rect 234342 287263 234398 287272
rect 234066 274544 234122 274553
rect 234066 274479 234122 274488
rect 233976 261520 234028 261526
rect 233976 261462 234028 261468
rect 233884 213988 233936 213994
rect 233884 213930 233936 213936
rect 233146 194848 233202 194857
rect 233146 194783 233202 194792
rect 232962 140176 233018 140185
rect 232962 140111 233018 140120
rect 232778 139768 232834 139777
rect 232778 139703 232834 139712
rect 233146 139088 233202 139097
rect 233146 139023 233202 139032
rect 233160 138922 233188 139023
rect 233148 138916 233200 138922
rect 233148 138858 233200 138864
rect 232502 138272 232558 138281
rect 232502 138207 232558 138216
rect 233896 138145 233924 213930
rect 233988 201482 234016 261462
rect 233976 201476 234028 201482
rect 233976 201418 234028 201424
rect 234540 195945 234568 388447
rect 235538 388376 235594 388385
rect 235538 388311 235594 388320
rect 235078 377904 235134 377913
rect 235078 377839 235134 377848
rect 235092 326505 235120 377839
rect 235446 374776 235502 374785
rect 235446 374711 235502 374720
rect 235354 359408 235410 359417
rect 235354 359343 235410 359352
rect 235262 354104 235318 354113
rect 235262 354039 235318 354048
rect 235170 350024 235226 350033
rect 235170 349959 235226 349968
rect 235078 326496 235134 326505
rect 235078 326431 235134 326440
rect 235184 304745 235212 349959
rect 235170 304736 235226 304745
rect 235170 304671 235226 304680
rect 235276 303521 235304 354039
rect 235368 305833 235396 359343
rect 235354 305824 235410 305833
rect 235354 305759 235410 305768
rect 235262 303512 235318 303521
rect 235262 303447 235318 303456
rect 235460 301481 235488 374711
rect 235446 301472 235502 301481
rect 235446 301407 235502 301416
rect 235552 300393 235580 388311
rect 237668 386889 237696 390116
rect 239218 387424 239274 387433
rect 239218 387359 239274 387368
rect 236458 386880 236514 386889
rect 236458 386815 236514 386824
rect 237654 386880 237710 386889
rect 237654 386815 237710 386824
rect 239034 386880 239090 386889
rect 239034 386815 239090 386824
rect 235814 356688 235870 356697
rect 235814 356623 235870 356632
rect 235630 343768 235686 343777
rect 235630 343703 235686 343712
rect 235538 300384 235594 300393
rect 235538 300319 235594 300328
rect 235538 207088 235594 207097
rect 235538 207023 235594 207032
rect 234894 206408 234950 206417
rect 234894 206343 234950 206352
rect 234526 195936 234582 195945
rect 234526 195871 234582 195880
rect 234908 151814 234936 206343
rect 235262 201512 235318 201521
rect 235262 201447 235318 201456
rect 234908 151786 235120 151814
rect 235092 138281 235120 151786
rect 235276 139913 235304 201447
rect 235448 197668 235500 197674
rect 235448 197610 235500 197616
rect 235356 197532 235408 197538
rect 235356 197474 235408 197480
rect 235368 140350 235396 197474
rect 235356 140344 235408 140350
rect 235356 140286 235408 140292
rect 235460 140282 235488 197610
rect 235552 192681 235580 207023
rect 235644 204921 235672 343703
rect 235724 339516 235776 339522
rect 235724 339458 235776 339464
rect 235630 204912 235686 204921
rect 235630 204847 235686 204856
rect 235538 192672 235594 192681
rect 235538 192607 235594 192616
rect 235736 184929 235764 339458
rect 235828 187241 235856 356623
rect 235906 348528 235962 348537
rect 235906 348463 235962 348472
rect 235814 187232 235870 187241
rect 235814 187167 235870 187176
rect 235722 184920 235778 184929
rect 235722 184855 235778 184864
rect 235920 143721 235948 348463
rect 236472 329769 236500 386815
rect 238574 376000 238630 376009
rect 238574 375935 238630 375944
rect 236826 369200 236882 369209
rect 236826 369135 236882 369144
rect 236734 362264 236790 362273
rect 236734 362199 236790 362208
rect 236550 345672 236606 345681
rect 236550 345607 236606 345616
rect 236458 329760 236514 329769
rect 236458 329695 236514 329704
rect 236564 310185 236592 345607
rect 236644 341624 236696 341630
rect 236644 341566 236696 341572
rect 236550 310176 236606 310185
rect 236550 310111 236606 310120
rect 236656 299305 236684 341566
rect 236748 315625 236776 362199
rect 236840 321065 236868 369135
rect 237930 369064 237986 369073
rect 237930 368999 237986 369008
rect 237286 355328 237342 355337
rect 237286 355263 237342 355272
rect 237194 353968 237250 353977
rect 237194 353903 237250 353912
rect 237010 351112 237066 351121
rect 237010 351047 237066 351056
rect 236920 341556 236972 341562
rect 236920 341498 236972 341504
rect 236826 321056 236882 321065
rect 236826 320991 236882 321000
rect 236734 315616 236790 315625
rect 236734 315551 236790 315560
rect 236932 312361 236960 341498
rect 236918 312352 236974 312361
rect 236918 312287 236974 312296
rect 236642 299296 236698 299305
rect 236642 299231 236698 299240
rect 237024 289785 237052 351047
rect 237104 340264 237156 340270
rect 237104 340206 237156 340212
rect 237010 289776 237066 289785
rect 237010 289711 237066 289720
rect 237116 191593 237144 340206
rect 237102 191584 237158 191593
rect 237102 191519 237158 191528
rect 237208 190369 237236 353903
rect 237194 190360 237250 190369
rect 237194 190295 237250 190304
rect 237300 146985 237328 355263
rect 237472 341760 237524 341766
rect 237472 341702 237524 341708
rect 237380 341488 237432 341494
rect 237378 341456 237380 341465
rect 237432 341456 237434 341465
rect 237378 341391 237434 341400
rect 237484 341057 237512 341702
rect 237746 341456 237802 341465
rect 237746 341391 237802 341400
rect 237470 341048 237526 341057
rect 237470 340983 237526 340992
rect 237470 340368 237526 340377
rect 237470 340303 237526 340312
rect 237484 340134 237512 340303
rect 237472 340128 237524 340134
rect 237378 340096 237434 340105
rect 237472 340070 237524 340076
rect 237378 340031 237434 340040
rect 237564 340060 237616 340066
rect 237392 339862 237420 340031
rect 237564 340002 237616 340008
rect 237380 339856 237432 339862
rect 237380 339798 237432 339804
rect 237576 339697 237604 340002
rect 237562 339688 237618 339697
rect 237562 339623 237618 339632
rect 237654 333296 237710 333305
rect 237654 333231 237710 333240
rect 237668 275369 237696 333231
rect 237760 285161 237788 341391
rect 237838 340096 237894 340105
rect 237838 340031 237894 340040
rect 237852 291689 237880 340031
rect 237944 331945 237972 368999
rect 238482 351248 238538 351257
rect 238482 351183 238538 351192
rect 238022 345944 238078 345953
rect 238022 345879 238078 345888
rect 238036 345014 238064 345879
rect 238036 344986 238340 345014
rect 238206 341592 238262 341601
rect 238036 341550 238206 341578
rect 238036 337414 238064 341550
rect 238206 341527 238262 341536
rect 238206 340368 238262 340377
rect 238206 340303 238262 340312
rect 238114 340232 238170 340241
rect 238114 340167 238170 340176
rect 238024 337408 238076 337414
rect 238024 337350 238076 337356
rect 237930 331936 237986 331945
rect 237930 331871 237986 331880
rect 237930 331120 237986 331129
rect 237930 331055 237986 331064
rect 237838 291680 237894 291689
rect 237838 291615 237894 291624
rect 237746 285152 237802 285161
rect 237746 285087 237802 285096
rect 237944 279721 237972 331055
rect 238022 329760 238078 329769
rect 238022 329695 238078 329704
rect 237930 279712 237986 279721
rect 237930 279647 237986 279656
rect 237654 275360 237710 275369
rect 237654 275295 237710 275304
rect 237378 274544 237434 274553
rect 237378 274479 237434 274488
rect 237392 272105 237420 274479
rect 238036 273193 238064 329695
rect 238128 289513 238156 340167
rect 238114 289504 238170 289513
rect 238114 289439 238170 289448
rect 238220 288425 238248 340303
rect 238312 292777 238340 344986
rect 238392 340332 238444 340338
rect 238392 340274 238444 340280
rect 238404 337521 238432 340274
rect 238390 337512 238446 337521
rect 238390 337447 238446 337456
rect 238392 337408 238444 337414
rect 238392 337350 238444 337356
rect 238298 292768 238354 292777
rect 238298 292703 238354 292712
rect 238206 288416 238262 288425
rect 238206 288351 238262 288360
rect 238404 286249 238432 337350
rect 238496 330857 238524 351183
rect 238588 333033 238616 375935
rect 238666 339416 238722 339425
rect 238666 339351 238722 339360
rect 238574 333024 238630 333033
rect 238574 332959 238630 332968
rect 238482 330848 238538 330857
rect 238482 330783 238538 330792
rect 238390 286240 238446 286249
rect 238390 286175 238446 286184
rect 238680 274281 238708 339351
rect 239048 333305 239076 386815
rect 239126 341728 239182 341737
rect 239126 341663 239182 341672
rect 239140 338570 239168 341663
rect 239128 338564 239180 338570
rect 239128 338506 239180 338512
rect 239034 333296 239090 333305
rect 239034 333231 239090 333240
rect 239232 331129 239260 387359
rect 239586 346080 239642 346089
rect 239586 346015 239642 346024
rect 239494 344312 239550 344321
rect 239494 344247 239550 344256
rect 239402 342952 239458 342961
rect 239402 342887 239458 342896
rect 239310 340640 239366 340649
rect 239310 340575 239366 340584
rect 239218 331120 239274 331129
rect 239218 331055 239274 331064
rect 239324 280809 239352 340575
rect 239416 282849 239444 342887
rect 239402 282840 239458 282849
rect 239402 282775 239458 282784
rect 239508 281897 239536 344247
rect 239600 284073 239628 346015
rect 240048 342712 240100 342718
rect 240048 342654 240100 342660
rect 240060 342281 240088 342654
rect 240046 342272 240102 342281
rect 240046 342207 240102 342216
rect 240048 341828 240100 341834
rect 240048 341770 240100 341776
rect 240060 340921 240088 341770
rect 240784 341420 240836 341426
rect 240784 341362 240836 341368
rect 240046 340912 240102 340921
rect 240046 340847 240102 340856
rect 239954 340776 240010 340785
rect 239954 340711 240010 340720
rect 239678 340504 239734 340513
rect 239678 340439 239734 340448
rect 239586 284064 239642 284073
rect 239586 283999 239642 284008
rect 239494 281888 239550 281897
rect 239494 281823 239550 281832
rect 239310 280800 239366 280809
rect 239310 280735 239366 280744
rect 239692 276389 239720 340439
rect 239864 340400 239916 340406
rect 239864 340342 239916 340348
rect 239876 339833 239904 340342
rect 239968 339998 239996 340711
rect 239956 339992 240008 339998
rect 239956 339934 240008 339940
rect 240046 339960 240102 339969
rect 240796 339932 240824 341362
rect 240046 339895 240048 339904
rect 240100 339895 240102 339904
rect 240048 339866 240100 339872
rect 239862 339824 239918 339833
rect 240046 339824 240102 339833
rect 239862 339759 239918 339768
rect 239968 339782 240046 339810
rect 239968 339402 239996 339782
rect 240046 339759 240102 339768
rect 241256 339425 241284 390116
rect 244844 386889 244872 390116
rect 244830 386880 244886 386889
rect 244830 386815 244886 386824
rect 248432 364334 248460 390116
rect 249890 387696 249946 387705
rect 249890 387631 249946 387640
rect 248432 364306 248552 364334
rect 241794 363760 241850 363769
rect 241794 363695 241850 363704
rect 241808 339932 241836 363695
rect 246302 358048 246358 358057
rect 246302 357983 246358 357992
rect 242808 345024 242860 345030
rect 242714 344992 242770 345001
rect 242808 344966 242860 344972
rect 242714 344927 242770 344936
rect 242728 340898 242756 344927
rect 242820 343777 242848 344966
rect 242806 343768 242862 343777
rect 242806 343703 242862 343712
rect 245842 343224 245898 343233
rect 245842 343159 245898 343168
rect 245658 343088 245714 343097
rect 245658 343023 245714 343032
rect 245672 342990 245700 343023
rect 245660 342984 245712 342990
rect 245660 342926 245712 342932
rect 243544 342848 243596 342854
rect 243544 342790 243596 342796
rect 244830 342816 244886 342825
rect 243556 342689 243584 342790
rect 244280 342780 244332 342786
rect 244830 342751 244886 342760
rect 244280 342722 244332 342728
rect 243542 342680 243598 342689
rect 243542 342615 243598 342624
rect 244292 342553 244320 342722
rect 244278 342544 244334 342553
rect 244278 342479 244334 342488
rect 243818 342272 243874 342281
rect 243818 342207 243874 342216
rect 242728 340870 242848 340898
rect 242820 339932 242848 340870
rect 243832 339932 243860 342207
rect 244844 339932 244872 342751
rect 245856 339932 245884 343159
rect 246316 342281 246344 357983
rect 247038 343632 247094 343641
rect 247038 343567 247094 343576
rect 247052 342922 247080 343567
rect 247866 343088 247922 343097
rect 247866 343023 247922 343032
rect 247040 342916 247092 342922
rect 247040 342858 247092 342864
rect 246854 342544 246910 342553
rect 246854 342479 246910 342488
rect 246302 342272 246358 342281
rect 246302 342207 246358 342216
rect 246868 339932 246896 342479
rect 247880 339932 247908 343023
rect 248524 340513 248552 364306
rect 249708 343052 249760 343058
rect 249708 342994 249760 343000
rect 248878 342680 248934 342689
rect 248878 342615 248934 342624
rect 248510 340504 248566 340513
rect 248510 340439 248566 340448
rect 248892 339932 248920 342615
rect 249720 342417 249748 342994
rect 249706 342408 249762 342417
rect 249706 342343 249762 342352
rect 249904 339932 249932 387631
rect 251914 387560 251970 387569
rect 251914 387495 251970 387504
rect 251086 343496 251142 343505
rect 251086 343431 251142 343440
rect 250902 343360 250958 343369
rect 250902 343295 250958 343304
rect 250916 339932 250944 343295
rect 251100 343126 251128 343431
rect 251088 343120 251140 343126
rect 251088 343062 251140 343068
rect 251928 339932 251956 387495
rect 252020 364334 252048 390116
rect 254950 369336 255006 369345
rect 254950 369271 255006 369280
rect 253938 367704 253994 367713
rect 253938 367639 253994 367648
rect 252020 364306 252232 364334
rect 252204 339969 252232 364306
rect 252926 344856 252982 344865
rect 252926 344791 252982 344800
rect 252190 339960 252246 339969
rect 252940 339932 252968 344791
rect 253202 344584 253258 344593
rect 253202 344519 253258 344528
rect 253216 343874 253244 344519
rect 253204 343868 253256 343874
rect 253204 343810 253256 343816
rect 253952 339932 253980 367639
rect 254964 339932 254992 369271
rect 255318 344176 255374 344185
rect 255318 344111 255374 344120
rect 255332 343806 255360 344111
rect 255320 343800 255372 343806
rect 255320 343742 255372 343748
rect 255608 341737 255636 390116
rect 259196 387433 259224 390116
rect 259182 387424 259238 387433
rect 259182 387359 259238 387368
rect 256054 386880 256110 386889
rect 256054 386815 256110 386824
rect 255962 344720 256018 344729
rect 255962 344655 256018 344664
rect 255594 341728 255650 341737
rect 255594 341663 255650 341672
rect 255976 339932 256004 344655
rect 256068 343097 256096 386815
rect 258722 386744 258778 386753
rect 258722 386679 258778 386688
rect 257986 381712 258042 381721
rect 257986 381647 258042 381656
rect 256974 344584 257030 344593
rect 256974 344519 257030 344528
rect 256698 344448 256754 344457
rect 256698 344383 256754 344392
rect 256712 343942 256740 344383
rect 256700 343936 256752 343942
rect 256700 343878 256752 343884
rect 256054 343088 256110 343097
rect 256054 343023 256110 343032
rect 256988 339932 257016 344519
rect 258000 339932 258028 381647
rect 258736 343233 258764 386679
rect 260748 378140 260800 378146
rect 260748 378082 260800 378088
rect 260010 377224 260066 377233
rect 260010 377159 260066 377168
rect 258998 371920 259054 371929
rect 258998 371855 259054 371864
rect 258722 343224 258778 343233
rect 258722 343159 258778 343168
rect 259012 339932 259040 371855
rect 260024 339932 260052 377159
rect 260760 376825 260788 378082
rect 260746 376816 260802 376825
rect 260746 376751 260802 376760
rect 261022 373416 261078 373425
rect 261022 373351 261078 373360
rect 261036 339932 261064 373351
rect 262034 342272 262090 342281
rect 262034 342207 262090 342216
rect 262048 339932 262076 342207
rect 262784 340649 262812 390116
rect 265624 389836 265676 389842
rect 265624 389778 265676 389784
rect 265636 377466 265664 389778
rect 265624 377460 265676 377466
rect 265624 377402 265676 377408
rect 264242 370696 264298 370705
rect 264242 370631 264298 370640
rect 262862 359544 262918 359553
rect 262862 359479 262918 359488
rect 262876 342281 262904 359479
rect 264058 344448 264114 344457
rect 264058 344383 264114 344392
rect 263598 344040 263654 344049
rect 263598 343975 263600 343984
rect 263652 343975 263654 343984
rect 263600 343946 263652 343952
rect 262862 342272 262918 342281
rect 262862 342207 262918 342216
rect 263046 342272 263102 342281
rect 263046 342207 263102 342216
rect 262770 340640 262826 340649
rect 262770 340575 262826 340584
rect 263060 339932 263088 342207
rect 264072 339932 264100 344383
rect 264256 342281 264284 370631
rect 265070 366344 265126 366353
rect 265070 366279 265126 366288
rect 264242 342272 264298 342281
rect 264242 342207 264298 342216
rect 265084 339932 265112 366279
rect 266372 344321 266400 390116
rect 267094 365120 267150 365129
rect 267094 365055 267150 365064
rect 267002 360904 267058 360913
rect 267002 360839 267058 360848
rect 267016 345014 267044 360839
rect 266464 344986 267044 345014
rect 266358 344312 266414 344321
rect 266358 344247 266414 344256
rect 266464 342394 266492 344986
rect 266280 342366 266492 342394
rect 266280 339946 266308 342366
rect 266110 339918 266308 339946
rect 267108 339932 267136 365055
rect 268106 344312 268162 344321
rect 268106 344247 268162 344256
rect 268120 339932 268148 344247
rect 269960 342961 269988 390116
rect 272524 387728 272576 387734
rect 272524 387670 272576 387676
rect 270408 387592 270460 387598
rect 270408 387534 270460 387540
rect 270130 387424 270186 387433
rect 270130 387359 270186 387368
rect 269946 342952 270002 342961
rect 269946 342887 270002 342896
rect 269118 342272 269174 342281
rect 269118 342207 269174 342216
rect 269132 339932 269160 342207
rect 270144 339932 270172 387359
rect 270420 387297 270448 387534
rect 270406 387288 270462 387297
rect 270406 387223 270462 387232
rect 272536 387025 272564 387670
rect 273166 387288 273222 387297
rect 273166 387223 273222 387232
rect 272522 387016 272578 387025
rect 272522 386951 272578 386960
rect 271234 378856 271290 378865
rect 271234 378791 271290 378800
rect 271142 376272 271198 376281
rect 271142 376207 271198 376216
rect 271156 339932 271184 376207
rect 271248 342281 271276 378791
rect 272524 377460 272576 377466
rect 272524 377402 272576 377408
rect 272536 351218 272564 377402
rect 272524 351212 272576 351218
rect 272524 351154 272576 351160
rect 271234 342272 271290 342281
rect 271234 342207 271290 342216
rect 272154 342272 272210 342281
rect 272154 342207 272210 342216
rect 272168 339932 272196 342207
rect 273180 339932 273208 387223
rect 273548 346089 273576 390116
rect 274640 387660 274692 387666
rect 274640 387602 274692 387608
rect 274652 387161 274680 387602
rect 274638 387152 274694 387161
rect 274638 387087 274694 387096
rect 275190 387016 275246 387025
rect 275190 386951 275246 386960
rect 273902 362400 273958 362409
rect 273902 362335 273958 362344
rect 273534 346080 273590 346089
rect 273534 346015 273590 346024
rect 273916 342281 273944 362335
rect 274178 356824 274234 356833
rect 274178 356759 274234 356768
rect 273902 342272 273958 342281
rect 273902 342207 273958 342216
rect 274192 339932 274220 356759
rect 275204 339932 275232 386951
rect 276202 343224 276258 343233
rect 276202 343159 276258 343168
rect 276216 339932 276244 343159
rect 277136 341465 277164 390116
rect 277216 387184 277268 387190
rect 277216 387126 277268 387132
rect 277122 341456 277178 341465
rect 277122 341391 277178 341400
rect 277228 339932 277256 387126
rect 280252 343936 280304 343942
rect 280252 343878 280304 343884
rect 278226 343088 278282 343097
rect 278226 343023 278282 343032
rect 278240 339932 278268 343023
rect 279238 342952 279294 342961
rect 279238 342887 279294 342896
rect 279252 339932 279280 342887
rect 252190 339895 252246 339904
rect 239784 339374 239996 339402
rect 241242 339416 241298 339425
rect 239784 277454 239812 339374
rect 241242 339351 241298 339360
rect 239864 338564 239916 338570
rect 239864 338506 239916 338512
rect 239876 278565 239904 338506
rect 280158 338464 280214 338473
rect 280158 338399 280214 338408
rect 239862 278556 239918 278565
rect 239862 278491 239918 278500
rect 239862 277468 239918 277477
rect 239784 277426 239862 277454
rect 239862 277403 239918 277412
rect 239678 276380 239734 276389
rect 239678 276315 239734 276324
rect 238666 274272 238722 274281
rect 238666 274207 238722 274216
rect 238022 273184 238078 273193
rect 238022 273119 238078 273128
rect 237378 272096 237434 272105
rect 237378 272031 237434 272040
rect 238206 260128 238262 260137
rect 238206 260063 238262 260072
rect 238114 255640 238170 255649
rect 238114 255575 238170 255584
rect 238022 225176 238078 225185
rect 238022 225111 238078 225120
rect 237378 214296 237434 214305
rect 237378 214231 237434 214240
rect 237392 213994 237420 214231
rect 237380 213988 237432 213994
rect 237380 213930 237432 213936
rect 237380 201476 237432 201482
rect 237380 201418 237432 201424
rect 237392 201385 237420 201418
rect 237378 201376 237434 201385
rect 237378 201311 237434 201320
rect 237380 200048 237432 200054
rect 237380 199990 237432 199996
rect 237392 199209 237420 199990
rect 237378 199200 237434 199209
rect 237378 199135 237434 199144
rect 237286 146976 237342 146985
rect 237286 146911 237342 146920
rect 238036 146146 238064 225111
rect 238128 193905 238156 255575
rect 238220 200297 238248 260063
rect 280172 256057 280200 338399
rect 280264 263537 280292 343878
rect 280620 341828 280672 341834
rect 280620 341770 280672 341776
rect 280344 341760 280396 341766
rect 280344 341702 280396 341708
rect 280356 295225 280384 341702
rect 280436 340128 280488 340134
rect 280436 340070 280488 340076
rect 280342 295216 280398 295225
rect 280342 295151 280398 295160
rect 280448 293865 280476 340070
rect 280526 338600 280582 338609
rect 280526 338535 280582 338544
rect 280434 293856 280490 293865
rect 280434 293791 280490 293800
rect 280540 292505 280568 338535
rect 280632 296449 280660 341770
rect 280724 341601 280752 390116
rect 282182 384432 282238 384441
rect 282182 384367 282238 384376
rect 281540 342644 281592 342650
rect 281540 342586 281592 342592
rect 280710 341592 280766 341601
rect 280710 341527 280766 341536
rect 280712 341488 280764 341494
rect 280712 341430 280764 341436
rect 280724 297809 280752 341430
rect 280894 341184 280950 341193
rect 280894 341119 280950 341128
rect 280804 340060 280856 340066
rect 280804 340002 280856 340008
rect 280710 297800 280766 297809
rect 280710 297735 280766 297744
rect 280618 296440 280674 296449
rect 280618 296375 280674 296384
rect 280816 296041 280844 340002
rect 280908 299441 280936 341119
rect 280988 340400 281040 340406
rect 280988 340342 281040 340348
rect 280894 299432 280950 299441
rect 280894 299367 280950 299376
rect 281000 298081 281028 340342
rect 280986 298072 281042 298081
rect 280986 298007 281042 298016
rect 280802 296032 280858 296041
rect 280802 295967 280858 295976
rect 280526 292496 280582 292505
rect 280526 292431 280582 292440
rect 281552 289513 281580 342586
rect 281724 339788 281776 339794
rect 281724 339730 281776 339736
rect 281632 339448 281684 339454
rect 281632 339390 281684 339396
rect 281644 291145 281672 339390
rect 281736 293593 281764 339730
rect 282196 319569 282224 384367
rect 282274 383208 282330 383217
rect 282274 383143 282330 383152
rect 282288 323649 282316 383143
rect 282828 380860 282880 380866
rect 282828 380802 282880 380808
rect 282840 379545 282868 380802
rect 282826 379536 282882 379545
rect 282826 379471 282882 379480
rect 282828 378072 282880 378078
rect 282828 378014 282880 378020
rect 282840 376825 282868 378014
rect 282826 376816 282882 376825
rect 282826 376751 282882 376760
rect 282918 376136 282974 376145
rect 282918 376071 282974 376080
rect 282366 338872 282422 338881
rect 282366 338807 282422 338816
rect 282274 323640 282330 323649
rect 282274 323575 282330 323584
rect 282182 319560 282238 319569
rect 282182 319495 282238 319504
rect 282380 317121 282408 338807
rect 282458 331800 282514 331809
rect 282458 331735 282514 331744
rect 282366 317112 282422 317121
rect 282366 317047 282422 317056
rect 282472 315489 282500 331735
rect 282550 330440 282606 330449
rect 282550 330375 282606 330384
rect 282458 315480 282514 315489
rect 282458 315415 282514 315424
rect 282564 313857 282592 330375
rect 282550 313848 282606 313857
rect 282550 313783 282606 313792
rect 282184 299464 282236 299470
rect 282182 299432 282184 299441
rect 282236 299432 282238 299441
rect 282182 299367 282238 299376
rect 281722 293584 281778 293593
rect 281722 293519 281778 293528
rect 281630 291136 281686 291145
rect 281630 291071 281686 291080
rect 282184 289808 282236 289814
rect 282182 289776 282184 289785
rect 282236 289776 282238 289785
rect 282182 289711 282238 289720
rect 281538 289504 281594 289513
rect 281538 289439 281594 289448
rect 282092 288380 282144 288386
rect 282092 288322 282144 288328
rect 282104 288289 282132 288322
rect 282736 288312 282788 288318
rect 282090 288280 282146 288289
rect 282736 288254 282788 288260
rect 282090 288215 282146 288224
rect 282748 288017 282776 288254
rect 282734 288008 282790 288017
rect 282734 287943 282790 287952
rect 282644 286748 282696 286754
rect 282644 286690 282696 286696
rect 282656 286657 282684 286690
rect 282642 286648 282698 286657
rect 282642 286583 282698 286592
rect 281540 285660 281592 285666
rect 281540 285602 281592 285608
rect 281552 285569 281580 285602
rect 282644 285592 282696 285598
rect 281538 285560 281594 285569
rect 281538 285495 281594 285504
rect 282642 285560 282644 285569
rect 282696 285560 282698 285569
rect 282642 285495 282698 285504
rect 282092 284300 282144 284306
rect 282092 284242 282144 284248
rect 282104 284209 282132 284242
rect 282090 284200 282146 284209
rect 282090 284135 282146 284144
rect 282000 281512 282052 281518
rect 281998 281480 282000 281489
rect 282052 281480 282054 281489
rect 281998 281415 282054 281424
rect 282000 280152 282052 280158
rect 282000 280094 282052 280100
rect 282012 279721 282040 280094
rect 281998 279712 282054 279721
rect 281998 279647 282054 279656
rect 282826 277808 282882 277817
rect 282826 277743 282882 277752
rect 282840 277506 282868 277743
rect 282828 277500 282880 277506
rect 282828 277442 282880 277448
rect 282734 277400 282790 277409
rect 282734 277335 282790 277344
rect 282748 276078 282776 277335
rect 282826 276312 282882 276321
rect 282826 276247 282882 276256
rect 282840 276146 282868 276247
rect 282828 276140 282880 276146
rect 282828 276082 282880 276088
rect 282736 276072 282788 276078
rect 282736 276014 282788 276020
rect 282826 275224 282882 275233
rect 282826 275159 282882 275168
rect 282840 274718 282868 275159
rect 282828 274712 282880 274718
rect 282828 274654 282880 274660
rect 282734 273728 282790 273737
rect 282734 273663 282790 273672
rect 282748 273290 282776 273663
rect 282828 273352 282880 273358
rect 282826 273320 282828 273329
rect 282880 273320 282882 273329
rect 282736 273284 282788 273290
rect 282826 273255 282882 273264
rect 282736 273226 282788 273232
rect 282826 272232 282882 272241
rect 282826 272167 282882 272176
rect 282840 271930 282868 272167
rect 282828 271924 282880 271930
rect 282828 271866 282880 271872
rect 282734 271144 282790 271153
rect 282734 271079 282790 271088
rect 282748 270570 282776 271079
rect 282826 270736 282882 270745
rect 282826 270671 282882 270680
rect 282840 270638 282868 270671
rect 282828 270632 282880 270638
rect 282828 270574 282880 270580
rect 282736 270564 282788 270570
rect 282736 270506 282788 270512
rect 281908 270496 281960 270502
rect 281908 270438 281960 270444
rect 281920 270065 281948 270438
rect 281906 270056 281962 270065
rect 281906 269991 281962 270000
rect 281908 267708 281960 267714
rect 281908 267650 281960 267656
rect 281920 267617 281948 267650
rect 281906 267608 281962 267617
rect 281906 267543 281962 267552
rect 281816 266348 281868 266354
rect 281816 266290 281868 266296
rect 281828 265985 281856 266290
rect 281814 265976 281870 265985
rect 281814 265911 281870 265920
rect 280250 263528 280306 263537
rect 280250 263463 280306 263472
rect 282828 262200 282880 262206
rect 282828 262142 282880 262148
rect 282840 262041 282868 262142
rect 282826 262032 282882 262041
rect 282826 261967 282882 261976
rect 282552 260840 282604 260846
rect 282550 260808 282552 260817
rect 282604 260808 282606 260817
rect 282550 260743 282606 260752
rect 282552 257508 282604 257514
rect 282552 257450 282604 257456
rect 282564 257417 282592 257450
rect 282550 257408 282606 257417
rect 282550 257343 282606 257352
rect 282828 256692 282880 256698
rect 282828 256634 282880 256640
rect 282840 256465 282868 256634
rect 282826 256456 282882 256465
rect 282826 256391 282882 256400
rect 280158 256048 280214 256057
rect 280158 255983 280214 255992
rect 282828 253904 282880 253910
rect 282828 253846 282880 253852
rect 282840 253473 282868 253846
rect 282826 253464 282882 253473
rect 282826 253399 282882 253408
rect 282826 242992 282882 243001
rect 282826 242927 282828 242936
rect 282880 242927 282882 242936
rect 282828 242898 282880 242904
rect 281538 239320 281594 239329
rect 281538 239255 281594 239264
rect 280158 237416 280214 237425
rect 280158 237351 280214 237360
rect 238666 216744 238722 216753
rect 238666 216679 238722 216688
rect 238390 204912 238446 204921
rect 238390 204847 238446 204856
rect 238206 200288 238262 200297
rect 238206 200223 238262 200232
rect 238300 197464 238352 197470
rect 238300 197406 238352 197412
rect 238208 197396 238260 197402
rect 238208 197338 238260 197344
rect 238114 193896 238170 193905
rect 238114 193831 238170 193840
rect 238220 151814 238248 197338
rect 237852 146118 238064 146146
rect 238128 151786 238248 151814
rect 235906 143712 235962 143721
rect 235906 143647 235962 143656
rect 236828 142044 236880 142050
rect 236828 141986 236880 141992
rect 235906 140720 235962 140729
rect 235906 140655 235962 140664
rect 235448 140276 235500 140282
rect 235448 140218 235500 140224
rect 235920 140214 235948 140655
rect 235908 140208 235960 140214
rect 235908 140150 235960 140156
rect 235262 139904 235318 139913
rect 235262 139839 235318 139848
rect 235722 139360 235778 139369
rect 235722 139295 235778 139304
rect 235632 138984 235684 138990
rect 235632 138926 235684 138932
rect 235644 138825 235672 138926
rect 235630 138816 235686 138825
rect 235630 138751 235686 138760
rect 235736 138650 235764 139295
rect 236840 139233 236868 141986
rect 237746 140720 237802 140729
rect 237746 140655 237802 140664
rect 237760 140622 237788 140655
rect 237748 140616 237800 140622
rect 237748 140558 237800 140564
rect 236826 139224 236882 139233
rect 236826 139159 236882 139168
rect 235908 139052 235960 139058
rect 235908 138994 235960 139000
rect 235920 138961 235948 138994
rect 235906 138952 235962 138961
rect 235906 138887 235962 138896
rect 235816 138780 235868 138786
rect 235816 138722 235868 138728
rect 235724 138644 235776 138650
rect 235724 138586 235776 138592
rect 235828 138553 235856 138722
rect 235908 138712 235960 138718
rect 235906 138680 235908 138689
rect 235960 138680 235962 138689
rect 235906 138615 235962 138624
rect 235814 138544 235870 138553
rect 235814 138479 235870 138488
rect 235078 138272 235134 138281
rect 235078 138207 235134 138216
rect 233882 138136 233938 138145
rect 233882 138071 233938 138080
rect 237852 138014 237880 146118
rect 238128 146010 238156 151786
rect 238036 145982 238156 146010
rect 238036 140146 238064 145982
rect 238312 145874 238340 197406
rect 238404 197033 238432 204847
rect 238680 203561 238708 216679
rect 238666 203552 238722 203561
rect 238666 203487 238722 203496
rect 280066 201512 280122 201521
rect 280066 201447 280122 201456
rect 238668 197736 238720 197742
rect 238668 197678 238720 197684
rect 238484 197600 238536 197606
rect 238484 197542 238536 197548
rect 238390 197024 238446 197033
rect 238390 196959 238446 196968
rect 238496 151814 238524 197542
rect 238574 183832 238630 183841
rect 238574 183767 238630 183776
rect 238128 145846 238340 145874
rect 238404 151786 238524 151814
rect 238024 140140 238076 140146
rect 238024 140082 238076 140088
rect 238128 140078 238156 145846
rect 238206 145752 238262 145761
rect 238206 145687 238262 145696
rect 238116 140072 238168 140078
rect 238116 140014 238168 140020
rect 238220 139398 238248 145687
rect 238404 141817 238432 151786
rect 238588 147674 238616 183767
rect 238496 147646 238616 147674
rect 238390 141808 238446 141817
rect 238390 141743 238446 141752
rect 238496 141522 238524 147646
rect 238680 144650 238708 197678
rect 239770 178460 239826 178469
rect 239770 178395 239826 178404
rect 238588 144622 238708 144650
rect 238588 141681 238616 144622
rect 238574 141672 238630 141681
rect 238574 141607 238630 141616
rect 238496 141494 238616 141522
rect 238482 140720 238538 140729
rect 238482 140655 238484 140664
rect 238536 140655 238538 140664
rect 238484 140626 238536 140632
rect 238588 140554 238616 141494
rect 239586 141400 239642 141409
rect 239586 141335 239642 141344
rect 238576 140548 238628 140554
rect 238576 140490 238628 140496
rect 239600 140418 239628 141335
rect 239678 140720 239734 140729
rect 239678 140655 239734 140664
rect 239692 140486 239720 140655
rect 239680 140480 239732 140486
rect 239680 140422 239732 140428
rect 239588 140412 239640 140418
rect 239588 140354 239640 140360
rect 238208 139392 238260 139398
rect 238208 139334 238260 139340
rect 238760 138848 238812 138854
rect 238760 138790 238812 138796
rect 238772 138281 238800 138790
rect 238758 138272 238814 138281
rect 238758 138207 238814 138216
rect 239784 138014 239812 178395
rect 239862 177372 239918 177381
rect 239862 177307 239918 177316
rect 237852 137986 238064 138014
rect 237380 137964 237432 137970
rect 237380 137906 237432 137912
rect 233148 137692 233200 137698
rect 233148 137634 233200 137640
rect 233160 137057 233188 137634
rect 233146 137048 233202 137057
rect 233146 136983 233202 136992
rect 237392 136921 237420 137906
rect 237378 136912 237434 136921
rect 237378 136847 237434 136856
rect 233422 133376 233478 133385
rect 233422 133311 233478 133320
rect 231122 28384 231178 28393
rect 231122 28319 231178 28328
rect 229834 3768 229890 3777
rect 229834 3703 229890 3712
rect 229848 480 229876 3703
rect 233436 480 233464 133311
rect 238036 112441 238064 137986
rect 239692 137986 239812 138014
rect 239692 135969 239720 137986
rect 239678 135960 239734 135969
rect 239678 135895 239734 135904
rect 238022 112432 238078 112441
rect 238022 112367 238078 112376
rect 239876 33153 239904 177307
rect 266910 140584 266966 140593
rect 266910 140519 266966 140528
rect 275282 140584 275338 140593
rect 275282 140519 275338 140528
rect 240782 139632 240838 139641
rect 240782 139567 240838 139576
rect 240796 139330 240824 139567
rect 240784 139324 240836 139330
rect 240784 139266 240836 139272
rect 239862 33144 239918 33153
rect 239862 33079 239918 33088
rect 241440 4865 241468 140148
rect 242636 6225 242664 140148
rect 243832 137630 243860 140148
rect 245028 137902 245056 140148
rect 245016 137896 245068 137902
rect 245016 137838 245068 137844
rect 246224 137834 246252 140148
rect 247040 137896 247092 137902
rect 247040 137838 247092 137844
rect 246212 137828 246264 137834
rect 246212 137770 246264 137776
rect 243820 137624 243872 137630
rect 243820 137566 243872 137572
rect 247052 136785 247080 137838
rect 247420 137766 247448 140148
rect 247408 137760 247460 137766
rect 247408 137702 247460 137708
rect 248616 137698 248644 140148
rect 249812 137970 249840 140148
rect 249800 137964 249852 137970
rect 249800 137906 249852 137912
rect 251008 137902 251036 140148
rect 251180 138576 251232 138582
rect 251180 138518 251232 138524
rect 250996 137896 251048 137902
rect 250996 137838 251048 137844
rect 248604 137692 248656 137698
rect 248604 137634 248656 137640
rect 247590 137184 247646 137193
rect 247590 137119 247646 137128
rect 247038 136776 247094 136785
rect 247038 136711 247094 136720
rect 244094 136368 244150 136377
rect 244094 136303 244150 136312
rect 242622 6216 242678 6225
rect 242622 6151 242678 6160
rect 241426 4856 241482 4865
rect 241426 4791 241482 4800
rect 241428 4140 241480 4146
rect 241428 4082 241480 4088
rect 237010 3904 237066 3913
rect 237010 3839 237066 3848
rect 237024 480 237052 3839
rect 240506 3224 240562 3233
rect 240506 3159 240562 3168
rect 240520 480 240548 3159
rect 241440 2825 241468 4082
rect 241426 2816 241482 2825
rect 241426 2751 241482 2760
rect 244108 480 244136 136303
rect 246302 134872 246358 134881
rect 246302 134807 246358 134816
rect 246316 3233 246344 134807
rect 246302 3224 246358 3233
rect 246302 3159 246358 3168
rect 247604 480 247632 137119
rect 251192 480 251220 138518
rect 252204 137329 252232 140148
rect 252190 137320 252246 137329
rect 252190 137255 252246 137264
rect 253400 6361 253428 140148
rect 254596 38185 254624 140148
rect 254674 137320 254730 137329
rect 254674 137255 254730 137264
rect 254582 38176 254638 38185
rect 254582 38111 254638 38120
rect 253386 6352 253442 6361
rect 253386 6287 253442 6296
rect 254688 480 254716 137255
rect 255792 21593 255820 140148
rect 256988 25673 257016 140148
rect 256974 25664 257030 25673
rect 256974 25599 257030 25608
rect 258184 22817 258212 140148
rect 258722 69456 258778 69465
rect 258722 69391 258778 69400
rect 258170 22808 258226 22817
rect 258170 22743 258226 22752
rect 255778 21584 255834 21593
rect 255778 21519 255834 21528
rect 258736 6225 258764 69391
rect 259380 36689 259408 140148
rect 260102 54496 260158 54505
rect 260102 54431 260158 54440
rect 259366 36680 259422 36689
rect 259366 36615 259422 36624
rect 258722 6216 258778 6225
rect 258722 6151 258778 6160
rect 260116 4865 260144 54431
rect 260576 33969 260604 140148
rect 261772 137986 261800 140148
rect 261680 137958 261800 137986
rect 262126 138000 262182 138009
rect 262310 138000 262366 138009
rect 260562 33960 260618 33969
rect 260562 33895 260618 33904
rect 261680 6497 261708 137958
rect 262126 137935 262128 137944
rect 262180 137935 262182 137944
rect 262232 137958 262310 137986
rect 262128 137906 262180 137912
rect 262232 137850 262260 137958
rect 262310 137935 262366 137944
rect 261772 137822 262260 137850
rect 261666 6488 261722 6497
rect 261666 6423 261722 6432
rect 260102 4856 260158 4865
rect 260102 4791 260158 4800
rect 258262 3224 258318 3233
rect 258262 3159 258318 3168
rect 258276 480 258304 3159
rect 261772 480 261800 137822
rect 262968 6633 262996 140148
rect 264164 6769 264192 140148
rect 265360 35329 265388 140148
rect 266556 93129 266584 140148
rect 266924 140010 266952 140519
rect 266912 140004 266964 140010
rect 266912 139946 266964 139952
rect 267002 139632 267058 139641
rect 267002 139567 267058 139576
rect 266542 93120 266598 93129
rect 266542 93055 266598 93064
rect 265346 35320 265402 35329
rect 265346 35255 265402 35264
rect 264150 6760 264206 6769
rect 264150 6695 264206 6704
rect 262954 6624 263010 6633
rect 262954 6559 263010 6568
rect 264980 4072 265032 4078
rect 264980 4014 265032 4020
rect 264992 2961 265020 4014
rect 267016 3233 267044 139567
rect 267752 108361 267780 140148
rect 268948 118017 268976 140148
rect 268934 118008 268990 118017
rect 268934 117943 268990 117952
rect 267738 108352 267794 108361
rect 267738 108287 267794 108296
rect 270144 106865 270172 140148
rect 271144 136672 271196 136678
rect 271144 136614 271196 136620
rect 270130 106856 270186 106865
rect 270130 106791 270186 106800
rect 271156 105505 271184 136614
rect 271142 105496 271198 105505
rect 271142 105431 271198 105440
rect 271340 94489 271368 140148
rect 272536 136678 272564 140148
rect 272524 136672 272576 136678
rect 272524 136614 272576 136620
rect 273732 95849 273760 140148
rect 274928 97345 274956 140148
rect 274914 97336 274970 97345
rect 274914 97271 274970 97280
rect 273718 95840 273774 95849
rect 273718 95775 273774 95784
rect 271326 94480 271382 94489
rect 271326 94415 271382 94424
rect 273902 85912 273958 85921
rect 273902 85847 273958 85856
rect 271142 85776 271198 85785
rect 271142 85711 271198 85720
rect 267186 46336 267242 46345
rect 267186 46271 267242 46280
rect 267200 4049 267228 46271
rect 267186 4040 267242 4049
rect 267186 3975 267242 3984
rect 268842 4040 268898 4049
rect 268842 3975 268898 3984
rect 267002 3224 267058 3233
rect 267002 3159 267058 3168
rect 265346 3088 265402 3097
rect 265346 3023 265402 3032
rect 264978 2952 265034 2961
rect 264978 2887 265034 2896
rect 265360 480 265388 3023
rect 268856 480 268884 3975
rect 271156 3233 271184 85711
rect 273916 3233 273944 85847
rect 271142 3224 271198 3233
rect 271142 3159 271198 3168
rect 272430 3224 272486 3233
rect 272430 3159 272486 3168
rect 273902 3224 273958 3233
rect 273902 3159 273958 3168
rect 272444 480 272472 3159
rect 275296 3097 275324 140519
rect 276124 137465 276152 140148
rect 277320 137601 277348 140148
rect 277306 137592 277362 137601
rect 277306 137527 277362 137536
rect 276110 137456 276166 137465
rect 276110 137391 276166 137400
rect 278516 104281 278544 140148
rect 278502 104272 278558 104281
rect 278502 104207 278558 104216
rect 280080 102785 280108 201447
rect 280172 137329 280200 237351
rect 280342 236056 280398 236065
rect 280342 235991 280398 236000
rect 280250 234696 280306 234705
rect 280250 234631 280306 234640
rect 280158 137320 280214 137329
rect 280158 137255 280214 137264
rect 280264 136377 280292 234631
rect 280356 138582 280384 235991
rect 280526 225040 280582 225049
rect 280526 224975 280582 224984
rect 280434 222864 280490 222873
rect 280434 222799 280490 222808
rect 280344 138576 280396 138582
rect 280344 138518 280396 138524
rect 280250 136368 280306 136377
rect 280250 136303 280306 136312
rect 280448 134745 280476 222799
rect 280540 140049 280568 224975
rect 280802 216744 280858 216753
rect 280802 216679 280858 216688
rect 280618 213208 280674 213217
rect 280618 213143 280674 213152
rect 280526 140040 280582 140049
rect 280526 139975 280582 139984
rect 280434 134736 280490 134745
rect 280434 134671 280490 134680
rect 280632 129169 280660 213143
rect 280618 129160 280674 129169
rect 280618 129095 280674 129104
rect 280066 102776 280122 102785
rect 280066 102711 280122 102720
rect 278042 32464 278098 32473
rect 278042 32399 278098 32408
rect 277858 4040 277914 4049
rect 277858 3975 277914 3984
rect 277872 3505 277900 3975
rect 278056 3505 278084 32399
rect 280816 3777 280844 216679
rect 280986 205728 281042 205737
rect 280986 205663 281042 205672
rect 281000 3913 281028 205663
rect 281170 204232 281226 204241
rect 281170 204167 281226 204176
rect 280986 3904 281042 3913
rect 280986 3839 281042 3848
rect 280802 3768 280858 3777
rect 280802 3703 280858 3712
rect 281184 3641 281212 204167
rect 281354 196072 281410 196081
rect 281354 196007 281410 196016
rect 281368 4049 281396 196007
rect 281552 140593 281580 239255
rect 281814 237688 281870 237697
rect 281814 237623 281870 237632
rect 281722 235240 281778 235249
rect 281722 235175 281778 235184
rect 281630 233608 281686 233617
rect 281630 233543 281686 233552
rect 281538 140584 281594 140593
rect 281538 140519 281594 140528
rect 281644 134881 281672 233543
rect 281736 137193 281764 235175
rect 281828 139641 281856 237623
rect 281998 233336 282054 233345
rect 281998 233271 282054 233280
rect 281906 231160 281962 231169
rect 281906 231095 281962 231104
rect 281920 216753 281948 231095
rect 281906 216744 281962 216753
rect 281906 216679 281962 216688
rect 281906 212664 281962 212673
rect 281906 212599 281962 212608
rect 281814 139632 281870 139641
rect 281814 139567 281870 139576
rect 281722 137184 281778 137193
rect 281722 137119 281778 137128
rect 281630 134872 281686 134881
rect 281630 134807 281686 134816
rect 281920 116657 281948 212599
rect 282012 205737 282040 233271
rect 282182 229256 282238 229265
rect 282182 229191 282238 229200
rect 282196 229158 282224 229191
rect 282184 229152 282236 229158
rect 282184 229094 282236 229100
rect 282274 227896 282330 227905
rect 282274 227831 282330 227840
rect 282288 227798 282316 227831
rect 282276 227792 282328 227798
rect 282276 227734 282328 227740
rect 282090 225312 282146 225321
rect 282090 225247 282146 225256
rect 281998 205728 282054 205737
rect 281998 205663 282054 205672
rect 281998 203280 282054 203289
rect 281998 203215 282054 203224
rect 281906 116648 281962 116657
rect 281906 116583 281962 116592
rect 282012 108497 282040 203215
rect 282104 138650 282132 225247
rect 282182 220960 282238 220969
rect 282182 220895 282238 220904
rect 282196 139126 282224 220895
rect 282458 219872 282514 219881
rect 282458 219807 282514 219816
rect 282366 218104 282422 218113
rect 282366 218039 282422 218048
rect 282380 196081 282408 218039
rect 282472 204241 282500 219807
rect 282828 219496 282880 219502
rect 282826 219464 282828 219473
rect 282880 219464 282882 219473
rect 282826 219399 282882 219408
rect 282826 211712 282882 211721
rect 282826 211647 282882 211656
rect 282840 211206 282868 211647
rect 282828 211200 282880 211206
rect 282828 211142 282880 211148
rect 282826 204912 282882 204921
rect 282826 204847 282882 204856
rect 282840 204338 282868 204847
rect 282828 204332 282880 204338
rect 282828 204274 282880 204280
rect 282458 204232 282514 204241
rect 282458 204167 282514 204176
rect 282366 196072 282422 196081
rect 282366 196007 282422 196016
rect 282274 193352 282330 193361
rect 282274 193287 282330 193296
rect 282184 139120 282236 139126
rect 282184 139062 282236 139068
rect 282092 138644 282144 138650
rect 282092 138586 282144 138592
rect 282288 133249 282316 193287
rect 282366 190632 282422 190641
rect 282366 190567 282422 190576
rect 282380 171714 282408 190567
rect 282458 178120 282514 178129
rect 282458 178055 282460 178064
rect 282512 178055 282514 178064
rect 282460 178026 282512 178032
rect 282826 176896 282882 176905
rect 282826 176831 282882 176840
rect 282840 176730 282868 176831
rect 282828 176724 282880 176730
rect 282828 176666 282880 176672
rect 282932 173641 282960 376071
rect 284312 361049 284340 390116
rect 284298 361040 284354 361049
rect 284298 360975 284354 360984
rect 287704 351212 287756 351218
rect 287704 351154 287756 351160
rect 284300 344004 284352 344010
rect 284300 343946 284352 343952
rect 283196 343868 283248 343874
rect 283196 343810 283248 343816
rect 283104 342984 283156 342990
rect 283104 342926 283156 342932
rect 283012 342712 283064 342718
rect 283012 342654 283064 342660
rect 283024 255105 283052 342654
rect 283116 267345 283144 342926
rect 283208 270473 283236 343810
rect 283288 343052 283340 343058
rect 283288 342994 283340 343000
rect 283194 270464 283250 270473
rect 283194 270399 283250 270408
rect 283300 268977 283328 342994
rect 283564 342440 283616 342446
rect 283564 342382 283616 342388
rect 283472 341216 283524 341222
rect 283472 341158 283524 341164
rect 283380 339720 283432 339726
rect 283380 339662 283432 339668
rect 283392 280129 283420 339662
rect 283484 282713 283512 341158
rect 283576 283665 283604 342382
rect 283656 339652 283708 339658
rect 283656 339594 283708 339600
rect 283562 283656 283618 283665
rect 283562 283591 283618 283600
rect 283470 282704 283526 282713
rect 283470 282639 283526 282648
rect 283668 281081 283696 339594
rect 283748 339584 283800 339590
rect 283748 339526 283800 339532
rect 283760 285666 283788 339526
rect 283748 285660 283800 285666
rect 283748 285602 283800 285608
rect 283654 281072 283710 281081
rect 283654 281007 283710 281016
rect 283378 280120 283434 280129
rect 283378 280055 283434 280064
rect 283286 268968 283342 268977
rect 283286 268903 283342 268912
rect 283102 267336 283158 267345
rect 283102 267271 283158 267280
rect 284312 266354 284340 343946
rect 287520 343800 287572 343806
rect 287520 343742 287572 343748
rect 285956 343732 286008 343738
rect 285956 343674 286008 343680
rect 284392 343120 284444 343126
rect 284392 343062 284444 343068
rect 284404 267714 284432 343062
rect 284484 342916 284536 342922
rect 284484 342858 284536 342864
rect 284496 270502 284524 342858
rect 285680 342848 285732 342854
rect 285680 342790 285732 342796
rect 284944 342576 284996 342582
rect 284944 342518 284996 342524
rect 284852 342508 284904 342514
rect 284852 342450 284904 342456
rect 284760 341352 284812 341358
rect 284760 341294 284812 341300
rect 284576 341284 284628 341290
rect 284576 341226 284628 341232
rect 284588 281518 284616 341226
rect 284668 339856 284720 339862
rect 284668 339798 284720 339804
rect 284576 281512 284628 281518
rect 284576 281454 284628 281460
rect 284680 280158 284708 339798
rect 284772 284306 284800 341294
rect 284864 288386 284892 342450
rect 284956 289814 284984 342518
rect 285036 339992 285088 339998
rect 285036 339934 285088 339940
rect 285048 299470 285076 339934
rect 285036 299464 285088 299470
rect 285036 299406 285088 299412
rect 284944 289808 284996 289814
rect 284944 289750 284996 289756
rect 284852 288380 284904 288386
rect 284852 288322 284904 288328
rect 284760 284300 284812 284306
rect 284760 284242 284812 284248
rect 284668 280152 284720 280158
rect 284668 280094 284720 280100
rect 284484 270496 284536 270502
rect 284484 270438 284536 270444
rect 284392 267708 284444 267714
rect 284392 267650 284444 267656
rect 284300 266348 284352 266354
rect 284300 266290 284352 266296
rect 285692 260846 285720 342790
rect 285864 342304 285916 342310
rect 285864 342246 285916 342252
rect 285772 339924 285824 339930
rect 285772 339866 285824 339872
rect 285680 260840 285732 260846
rect 285680 260782 285732 260788
rect 285784 257514 285812 339866
rect 285876 285598 285904 342246
rect 285968 286754 285996 343674
rect 286048 343664 286100 343670
rect 286048 343606 286100 343612
rect 286060 288318 286088 343606
rect 287428 342372 287480 342378
rect 287428 342314 287480 342320
rect 287060 341692 287112 341698
rect 287060 341634 287112 341640
rect 286048 288312 286100 288318
rect 286048 288254 286100 288260
rect 285956 286748 286008 286754
rect 285956 286690 286008 286696
rect 285864 285592 285916 285598
rect 285864 285534 285916 285540
rect 285772 257508 285824 257514
rect 285772 257450 285824 257456
rect 283010 255096 283066 255105
rect 283010 255031 283066 255040
rect 285862 238912 285918 238921
rect 285862 238847 285918 238856
rect 283102 230616 283158 230625
rect 283102 230551 283158 230560
rect 283010 191040 283066 191049
rect 283010 190975 283066 190984
rect 282918 173632 282974 173641
rect 282918 173567 282974 173576
rect 282828 172508 282880 172514
rect 282828 172450 282880 172456
rect 282736 172440 282788 172446
rect 282736 172382 282788 172388
rect 282748 171873 282776 172382
rect 282840 172281 282868 172450
rect 282826 172272 282882 172281
rect 282826 172207 282882 172216
rect 282734 171864 282790 171873
rect 282734 171799 282790 171808
rect 282380 171686 282960 171714
rect 282828 171080 282880 171086
rect 282828 171022 282880 171028
rect 282840 170785 282868 171022
rect 282826 170776 282882 170785
rect 282826 170711 282882 170720
rect 282828 169720 282880 169726
rect 282826 169688 282828 169697
rect 282880 169688 282882 169697
rect 282826 169623 282882 169632
rect 282828 169584 282880 169590
rect 282828 169526 282880 169532
rect 282840 169289 282868 169526
rect 282826 169280 282882 169289
rect 282826 169215 282882 169224
rect 282736 168360 282788 168366
rect 282736 168302 282788 168308
rect 282748 167793 282776 168302
rect 282828 168292 282880 168298
rect 282828 168234 282880 168240
rect 282840 168201 282868 168234
rect 282826 168192 282882 168201
rect 282826 168127 282882 168136
rect 282734 167784 282790 167793
rect 282734 167719 282790 167728
rect 282274 133240 282330 133249
rect 282274 133175 282330 133184
rect 281998 108488 282054 108497
rect 281998 108423 282054 108432
rect 282182 43616 282238 43625
rect 282182 43551 282238 43560
rect 281354 4040 281410 4049
rect 281354 3975 281410 3984
rect 281170 3632 281226 3641
rect 281170 3567 281226 3576
rect 282196 3505 282224 43551
rect 282932 4146 282960 171686
rect 283024 14793 283052 190975
rect 283116 123593 283144 230551
rect 284482 229528 284538 229537
rect 284482 229463 284538 229472
rect 283286 222320 283342 222329
rect 283286 222255 283342 222264
rect 283194 214024 283250 214033
rect 283194 213959 283250 213968
rect 283102 123584 283158 123593
rect 283102 123519 283158 123528
rect 283208 111081 283236 213959
rect 283300 129305 283328 222255
rect 283378 221368 283434 221377
rect 283378 221303 283434 221312
rect 283392 138922 283420 221303
rect 283470 216744 283526 216753
rect 283470 216679 283526 216688
rect 283380 138916 283432 138922
rect 283380 138858 283432 138864
rect 283484 136241 283512 216679
rect 283562 215656 283618 215665
rect 283562 215591 283618 215600
rect 283470 136232 283526 136241
rect 283470 136167 283526 136176
rect 283576 136105 283604 215591
rect 284390 215384 284446 215393
rect 284390 215319 284446 215328
rect 283654 207496 283710 207505
rect 283654 207431 283710 207440
rect 283562 136096 283618 136105
rect 283562 136031 283618 136040
rect 283668 134609 283696 207431
rect 284298 193624 284354 193633
rect 284298 193559 284354 193568
rect 283748 178084 283800 178090
rect 283748 178026 283800 178032
rect 283760 140010 283788 178026
rect 283748 140004 283800 140010
rect 283748 139946 283800 139952
rect 283654 134600 283710 134609
rect 283654 134535 283710 134544
rect 283286 129296 283342 129305
rect 283286 129231 283342 129240
rect 283194 111072 283250 111081
rect 283194 111007 283250 111016
rect 284312 50289 284340 193559
rect 284404 109721 284432 215319
rect 284496 124953 284524 229463
rect 284944 229152 284996 229158
rect 284944 229094 284996 229100
rect 284666 227080 284722 227089
rect 284666 227015 284722 227024
rect 284574 203008 284630 203017
rect 284574 202943 284630 202952
rect 284482 124944 284538 124953
rect 284482 124879 284538 124888
rect 284390 109712 284446 109721
rect 284390 109647 284446 109656
rect 284588 98841 284616 202943
rect 284680 126449 284708 227015
rect 284758 226400 284814 226409
rect 284758 226335 284814 226344
rect 284772 132025 284800 226335
rect 284850 223680 284906 223689
rect 284850 223615 284906 223624
rect 284758 132016 284814 132025
rect 284758 131951 284814 131960
rect 284864 131889 284892 223615
rect 284956 138718 284984 229094
rect 285128 227792 285180 227798
rect 285128 227734 285180 227740
rect 285034 208992 285090 209001
rect 285034 208927 285090 208936
rect 284944 138712 284996 138718
rect 284944 138654 284996 138660
rect 284850 131880 284906 131889
rect 284850 131815 284906 131824
rect 284666 126440 284722 126449
rect 284666 126375 284722 126384
rect 285048 119513 285076 208927
rect 285140 138786 285168 227734
rect 285770 197432 285826 197441
rect 285770 197367 285826 197376
rect 285678 196072 285734 196081
rect 285678 196007 285734 196016
rect 285128 138780 285180 138786
rect 285128 138722 285180 138728
rect 285034 119504 285090 119513
rect 285034 119439 285090 119448
rect 284574 98832 284630 98841
rect 284574 98767 284630 98776
rect 284298 50280 284354 50289
rect 284298 50215 284354 50224
rect 285692 21457 285720 196007
rect 285784 32609 285812 197367
rect 285876 138009 285904 238847
rect 285954 231976 286010 231985
rect 285954 231911 286010 231920
rect 285862 138000 285918 138009
rect 285862 137935 285918 137944
rect 285968 133385 285996 231911
rect 286046 204368 286102 204377
rect 286046 204303 286102 204312
rect 285954 133376 286010 133385
rect 285954 133311 286010 133320
rect 286060 123457 286088 204303
rect 286322 201784 286378 201793
rect 286322 201719 286378 201728
rect 286138 200424 286194 200433
rect 286138 200359 286194 200368
rect 286046 123448 286102 123457
rect 286046 123383 286102 123392
rect 286152 119377 286180 200359
rect 286230 199336 286286 199345
rect 286230 199271 286286 199280
rect 286244 124817 286272 199271
rect 286336 131753 286364 201719
rect 286414 198792 286470 198801
rect 286414 198727 286470 198736
rect 286322 131744 286378 131753
rect 286322 131679 286378 131688
rect 286428 130393 286456 198727
rect 286506 197704 286562 197713
rect 286506 197639 286562 197648
rect 286414 130384 286470 130393
rect 286414 130319 286470 130328
rect 286520 129033 286548 197639
rect 287072 169590 287100 341634
rect 287152 274712 287204 274718
rect 287152 274654 287204 274660
rect 287060 169584 287112 169590
rect 287060 169526 287112 169532
rect 287164 138990 287192 274654
rect 287244 273352 287296 273358
rect 287244 273294 287296 273300
rect 287256 140146 287284 273294
rect 287336 271924 287388 271930
rect 287336 271866 287388 271872
rect 287244 140140 287296 140146
rect 287244 140082 287296 140088
rect 287348 140078 287376 271866
rect 287440 253910 287468 342314
rect 287532 256698 287560 343742
rect 287612 342780 287664 342786
rect 287612 342722 287664 342728
rect 287624 262206 287652 342722
rect 287612 262200 287664 262206
rect 287612 262142 287664 262148
rect 287520 256692 287572 256698
rect 287520 256634 287572 256640
rect 287428 253904 287480 253910
rect 287428 253846 287480 253852
rect 287518 207224 287574 207233
rect 287518 207159 287574 207168
rect 287426 206408 287482 206417
rect 287426 206343 287482 206352
rect 287336 140072 287388 140078
rect 287336 140014 287388 140020
rect 287152 138984 287204 138990
rect 287152 138926 287204 138932
rect 286506 129024 286562 129033
rect 286506 128959 286562 128968
rect 286230 124808 286286 124817
rect 286230 124743 286286 124752
rect 286138 119368 286194 119377
rect 286138 119303 286194 119312
rect 287440 90409 287468 206343
rect 287532 100201 287560 207159
rect 287716 187746 287744 351154
rect 287900 340377 287928 390116
rect 288532 345704 288584 345710
rect 288532 345646 288584 345652
rect 287886 340368 287942 340377
rect 287886 340303 287942 340312
rect 288438 217832 288494 217841
rect 288438 217767 288494 217776
rect 287794 188456 287850 188465
rect 287794 188391 287850 188400
rect 287704 187740 287756 187746
rect 287704 187682 287756 187688
rect 287610 187640 287666 187649
rect 287610 187575 287666 187584
rect 287624 104145 287652 187575
rect 287702 186824 287758 186833
rect 287702 186759 287758 186768
rect 287716 120737 287744 186759
rect 287808 122097 287836 188391
rect 287886 186008 287942 186017
rect 287886 185943 287942 185952
rect 287794 122088 287850 122097
rect 287794 122023 287850 122032
rect 287702 120728 287758 120737
rect 287702 120663 287758 120672
rect 287610 104136 287666 104145
rect 287610 104071 287666 104080
rect 287900 101425 287928 185943
rect 287886 101416 287942 101425
rect 287886 101351 287942 101360
rect 287518 100192 287574 100201
rect 287518 100127 287574 100136
rect 287426 90400 287482 90409
rect 287426 90335 287482 90344
rect 287704 87100 287756 87106
rect 287704 87042 287756 87048
rect 285770 32600 285826 32609
rect 285770 32535 285826 32544
rect 285678 21448 285734 21457
rect 285678 21383 285734 21392
rect 283010 14784 283066 14793
rect 283010 14719 283066 14728
rect 286598 6216 286654 6225
rect 286598 6151 286654 6160
rect 283102 4856 283158 4865
rect 283102 4791 283158 4800
rect 282920 4140 282972 4146
rect 282920 4082 282972 4088
rect 277858 3496 277914 3505
rect 277858 3431 277914 3440
rect 278042 3496 278098 3505
rect 278042 3431 278098 3440
rect 279514 3496 279570 3505
rect 279514 3431 279570 3440
rect 282182 3496 282238 3505
rect 282182 3431 282238 3440
rect 276018 3224 276074 3233
rect 276018 3159 276074 3168
rect 275282 3088 275338 3097
rect 275282 3023 275338 3032
rect 276032 480 276060 3159
rect 279528 480 279556 3431
rect 283116 480 283144 4791
rect 286612 480 286640 6151
rect 287716 4826 287744 87042
rect 287704 4820 287756 4826
rect 287704 4762 287756 4768
rect 288452 3369 288480 217767
rect 288544 168298 288572 345646
rect 291384 341148 291436 341154
rect 291384 341090 291436 341096
rect 291292 341080 291344 341086
rect 291292 341022 291344 341028
rect 288624 277500 288676 277506
rect 288624 277442 288676 277448
rect 288532 168292 288584 168298
rect 288532 168234 288584 168240
rect 288636 137970 288664 277442
rect 288716 276140 288768 276146
rect 288716 276082 288768 276088
rect 288728 139058 288756 276082
rect 289912 276072 289964 276078
rect 289912 276014 289964 276020
rect 288806 274952 288862 274961
rect 288806 274887 288862 274896
rect 288820 140321 288848 274887
rect 288900 242956 288952 242962
rect 288900 242898 288952 242904
rect 288806 140312 288862 140321
rect 288806 140247 288862 140256
rect 288716 139052 288768 139058
rect 288716 138994 288768 139000
rect 288912 138854 288940 242898
rect 288992 211200 289044 211206
rect 288992 211142 289044 211148
rect 289004 139262 289032 211142
rect 289818 190088 289874 190097
rect 289818 190023 289874 190032
rect 289082 181112 289138 181121
rect 289082 181047 289138 181056
rect 289096 139505 289124 181047
rect 289176 176724 289228 176730
rect 289176 176666 289228 176672
rect 289188 140214 289216 176666
rect 289176 140208 289228 140214
rect 289176 140150 289228 140156
rect 289082 139496 289138 139505
rect 289082 139431 289138 139440
rect 288992 139256 289044 139262
rect 288992 139198 289044 139204
rect 288900 138848 288952 138854
rect 288900 138790 288952 138796
rect 288624 137964 288676 137970
rect 288624 137906 288676 137912
rect 289832 49201 289860 190023
rect 289924 141681 289952 276014
rect 290004 273284 290056 273290
rect 290004 273226 290056 273232
rect 290016 141817 290044 273226
rect 290094 250336 290150 250345
rect 290094 250271 290150 250280
rect 290002 141808 290058 141817
rect 290002 141743 290058 141752
rect 289910 141672 289966 141681
rect 289910 141607 289966 141616
rect 290108 138417 290136 250271
rect 290186 249520 290242 249529
rect 290186 249455 290242 249464
rect 290200 139233 290228 249455
rect 290278 247888 290334 247897
rect 290278 247823 290334 247832
rect 290292 141409 290320 247823
rect 290370 240680 290426 240689
rect 290370 240615 290426 240624
rect 290278 141400 290334 141409
rect 290278 141335 290334 141344
rect 290384 139913 290412 240615
rect 290464 219496 290516 219502
rect 290464 219438 290516 219444
rect 290370 139904 290426 139913
rect 290370 139839 290426 139848
rect 290186 139224 290242 139233
rect 290476 139194 290504 219438
rect 291200 187740 291252 187746
rect 291200 187682 291252 187688
rect 291212 168366 291240 187682
rect 291304 169726 291332 341022
rect 291396 172446 291424 341090
rect 291488 340241 291516 390116
rect 295076 362545 295104 390116
rect 295062 362536 295118 362545
rect 295062 362471 295118 362480
rect 291844 341420 291896 341426
rect 291844 341362 291896 341368
rect 291474 340232 291530 340241
rect 291474 340167 291530 340176
rect 291568 270632 291620 270638
rect 291568 270574 291620 270580
rect 291476 270564 291528 270570
rect 291476 270506 291528 270512
rect 291384 172440 291436 172446
rect 291384 172382 291436 172388
rect 291292 169720 291344 169726
rect 291292 169662 291344 169668
rect 291200 168360 291252 168366
rect 291200 168302 291252 168308
rect 291488 140282 291516 270506
rect 291580 140350 291608 270574
rect 291658 247072 291714 247081
rect 291658 247007 291714 247016
rect 291568 140344 291620 140350
rect 291568 140286 291620 140292
rect 291476 140276 291528 140282
rect 291476 140218 291528 140224
rect 291672 140185 291700 247007
rect 291752 204332 291804 204338
rect 291752 204274 291804 204280
rect 291658 140176 291714 140185
rect 291658 140111 291714 140120
rect 290186 139159 290242 139168
rect 290464 139188 290516 139194
rect 290464 139130 290516 139136
rect 290094 138408 290150 138417
rect 290094 138343 290150 138352
rect 289818 49192 289874 49201
rect 289818 49127 289874 49136
rect 289082 49056 289138 49065
rect 289082 48991 289138 49000
rect 289096 3369 289124 48991
rect 290186 9072 290242 9081
rect 290186 9007 290242 9016
rect 288438 3360 288494 3369
rect 288438 3295 288494 3304
rect 289082 3360 289138 3369
rect 289082 3295 289138 3304
rect 290200 480 290228 9007
rect 291764 4078 291792 204274
rect 291856 6866 291884 341362
rect 295340 341012 295392 341018
rect 295340 340954 295392 340960
rect 292580 340944 292632 340950
rect 292580 340886 292632 340892
rect 292592 171086 292620 340886
rect 292670 251288 292726 251297
rect 292670 251223 292726 251232
rect 292580 171080 292632 171086
rect 292580 171022 292632 171028
rect 292684 141953 292712 251223
rect 295352 172514 295380 340954
rect 298664 340105 298692 390116
rect 302252 345953 302280 390116
rect 305840 382809 305868 390116
rect 305826 382800 305882 382809
rect 305826 382735 305882 382744
rect 309428 356969 309456 390116
rect 309414 356960 309470 356969
rect 309414 356895 309470 356904
rect 313016 352617 313044 390116
rect 313002 352608 313058 352617
rect 313002 352543 313058 352552
rect 316604 351393 316632 390116
rect 320192 355473 320220 390116
rect 320178 355464 320234 355473
rect 320178 355399 320234 355408
rect 316590 351384 316646 351393
rect 316590 351319 316646 351328
rect 302238 345944 302294 345953
rect 302238 345879 302294 345888
rect 323780 345001 323808 390116
rect 327368 358057 327396 390116
rect 327354 358048 327410 358057
rect 327354 357983 327410 357992
rect 323766 344992 323822 345001
rect 323766 344927 323822 344936
rect 330956 342825 330984 390116
rect 334544 386753 334572 390116
rect 334530 386744 334586 386753
rect 334530 386679 334586 386688
rect 330942 342816 330998 342825
rect 330942 342751 330998 342760
rect 338132 342553 338160 390116
rect 341720 386889 341748 390116
rect 341706 386880 341762 386889
rect 341706 386815 341762 386824
rect 345308 342689 345336 390116
rect 348896 387705 348924 390116
rect 348882 387696 348938 387705
rect 348882 387631 348938 387640
rect 352484 343369 352512 390116
rect 356072 387569 356100 390116
rect 356058 387560 356114 387569
rect 356058 387495 356114 387504
rect 359660 344865 359688 390116
rect 363248 367713 363276 390116
rect 366836 369345 366864 390116
rect 366822 369336 366878 369345
rect 366822 369271 366878 369280
rect 363234 367704 363290 367713
rect 363234 367639 363290 367648
rect 359646 344856 359702 344865
rect 359646 344791 359702 344800
rect 370424 344729 370452 390116
rect 370410 344720 370466 344729
rect 370410 344655 370466 344664
rect 374012 344593 374040 390116
rect 377600 381721 377628 390116
rect 377586 381712 377642 381721
rect 377586 381647 377642 381656
rect 381188 371929 381216 390116
rect 384776 377233 384804 390116
rect 384762 377224 384818 377233
rect 384762 377159 384818 377168
rect 388364 373425 388392 390116
rect 388350 373416 388406 373425
rect 388350 373351 388406 373360
rect 381174 371920 381230 371929
rect 381174 371855 381230 371864
rect 391952 359553 391980 390116
rect 392582 387152 392638 387161
rect 392582 387087 392638 387096
rect 391938 359544 391994 359553
rect 391938 359479 391994 359488
rect 373998 344584 374054 344593
rect 373998 344519 374054 344528
rect 352470 343360 352526 343369
rect 352470 343295 352526 343304
rect 392596 343233 392624 387087
rect 395540 370705 395568 390116
rect 395526 370696 395582 370705
rect 395526 370631 395582 370640
rect 399128 344457 399156 390116
rect 402716 366353 402744 390116
rect 402702 366344 402758 366353
rect 402702 366279 402758 366288
rect 406304 360913 406332 390116
rect 409892 365129 409920 390116
rect 409878 365120 409934 365129
rect 409878 365055 409934 365064
rect 406290 360904 406346 360913
rect 406290 360839 406346 360848
rect 410524 347064 410576 347070
rect 410524 347006 410576 347012
rect 410536 345030 410564 347006
rect 410524 345024 410576 345030
rect 410524 344966 410576 344972
rect 399114 344448 399170 344457
rect 399114 344383 399170 344392
rect 413480 344321 413508 390116
rect 417068 378865 417096 390116
rect 417422 387560 417478 387569
rect 417422 387495 417478 387504
rect 417054 378856 417110 378865
rect 417054 378791 417110 378800
rect 413466 344312 413522 344321
rect 413466 344247 413522 344256
rect 392582 343224 392638 343233
rect 392582 343159 392638 343168
rect 417436 343097 417464 387495
rect 420656 387433 420684 390116
rect 420642 387424 420698 387433
rect 420642 387359 420698 387368
rect 424244 376281 424272 390116
rect 424230 376272 424286 376281
rect 424230 376207 424286 376216
rect 426348 369980 426400 369986
rect 426348 369922 426400 369928
rect 426360 367810 426388 369922
rect 420184 367804 420236 367810
rect 420184 367746 420236 367752
rect 426348 367804 426400 367810
rect 426348 367746 426400 367752
rect 420196 358766 420224 367746
rect 427832 362409 427860 390116
rect 431420 387297 431448 390116
rect 431406 387288 431462 387297
rect 431406 387223 431462 387232
rect 427912 373312 427964 373318
rect 427912 373254 427964 373260
rect 427924 369986 427952 373254
rect 427912 369980 427964 369986
rect 427912 369922 427964 369928
rect 427818 362400 427874 362409
rect 427818 362335 427874 362344
rect 417516 358760 417568 358766
rect 417516 358702 417568 358708
rect 420184 358760 420236 358766
rect 420184 358702 420236 358708
rect 417528 347070 417556 358702
rect 435008 356833 435036 390116
rect 438596 387025 438624 390116
rect 442184 387161 442212 390116
rect 445772 387190 445800 390116
rect 449360 387569 449388 390116
rect 452948 387705 452976 390116
rect 452934 387696 452990 387705
rect 452934 387631 452990 387640
rect 449346 387560 449402 387569
rect 449346 387495 449402 387504
rect 445760 387184 445812 387190
rect 442170 387152 442226 387161
rect 445760 387126 445812 387132
rect 442170 387087 442226 387096
rect 438582 387016 438638 387025
rect 438582 386951 438638 386960
rect 452948 384305 452976 387631
rect 456536 386889 456564 390116
rect 460124 386918 460152 390116
rect 458824 386912 458876 386918
rect 454682 386880 454738 386889
rect 454682 386815 454738 386824
rect 456522 386880 456578 386889
rect 458824 386854 458876 386860
rect 460112 386912 460164 386918
rect 460112 386854 460164 386860
rect 456522 386815 456578 386824
rect 452934 384296 452990 384305
rect 452934 384231 452990 384240
rect 449900 382968 449952 382974
rect 449900 382910 449952 382916
rect 449912 376038 449940 382910
rect 438768 376032 438820 376038
rect 438768 375974 438820 375980
rect 449900 376032 449952 376038
rect 449900 375974 449952 375980
rect 438780 373318 438808 375974
rect 438768 373312 438820 373318
rect 438768 373254 438820 373260
rect 454696 363769 454724 386815
rect 454682 363760 454738 363769
rect 454682 363695 454738 363704
rect 434994 356824 435050 356833
rect 434994 356759 435050 356768
rect 458178 356008 458234 356017
rect 458178 355943 458234 355952
rect 458192 349874 458220 355943
rect 457456 349846 458220 349874
rect 456798 347712 456854 347721
rect 456798 347647 456854 347656
rect 417516 347064 417568 347070
rect 417516 347006 417568 347012
rect 417422 343088 417478 343097
rect 417422 343023 417478 343032
rect 345294 342680 345350 342689
rect 345294 342615 345350 342624
rect 338118 342544 338174 342553
rect 338118 342479 338174 342488
rect 298650 340096 298706 340105
rect 298650 340031 298706 340040
rect 456812 339425 456840 347647
rect 453302 339416 453358 339425
rect 453302 339351 453358 339360
rect 456798 339416 456854 339425
rect 456798 339351 456854 339360
rect 453316 332489 453344 339351
rect 447782 332480 447838 332489
rect 447782 332415 447838 332424
rect 453302 332480 453358 332489
rect 453302 332415 453358 332424
rect 447796 270473 447824 332415
rect 457456 327049 457484 349846
rect 456062 327040 456118 327049
rect 456062 326975 456118 326984
rect 457442 327040 457498 327049
rect 457442 326975 457498 326984
rect 456076 318753 456104 326975
rect 454682 318744 454738 318753
rect 454682 318679 454738 318688
rect 456062 318744 456118 318753
rect 456062 318679 456118 318688
rect 442262 270464 442318 270473
rect 442262 270399 442318 270408
rect 447782 270464 447838 270473
rect 447782 270399 447838 270408
rect 442276 238785 442304 270399
rect 454696 253201 454724 318679
rect 451922 253192 451978 253201
rect 451922 253127 451978 253136
rect 454682 253192 454738 253201
rect 454682 253127 454738 253136
rect 440882 238776 440938 238785
rect 440882 238711 440938 238720
rect 442262 238776 442318 238785
rect 442262 238711 442318 238720
rect 440896 231849 440924 238711
rect 439502 231840 439558 231849
rect 439502 231775 439558 231784
rect 440882 231840 440938 231849
rect 440882 231775 440938 231784
rect 439516 191729 439544 231775
rect 451936 224913 451964 253127
rect 450542 224904 450598 224913
rect 450542 224839 450598 224848
rect 451922 224904 451978 224913
rect 451922 224839 451978 224848
rect 450556 204241 450584 224839
rect 449162 204232 449218 204241
rect 449162 204167 449218 204176
rect 450542 204232 450598 204241
rect 450542 204167 450598 204176
rect 449176 198801 449204 204167
rect 445390 198792 445446 198801
rect 445390 198727 445446 198736
rect 449162 198792 449218 198801
rect 449162 198727 449218 198736
rect 445404 194857 445432 198727
rect 442906 194848 442962 194857
rect 442906 194783 442962 194792
rect 445390 194848 445446 194857
rect 445390 194783 445446 194792
rect 436006 191720 436062 191729
rect 436006 191655 436062 191664
rect 439502 191720 439558 191729
rect 439502 191655 439558 191664
rect 434626 187776 434682 187785
rect 434626 187711 434682 187720
rect 429198 185600 429254 185609
rect 429198 185535 429254 185544
rect 428462 184920 428518 184929
rect 428462 184855 428518 184864
rect 426438 183152 426494 183161
rect 426438 183087 426494 183096
rect 426452 176746 426480 183087
rect 428476 179489 428504 184855
rect 429212 183161 429240 185535
rect 434640 184929 434668 187711
rect 436020 185609 436048 191655
rect 442920 190505 442948 194783
rect 442906 190496 442962 190505
rect 442906 190431 442962 190440
rect 436098 190360 436154 190369
rect 436098 190295 436154 190304
rect 436112 187785 436140 190295
rect 436098 187776 436154 187785
rect 436098 187711 436154 187720
rect 436006 185600 436062 185609
rect 436006 185535 436062 185544
rect 434626 184920 434682 184929
rect 434626 184855 434682 184864
rect 429198 183152 429254 183161
rect 429198 183087 429254 183096
rect 427082 179480 427138 179489
rect 427082 179415 427138 179424
rect 428462 179480 428518 179489
rect 428462 179415 428518 179424
rect 426360 176718 426480 176746
rect 425702 176080 425758 176089
rect 425702 176015 425758 176024
rect 421562 175944 421618 175953
rect 421562 175879 421618 175888
rect 295340 172508 295392 172514
rect 295340 172450 295392 172456
rect 421576 166433 421604 175879
rect 421562 166424 421618 166433
rect 421562 166359 421618 166368
rect 425716 165617 425744 176015
rect 426360 175953 426388 176718
rect 427096 176089 427124 179415
rect 427082 176080 427138 176089
rect 427082 176015 427138 176024
rect 426346 175944 426402 175953
rect 426346 175879 426402 175888
rect 425702 165608 425758 165617
rect 425702 165543 425758 165552
rect 292670 141944 292726 141953
rect 292670 141879 292726 141888
rect 458836 140418 458864 386854
rect 462962 368384 463018 368393
rect 462962 368319 463018 368328
rect 462976 359009 463004 368319
rect 462962 359000 463018 359009
rect 462962 358935 463018 358944
rect 459558 358728 459614 358737
rect 459558 358663 459614 358672
rect 459572 356017 459600 358663
rect 462318 357368 462374 357377
rect 462318 357303 462374 357312
rect 459558 356008 459614 356017
rect 459558 355943 459614 355952
rect 462332 350441 462360 357303
rect 458914 350432 458970 350441
rect 458914 350367 458970 350376
rect 462318 350432 462374 350441
rect 462318 350367 462374 350376
rect 458928 347721 458956 350367
rect 463712 348537 463740 390116
rect 467102 378040 467158 378049
rect 467102 377975 467158 377984
rect 467116 371521 467144 377975
rect 465078 371512 465134 371521
rect 465078 371447 465134 371456
rect 467102 371512 467158 371521
rect 467102 371447 467158 371456
rect 464342 371240 464398 371249
rect 464342 371175 464398 371184
rect 464356 357377 464384 371175
rect 465092 368506 465120 371447
rect 465000 368478 465120 368506
rect 465000 368393 465028 368478
rect 464986 368384 465042 368393
rect 464986 368319 465042 368328
rect 464342 357368 464398 357377
rect 464342 357303 464398 357312
rect 463698 348528 463754 348537
rect 463698 348463 463754 348472
rect 458914 347712 458970 347721
rect 458914 347647 458970 347656
rect 458824 140412 458876 140418
rect 458824 140354 458876 140360
rect 467300 139330 467328 390116
rect 469218 382800 469274 382809
rect 469218 382735 469274 382744
rect 469232 378049 469260 382735
rect 469218 378040 469274 378049
rect 469218 377975 469274 377984
rect 467838 375456 467894 375465
rect 467838 375391 467894 375400
rect 467852 371385 467880 375391
rect 467838 371376 467894 371385
rect 467838 371311 467894 371320
rect 470888 139398 470916 390116
rect 473174 388784 473230 388793
rect 473358 388784 473414 388793
rect 473174 388719 473230 388728
rect 473280 388742 473358 388770
rect 473188 388249 473216 388719
rect 473280 388521 473308 388742
rect 473358 388719 473414 388728
rect 473266 388512 473322 388521
rect 473542 388512 473598 388521
rect 473266 388447 473322 388456
rect 473372 388470 473542 388498
rect 473174 388240 473230 388249
rect 473174 388175 473230 388184
rect 471980 386368 472032 386374
rect 471980 386310 472032 386316
rect 471242 384704 471298 384713
rect 471242 384639 471298 384648
rect 471256 375465 471284 384639
rect 471992 382974 472020 386310
rect 473372 385098 473400 388470
rect 473542 388447 473598 388456
rect 473280 385070 473400 385098
rect 473280 384713 473308 385070
rect 473266 384704 473322 384713
rect 473266 384639 473322 384648
rect 471980 382968 472032 382974
rect 471980 382910 472032 382916
rect 471242 375456 471298 375465
rect 471242 375391 471298 375400
rect 474476 355337 474504 390116
rect 479536 389201 479564 449919
rect 479628 411913 479656 529926
rect 479708 520260 479760 520266
rect 479708 520202 479760 520208
rect 479614 411904 479670 411913
rect 479614 411839 479670 411848
rect 479614 403064 479670 403073
rect 479614 402999 479670 403008
rect 476118 389192 476174 389201
rect 474648 389156 474700 389162
rect 476118 389127 476174 389136
rect 479522 389192 479578 389201
rect 479522 389127 479578 389136
rect 474648 389098 474700 389104
rect 474660 387841 474688 389098
rect 476132 388521 476160 389127
rect 476118 388512 476174 388521
rect 476118 388447 476174 388456
rect 474646 387832 474702 387841
rect 474646 387767 474702 387776
rect 479628 386374 479656 402999
rect 479616 386368 479668 386374
rect 479616 386310 479668 386316
rect 479720 386073 479748 520202
rect 479904 501673 479932 538999
rect 479890 501664 479946 501673
rect 479890 501599 479946 501608
rect 479996 479913 480024 637599
rect 480180 528554 480208 657086
rect 480352 644768 480404 644774
rect 480352 644710 480404 644716
rect 480260 637832 480312 637838
rect 480260 637774 480312 637780
rect 480088 528526 480208 528554
rect 480088 518362 480116 528526
rect 480168 520056 480220 520062
rect 480168 519998 480220 520004
rect 480076 518356 480128 518362
rect 480076 518298 480128 518304
rect 480076 518016 480128 518022
rect 480076 517958 480128 517964
rect 480088 517585 480116 517958
rect 480074 517576 480130 517585
rect 480074 517511 480130 517520
rect 480180 516905 480208 519998
rect 480166 516896 480222 516905
rect 480166 516831 480222 516840
rect 479982 479904 480038 479913
rect 479982 479839 480038 479848
rect 480272 465769 480300 637774
rect 480364 474473 480392 644710
rect 480444 640620 480496 640626
rect 480444 640562 480496 640568
rect 480350 474464 480406 474473
rect 480350 474399 480406 474408
rect 480456 474065 480484 640562
rect 484044 600273 484072 657319
rect 484122 657248 484178 657257
rect 484122 657183 484178 657192
rect 484030 600264 484086 600273
rect 484030 600199 484086 600208
rect 484136 600001 484164 657183
rect 484214 657112 484270 657121
rect 484214 657047 484270 657056
rect 484122 599992 484178 600001
rect 484122 599927 484178 599936
rect 484228 563009 484256 657047
rect 484306 655616 484362 655625
rect 484306 655551 484362 655560
rect 484214 563000 484270 563009
rect 484214 562935 484270 562944
rect 482282 554568 482338 554577
rect 482282 554503 482338 554512
rect 481730 550488 481786 550497
rect 481730 550423 481786 550432
rect 480536 544400 480588 544406
rect 480536 544342 480588 544348
rect 480442 474056 480498 474065
rect 480442 473991 480498 474000
rect 480258 465760 480314 465769
rect 480258 465695 480314 465704
rect 480548 405657 480576 544342
rect 480628 541816 480680 541822
rect 480628 541758 480680 541764
rect 480534 405648 480590 405657
rect 480534 405583 480590 405592
rect 479798 405240 479854 405249
rect 479798 405175 479854 405184
rect 479812 388249 479840 405175
rect 480640 404297 480668 541758
rect 480720 538892 480772 538898
rect 480720 538834 480772 538840
rect 480626 404288 480682 404297
rect 480626 404223 480682 404232
rect 480732 402937 480760 538834
rect 480996 537600 481048 537606
rect 480996 537542 481048 537548
rect 480812 537532 480864 537538
rect 480812 537474 480864 537480
rect 480824 403753 480852 537474
rect 480904 534200 480956 534206
rect 480904 534142 480956 534148
rect 480810 403744 480866 403753
rect 480810 403679 480866 403688
rect 480718 402928 480774 402937
rect 480718 402863 480774 402872
rect 480916 402665 480944 534142
rect 481008 408241 481036 537542
rect 481086 532128 481142 532137
rect 481086 532063 481142 532072
rect 481100 413001 481128 532063
rect 481640 523796 481692 523802
rect 481640 523738 481692 523744
rect 481652 523161 481680 523738
rect 481638 523152 481694 523161
rect 481638 523087 481694 523096
rect 481640 518628 481692 518634
rect 481640 518570 481692 518576
rect 481652 511873 481680 518570
rect 481744 513369 481772 550423
rect 481822 542328 481878 542337
rect 481822 542263 481878 542272
rect 481836 514729 481864 542263
rect 482006 536480 482062 536489
rect 482006 536415 482062 536424
rect 481914 533896 481970 533905
rect 481914 533831 481970 533840
rect 481822 514720 481878 514729
rect 481822 514655 481878 514664
rect 481730 513360 481786 513369
rect 481730 513295 481786 513304
rect 481638 511864 481694 511873
rect 481638 511799 481694 511808
rect 481928 511601 481956 533831
rect 482020 515273 482048 536415
rect 482098 530496 482154 530505
rect 482098 530431 482154 530440
rect 482112 518634 482140 530431
rect 482190 523696 482246 523705
rect 482190 523631 482246 523640
rect 482100 518628 482152 518634
rect 482100 518570 482152 518576
rect 482100 518356 482152 518362
rect 482100 518298 482152 518304
rect 482006 515264 482062 515273
rect 482006 515199 482062 515208
rect 481914 511592 481970 511601
rect 481914 511527 481970 511536
rect 481640 510604 481692 510610
rect 481640 510546 481692 510552
rect 481652 507113 481680 510546
rect 482112 510542 482140 518298
rect 482204 515817 482232 523631
rect 482190 515808 482246 515817
rect 482190 515743 482246 515752
rect 482190 514856 482246 514865
rect 482190 514791 482246 514800
rect 482100 510536 482152 510542
rect 482100 510478 482152 510484
rect 481638 507104 481694 507113
rect 481638 507039 481694 507048
rect 482100 480208 482152 480214
rect 482100 480150 482152 480156
rect 482112 479369 482140 480150
rect 482098 479360 482154 479369
rect 482098 479295 482154 479304
rect 482100 478848 482152 478854
rect 482100 478790 482152 478796
rect 482112 478281 482140 478790
rect 482098 478272 482154 478281
rect 482098 478207 482154 478216
rect 482098 474736 482154 474745
rect 482098 474671 482100 474680
rect 482152 474671 482154 474680
rect 482100 474642 482152 474648
rect 482100 473340 482152 473346
rect 482100 473282 482152 473288
rect 482112 472297 482140 473282
rect 482098 472288 482154 472297
rect 482098 472223 482154 472232
rect 482100 471980 482152 471986
rect 482100 471922 482152 471928
rect 482008 471912 482060 471918
rect 482008 471854 482060 471860
rect 482020 471753 482048 471854
rect 482006 471744 482062 471753
rect 482006 471679 482062 471688
rect 482112 471209 482140 471922
rect 482098 471200 482154 471209
rect 482098 471135 482154 471144
rect 482100 470552 482152 470558
rect 482100 470494 482152 470500
rect 482008 470484 482060 470490
rect 482008 470426 482060 470432
rect 482020 470393 482048 470426
rect 482006 470384 482062 470393
rect 482006 470319 482062 470328
rect 482112 469577 482140 470494
rect 482098 469568 482154 469577
rect 482098 469503 482154 469512
rect 482100 469192 482152 469198
rect 482100 469134 482152 469140
rect 482008 469124 482060 469130
rect 482008 469066 482060 469072
rect 482020 468625 482048 469066
rect 482112 469033 482140 469134
rect 482098 469024 482154 469033
rect 482098 468959 482154 468968
rect 482006 468616 482062 468625
rect 482006 468551 482062 468560
rect 482100 467832 482152 467838
rect 482006 467800 482062 467809
rect 482100 467774 482152 467780
rect 482006 467735 482008 467744
rect 482060 467735 482062 467744
rect 482008 467706 482060 467712
rect 482112 466857 482140 467774
rect 482098 466848 482154 466857
rect 482098 466783 482154 466792
rect 482008 465044 482060 465050
rect 482008 464986 482060 464992
rect 482020 464681 482048 464986
rect 482100 464976 482152 464982
rect 482098 464944 482100 464953
rect 482152 464944 482154 464953
rect 482098 464879 482154 464888
rect 482100 464840 482152 464846
rect 482100 464782 482152 464788
rect 482006 464672 482062 464681
rect 482006 464607 482062 464616
rect 482112 464137 482140 464782
rect 482098 464128 482154 464137
rect 482098 464063 482154 464072
rect 482100 463684 482152 463690
rect 482100 463626 482152 463632
rect 482112 463457 482140 463626
rect 482098 463448 482154 463457
rect 482098 463383 482154 463392
rect 482100 463344 482152 463350
rect 482100 463286 482152 463292
rect 482112 463049 482140 463286
rect 482098 463040 482154 463049
rect 482098 462975 482154 462984
rect 482008 462324 482060 462330
rect 482008 462266 482060 462272
rect 481916 462256 481968 462262
rect 481916 462198 481968 462204
rect 481928 461417 481956 462198
rect 482020 461961 482048 462266
rect 482100 462188 482152 462194
rect 482100 462130 482152 462136
rect 482112 462097 482140 462130
rect 482098 462088 482154 462097
rect 482098 462023 482154 462032
rect 482006 461952 482062 461961
rect 482006 461887 482062 461896
rect 481914 461408 481970 461417
rect 481914 461343 481970 461352
rect 482100 460828 482152 460834
rect 482100 460770 482152 460776
rect 482112 460737 482140 460770
rect 482098 460728 482154 460737
rect 482098 460663 482154 460672
rect 482008 459536 482060 459542
rect 482008 459478 482060 459484
rect 482020 458697 482048 459478
rect 482100 459468 482152 459474
rect 482100 459410 482152 459416
rect 482112 459377 482140 459410
rect 482098 459368 482154 459377
rect 482098 459303 482154 459312
rect 482006 458688 482062 458697
rect 482006 458623 482062 458632
rect 482008 458176 482060 458182
rect 482008 458118 482060 458124
rect 482020 457609 482048 458118
rect 482100 458108 482152 458114
rect 482100 458050 482152 458056
rect 482112 458017 482140 458050
rect 482098 458008 482154 458017
rect 482098 457943 482154 457952
rect 482006 457600 482062 457609
rect 482006 457535 482062 457544
rect 482100 456748 482152 456754
rect 482100 456690 482152 456696
rect 482112 456657 482140 456690
rect 482098 456648 482154 456657
rect 482098 456583 482154 456592
rect 482008 455388 482060 455394
rect 482008 455330 482060 455336
rect 482020 454889 482048 455330
rect 482100 455320 482152 455326
rect 482098 455288 482100 455297
rect 482152 455288 482154 455297
rect 482098 455223 482154 455232
rect 482006 454880 482062 454889
rect 482006 454815 482062 454824
rect 482100 454028 482152 454034
rect 482100 453970 482152 453976
rect 482112 453801 482140 453970
rect 482098 453792 482154 453801
rect 482098 453727 482154 453736
rect 482100 452600 482152 452606
rect 482098 452568 482100 452577
rect 482152 452568 482154 452577
rect 482098 452503 482154 452512
rect 482100 452464 482152 452470
rect 482100 452406 482152 452412
rect 482112 451625 482140 452406
rect 482098 451616 482154 451625
rect 482098 451551 482154 451560
rect 482204 449993 482232 514791
rect 482296 510921 482324 554503
rect 483754 554160 483810 554169
rect 483754 554095 483810 554104
rect 483202 550216 483258 550225
rect 483202 550151 483258 550160
rect 482558 523560 482614 523569
rect 482558 523495 482614 523504
rect 482374 522200 482430 522209
rect 482374 522135 482430 522144
rect 482388 514185 482416 522135
rect 482466 520976 482522 520985
rect 482466 520911 482522 520920
rect 482374 514176 482430 514185
rect 482374 514111 482430 514120
rect 482374 512000 482430 512009
rect 482374 511935 482430 511944
rect 482282 510912 482338 510921
rect 482282 510847 482338 510856
rect 482282 510504 482338 510513
rect 482282 510439 482338 510448
rect 482190 449984 482246 449993
rect 482190 449919 482246 449928
rect 482192 449880 482244 449886
rect 482190 449848 482192 449857
rect 482244 449848 482246 449857
rect 482100 449812 482152 449818
rect 482190 449783 482246 449792
rect 482100 449754 482152 449760
rect 482112 449449 482140 449754
rect 482192 449744 482244 449750
rect 482192 449686 482244 449692
rect 482098 449440 482154 449449
rect 482098 449375 482154 449384
rect 482204 448905 482232 449686
rect 482190 448896 482246 448905
rect 482190 448831 482246 448840
rect 482192 448520 482244 448526
rect 482192 448462 482244 448468
rect 482100 448452 482152 448458
rect 482100 448394 482152 448400
rect 482112 447953 482140 448394
rect 482204 448361 482232 448462
rect 482190 448352 482246 448361
rect 482190 448287 482246 448296
rect 482098 447944 482154 447953
rect 482098 447879 482154 447888
rect 482008 447092 482060 447098
rect 482008 447034 482060 447040
rect 482020 446729 482048 447034
rect 482100 447024 482152 447030
rect 482100 446966 482152 446972
rect 482190 446992 482246 447001
rect 482006 446720 482062 446729
rect 482006 446655 482062 446664
rect 482112 446185 482140 446966
rect 482190 446927 482192 446936
rect 482244 446927 482246 446936
rect 482192 446898 482244 446904
rect 482098 446176 482154 446185
rect 482098 446111 482154 446120
rect 482100 445732 482152 445738
rect 482100 445674 482152 445680
rect 482112 445233 482140 445674
rect 482192 445664 482244 445670
rect 482192 445606 482244 445612
rect 482204 445505 482232 445606
rect 482190 445496 482246 445505
rect 482190 445431 482246 445440
rect 482098 445224 482154 445233
rect 482098 445159 482154 445168
rect 482192 444372 482244 444378
rect 482192 444314 482244 444320
rect 482100 444304 482152 444310
rect 482204 444281 482232 444314
rect 482100 444246 482152 444252
rect 482190 444272 482246 444281
rect 482112 444009 482140 444246
rect 482190 444207 482246 444216
rect 482098 444000 482154 444009
rect 482098 443935 482154 443944
rect 482192 442944 482244 442950
rect 482192 442886 482244 442892
rect 482204 442785 482232 442886
rect 482190 442776 482246 442785
rect 482190 442711 482246 442720
rect 482100 441584 482152 441590
rect 482100 441526 482152 441532
rect 482112 441289 482140 441526
rect 482192 441516 482244 441522
rect 482192 441458 482244 441464
rect 482098 441280 482154 441289
rect 482098 441215 482154 441224
rect 482204 440745 482232 441458
rect 482190 440736 482246 440745
rect 482190 440671 482246 440680
rect 482192 440224 482244 440230
rect 482192 440166 482244 440172
rect 482204 440065 482232 440166
rect 482190 440056 482246 440065
rect 482190 439991 482246 440000
rect 482100 438864 482152 438870
rect 482100 438806 482152 438812
rect 482190 438832 482246 438841
rect 482112 438569 482140 438806
rect 482190 438767 482192 438776
rect 482244 438767 482246 438776
rect 482192 438738 482244 438744
rect 482098 438560 482154 438569
rect 482098 438495 482154 438504
rect 482192 428256 482244 428262
rect 482192 428198 482244 428204
rect 482204 424561 482232 428198
rect 482190 424552 482246 424561
rect 482190 424487 482246 424496
rect 482192 418056 482244 418062
rect 482192 417998 482244 418004
rect 482204 417353 482232 417998
rect 482190 417344 482246 417353
rect 482190 417279 482246 417288
rect 482192 415336 482244 415342
rect 482192 415278 482244 415284
rect 482204 414633 482232 415278
rect 482190 414624 482246 414633
rect 482190 414559 482246 414568
rect 482192 413976 482244 413982
rect 482192 413918 482244 413924
rect 482204 413681 482232 413918
rect 482190 413672 482246 413681
rect 482190 413607 482246 413616
rect 481086 412992 481142 413001
rect 481086 412927 481142 412936
rect 482192 411188 482244 411194
rect 482192 411130 482244 411136
rect 482204 411097 482232 411130
rect 482190 411088 482246 411097
rect 482190 411023 482246 411032
rect 482192 410984 482244 410990
rect 482192 410926 482244 410932
rect 482204 410825 482232 410926
rect 482190 410816 482246 410825
rect 482190 410751 482246 410760
rect 482192 408400 482244 408406
rect 482190 408368 482192 408377
rect 482244 408368 482246 408377
rect 482190 408303 482246 408312
rect 480994 408232 481050 408241
rect 480994 408167 481050 408176
rect 482192 407040 482244 407046
rect 482192 406982 482244 406988
rect 482204 406609 482232 406982
rect 482190 406600 482246 406609
rect 482190 406535 482246 406544
rect 480902 402656 480958 402665
rect 480902 402591 480958 402600
rect 482192 400172 482244 400178
rect 482192 400114 482244 400120
rect 482204 399401 482232 400114
rect 482190 399392 482246 399401
rect 482190 399327 482246 399336
rect 482008 398812 482060 398818
rect 482008 398754 482060 398760
rect 482020 398449 482048 398754
rect 482192 398676 482244 398682
rect 482192 398618 482244 398624
rect 482006 398440 482062 398449
rect 482006 398375 482062 398384
rect 482204 397769 482232 398618
rect 482190 397760 482246 397769
rect 482190 397695 482246 397704
rect 482192 397384 482244 397390
rect 482192 397326 482244 397332
rect 482204 396681 482232 397326
rect 482190 396672 482246 396681
rect 482190 396607 482246 396616
rect 482192 396024 482244 396030
rect 482192 395966 482244 395972
rect 482204 395729 482232 395966
rect 482190 395720 482246 395729
rect 482190 395655 482246 395664
rect 482192 394664 482244 394670
rect 482192 394606 482244 394612
rect 482204 393961 482232 394606
rect 482190 393952 482246 393961
rect 482190 393887 482246 393896
rect 482192 393304 482244 393310
rect 482192 393246 482244 393252
rect 482100 393236 482152 393242
rect 482100 393178 482152 393184
rect 482112 392329 482140 393178
rect 482098 392320 482154 392329
rect 482098 392255 482154 392264
rect 482204 388385 482232 393246
rect 482190 388376 482246 388385
rect 482190 388311 482246 388320
rect 479798 388240 479854 388249
rect 479798 388175 479854 388184
rect 482296 387705 482324 510439
rect 482282 387696 482338 387705
rect 482282 387631 482338 387640
rect 477498 386064 477554 386073
rect 477498 385999 477554 386008
rect 479706 386064 479762 386073
rect 479706 385999 479762 386008
rect 477512 382809 477540 385999
rect 477498 382800 477554 382809
rect 477498 382735 477554 382744
rect 474462 355328 474518 355337
rect 474462 355263 474518 355272
rect 482388 164801 482416 511935
rect 482480 510377 482508 520911
rect 482572 513097 482600 523495
rect 482926 520840 482982 520849
rect 482926 520775 482982 520784
rect 482940 514865 482968 520775
rect 483020 519512 483072 519518
rect 483020 519454 483072 519460
rect 483032 519081 483060 519454
rect 483018 519072 483074 519081
rect 483018 519007 483074 519016
rect 483112 518084 483164 518090
rect 483112 518026 483164 518032
rect 483018 517576 483074 517585
rect 483018 517511 483074 517520
rect 482926 514856 482982 514865
rect 482926 514791 482982 514800
rect 482558 513088 482614 513097
rect 482558 513023 482614 513032
rect 482560 510536 482612 510542
rect 483032 510513 483060 517511
rect 483124 510610 483152 518026
rect 483112 510604 483164 510610
rect 483112 510546 483164 510552
rect 482560 510478 482612 510484
rect 483018 510504 483074 510513
rect 482466 510368 482522 510377
rect 482466 510303 482522 510312
rect 482466 495544 482522 495553
rect 482466 495479 482522 495488
rect 482480 342961 482508 495479
rect 482572 393122 482600 510478
rect 483018 510439 483074 510448
rect 482650 508600 482706 508609
rect 482650 508535 482706 508544
rect 482664 393310 482692 508535
rect 482836 506456 482888 506462
rect 482836 506398 482888 506404
rect 482848 506161 482876 506398
rect 482928 506388 482980 506394
rect 482928 506330 482980 506336
rect 482940 506297 482968 506330
rect 482926 506288 482982 506297
rect 482926 506223 482982 506232
rect 482834 506152 482890 506161
rect 482834 506087 482890 506096
rect 482836 500948 482888 500954
rect 482836 500890 482888 500896
rect 482848 500041 482876 500890
rect 482928 500880 482980 500886
rect 482928 500822 482980 500828
rect 482940 500585 482968 500822
rect 482926 500576 482982 500585
rect 482926 500511 482982 500520
rect 482834 500032 482890 500041
rect 482834 499967 482890 499976
rect 482834 494728 482890 494737
rect 482834 494663 482890 494672
rect 482742 492008 482798 492017
rect 482742 491943 482798 491952
rect 482652 393304 482704 393310
rect 482652 393246 482704 393252
rect 482572 393094 482692 393122
rect 482664 387598 482692 393094
rect 482652 387592 482704 387598
rect 482652 387534 482704 387540
rect 482756 383353 482784 491943
rect 482848 428262 482876 494663
rect 482926 491872 482982 491881
rect 482926 491807 482982 491816
rect 482836 428256 482888 428262
rect 482836 428198 482888 428204
rect 482836 425060 482888 425066
rect 482836 425002 482888 425008
rect 482848 424833 482876 425002
rect 482834 424824 482890 424833
rect 482834 424759 482890 424768
rect 482836 423632 482888 423638
rect 482836 423574 482888 423580
rect 482848 423473 482876 423574
rect 482834 423464 482890 423473
rect 482834 423399 482890 423408
rect 482836 423360 482888 423366
rect 482834 423328 482836 423337
rect 482888 423328 482890 423337
rect 482834 423263 482890 423272
rect 482836 418124 482888 418130
rect 482836 418066 482888 418072
rect 482848 418033 482876 418066
rect 482834 418024 482890 418033
rect 482834 417959 482890 417968
rect 482836 416764 482888 416770
rect 482836 416706 482888 416712
rect 482848 416673 482876 416706
rect 482834 416664 482890 416673
rect 482834 416599 482890 416608
rect 482836 415404 482888 415410
rect 482836 415346 482888 415352
rect 482848 415177 482876 415346
rect 482834 415168 482890 415177
rect 482834 415103 482890 415112
rect 482836 413908 482888 413914
rect 482836 413850 482888 413856
rect 482848 413817 482876 413850
rect 482834 413808 482890 413817
rect 482834 413743 482890 413752
rect 482836 412548 482888 412554
rect 482836 412490 482888 412496
rect 482848 412457 482876 412490
rect 482834 412448 482890 412457
rect 482834 412383 482890 412392
rect 482836 411256 482888 411262
rect 482836 411198 482888 411204
rect 482848 410417 482876 411198
rect 482834 410408 482890 410417
rect 482834 410343 482890 410352
rect 482836 409828 482888 409834
rect 482836 409770 482888 409776
rect 482848 409601 482876 409770
rect 482834 409592 482890 409601
rect 482834 409527 482890 409536
rect 482836 408468 482888 408474
rect 482836 408410 482888 408416
rect 482848 407561 482876 408410
rect 482834 407552 482890 407561
rect 482834 407487 482890 407496
rect 482836 407108 482888 407114
rect 482836 407050 482888 407056
rect 482848 406881 482876 407050
rect 482834 406872 482890 406881
rect 482834 406807 482890 406816
rect 482836 405680 482888 405686
rect 482836 405622 482888 405628
rect 482848 404841 482876 405622
rect 482834 404832 482890 404841
rect 482834 404767 482890 404776
rect 482836 402960 482888 402966
rect 482836 402902 482888 402908
rect 482848 402121 482876 402902
rect 482834 402112 482890 402121
rect 482834 402047 482890 402056
rect 482836 401600 482888 401606
rect 482836 401542 482888 401548
rect 482848 401441 482876 401542
rect 482834 401432 482890 401441
rect 482834 401367 482890 401376
rect 482836 401328 482888 401334
rect 482836 401270 482888 401276
rect 482848 401033 482876 401270
rect 482834 401024 482890 401033
rect 482834 400959 482890 400968
rect 482836 400104 482888 400110
rect 482836 400046 482888 400052
rect 482848 399945 482876 400046
rect 482834 399936 482890 399945
rect 482834 399871 482890 399880
rect 482836 398744 482888 398750
rect 482834 398712 482836 398721
rect 482888 398712 482890 398721
rect 482834 398647 482890 398656
rect 482836 397452 482888 397458
rect 482836 397394 482888 397400
rect 482848 397225 482876 397394
rect 482834 397216 482890 397225
rect 482834 397151 482890 397160
rect 482836 395956 482888 395962
rect 482836 395898 482888 395904
rect 482848 395865 482876 395898
rect 482834 395856 482890 395865
rect 482834 395791 482890 395800
rect 482836 394596 482888 394602
rect 482836 394538 482888 394544
rect 482848 394369 482876 394538
rect 482834 394360 482890 394369
rect 482834 394295 482890 394304
rect 482836 393304 482888 393310
rect 482834 393272 482836 393281
rect 482888 393272 482890 393281
rect 482940 393258 482968 491807
rect 483216 426737 483244 550151
rect 483294 541920 483350 541929
rect 483294 541855 483350 541864
rect 483202 426728 483258 426737
rect 483202 426663 483258 426672
rect 483308 426193 483336 541855
rect 483478 538928 483534 538937
rect 483478 538863 483534 538872
rect 483386 537840 483442 537849
rect 483386 537775 483442 537784
rect 483400 428369 483428 537775
rect 483492 430817 483520 538863
rect 483570 535392 483626 535401
rect 483570 535327 483626 535336
rect 483584 432177 483612 535327
rect 483662 530360 483718 530369
rect 483662 530295 483718 530304
rect 483676 436257 483704 530295
rect 483768 437073 483796 554095
rect 483846 545864 483902 545873
rect 483846 545799 483902 545808
rect 483754 437064 483810 437073
rect 483754 436999 483810 437008
rect 483662 436248 483718 436257
rect 483662 436183 483718 436192
rect 483570 432168 483626 432177
rect 483570 432103 483626 432112
rect 483478 430808 483534 430817
rect 483478 430743 483534 430752
rect 483386 428360 483442 428369
rect 483386 428295 483442 428304
rect 483294 426184 483350 426193
rect 483294 426119 483350 426128
rect 483860 421569 483888 545799
rect 484320 532137 484348 655551
rect 485608 599690 485636 657698
rect 485688 657212 485740 657218
rect 485688 657154 485740 657160
rect 485596 599684 485648 599690
rect 485596 599626 485648 599632
rect 485700 599622 485728 657154
rect 486700 643544 486752 643550
rect 486700 643486 486752 643492
rect 485962 640792 486018 640801
rect 485962 640727 486018 640736
rect 485872 640688 485924 640694
rect 485872 640630 485924 640636
rect 485780 639600 485832 639606
rect 485780 639542 485832 639548
rect 485792 639033 485820 639542
rect 485778 639024 485834 639033
rect 485778 638959 485834 638968
rect 485688 599616 485740 599622
rect 485688 599558 485740 599564
rect 485134 558512 485190 558521
rect 485134 558447 485190 558456
rect 484398 551576 484454 551585
rect 484398 551511 484454 551520
rect 484306 532128 484362 532137
rect 484306 532063 484362 532072
rect 484412 431089 484440 551511
rect 484490 548720 484546 548729
rect 484490 548655 484546 548664
rect 484398 431080 484454 431089
rect 484398 431015 484454 431024
rect 484504 429457 484532 548655
rect 484582 543280 484638 543289
rect 484582 543215 484638 543224
rect 484490 429448 484546 429457
rect 484490 429383 484546 429392
rect 484596 428913 484624 543215
rect 484674 540696 484730 540705
rect 484674 540631 484730 540640
rect 484688 430001 484716 540631
rect 484766 537976 484822 537985
rect 484766 537911 484822 537920
rect 484780 436529 484808 537911
rect 484950 532264 485006 532273
rect 484950 532199 485006 532208
rect 484858 526824 484914 526833
rect 484858 526759 484914 526768
rect 484766 436520 484822 436529
rect 484766 436455 484822 436464
rect 484674 429992 484730 430001
rect 484674 429927 484730 429936
rect 484582 428904 484638 428913
rect 484582 428839 484638 428848
rect 484872 428097 484900 526759
rect 484964 434897 484992 532199
rect 485042 525328 485098 525337
rect 485042 525263 485098 525272
rect 484950 434888 485006 434897
rect 484950 434823 485006 434832
rect 485056 432721 485084 525263
rect 485148 494737 485176 558447
rect 485780 546372 485832 546378
rect 485780 546314 485832 546320
rect 485792 545193 485820 546314
rect 485778 545184 485834 545193
rect 485778 545119 485834 545128
rect 485226 523968 485282 523977
rect 485226 523903 485282 523912
rect 485240 503441 485268 523903
rect 485226 503432 485282 503441
rect 485226 503367 485282 503376
rect 485134 494728 485190 494737
rect 485134 494663 485190 494672
rect 485884 474706 485912 640630
rect 485976 480049 486004 640727
rect 486148 547256 486200 547262
rect 486148 547198 486200 547204
rect 486056 538960 486108 538966
rect 486056 538902 486108 538908
rect 485962 480040 486018 480049
rect 485962 479975 486018 479984
rect 485872 474700 485924 474706
rect 485872 474642 485924 474648
rect 485042 432712 485098 432721
rect 485042 432647 485098 432656
rect 484858 428088 484914 428097
rect 484858 428023 484914 428032
rect 483846 421560 483902 421569
rect 483846 421495 483902 421504
rect 486068 411194 486096 538902
rect 486160 423366 486188 547198
rect 486330 544640 486386 544649
rect 486330 544575 486386 544584
rect 486238 541784 486294 541793
rect 486238 541719 486294 541728
rect 486148 423360 486200 423366
rect 486148 423302 486200 423308
rect 486252 422113 486280 541719
rect 486344 435441 486372 544575
rect 486422 533760 486478 533769
rect 486422 533695 486478 533704
rect 486330 435432 486386 435441
rect 486330 435367 486386 435376
rect 486436 433537 486464 533695
rect 486514 529680 486570 529689
rect 486514 529615 486570 529624
rect 486422 433528 486478 433537
rect 486422 433463 486478 433472
rect 486528 431633 486556 529615
rect 486606 526960 486662 526969
rect 486606 526895 486662 526904
rect 486620 433809 486648 526895
rect 486712 470490 486740 643486
rect 486988 599865 487016 657727
rect 501786 657727 501842 657736
rect 494796 657698 494848 657704
rect 487068 656940 487120 656946
rect 487068 656882 487120 656888
rect 499028 656940 499080 656946
rect 499028 656882 499080 656888
rect 486974 599856 487030 599865
rect 486974 599791 487030 599800
rect 487080 599758 487108 656882
rect 497646 656024 497702 656033
rect 497646 655959 497702 655968
rect 494886 655888 494942 655897
rect 494886 655823 494942 655832
rect 492126 655616 492182 655625
rect 492126 655551 492182 655560
rect 492140 654908 492168 655551
rect 494900 654908 494928 655823
rect 496266 655752 496322 655761
rect 496266 655687 496322 655696
rect 496280 654908 496308 655687
rect 497660 654908 497688 655959
rect 499040 654908 499068 656882
rect 501800 654908 501828 657727
rect 503166 657248 503222 657257
rect 507136 657218 507164 670686
rect 508516 657393 508544 700295
rect 527180 700266 527232 700272
rect 510068 657756 510120 657762
rect 510068 657698 510120 657704
rect 508502 657384 508558 657393
rect 508502 657319 508558 657328
rect 503166 657183 503222 657192
rect 507124 657212 507176 657218
rect 503180 654908 503208 657183
rect 507124 657154 507176 657160
rect 504546 657112 504602 657121
rect 504546 657047 504602 657056
rect 504560 654908 504588 657047
rect 505928 655716 505980 655722
rect 505928 655658 505980 655664
rect 505940 654908 505968 655658
rect 507136 654922 507164 657154
rect 508516 654922 508544 657319
rect 507136 654894 507334 654922
rect 508516 654894 508714 654922
rect 510080 654908 510108 657698
rect 512828 657688 512880 657694
rect 512828 657630 512880 657636
rect 514206 657656 514262 657665
rect 511448 657144 511500 657150
rect 511448 657086 511500 657092
rect 511460 654908 511488 657086
rect 512840 654908 512868 657630
rect 534906 657656 534962 657665
rect 514206 657591 514262 657600
rect 521108 657620 521160 657626
rect 514220 654908 514248 657591
rect 534906 657591 534962 657600
rect 521108 657562 521160 657568
rect 519728 657552 519780 657558
rect 515586 657520 515642 657529
rect 519728 657494 519780 657500
rect 515586 657455 515642 657464
rect 515600 654908 515628 657455
rect 518348 657280 518400 657286
rect 518348 657222 518400 657228
rect 516968 657076 517020 657082
rect 516968 657018 517020 657024
rect 516980 654908 517008 657018
rect 518360 654908 518388 657222
rect 519740 654908 519768 657494
rect 521120 654908 521148 657562
rect 532146 657520 532202 657529
rect 532146 657455 532202 657464
rect 529386 657384 529442 657393
rect 529386 657319 529442 657328
rect 528008 657076 528060 657082
rect 528008 657018 528060 657024
rect 526628 657008 526680 657014
rect 526628 656950 526680 656956
rect 525248 655648 525300 655654
rect 525248 655590 525300 655596
rect 522488 655580 522540 655586
rect 522488 655522 522540 655528
rect 522500 654908 522528 655522
rect 525260 654908 525288 655590
rect 526640 654908 526668 656950
rect 528020 654908 528048 657018
rect 529400 654908 529428 657319
rect 530766 657248 530822 657257
rect 530766 657183 530822 657192
rect 530780 654908 530808 657183
rect 532160 654908 532188 657455
rect 533528 657008 533580 657014
rect 533528 656950 533580 656956
rect 533540 654908 533568 656950
rect 534920 654908 534948 657591
rect 536286 657112 536342 657121
rect 536286 657047 536342 657056
rect 536300 654908 536328 657047
rect 537666 656976 537722 656985
rect 537666 656911 537722 656920
rect 539048 656940 539100 656946
rect 537680 654908 537708 656911
rect 539048 656882 539100 656888
rect 539060 654908 539088 656882
rect 540336 655716 540388 655722
rect 540336 655658 540388 655664
rect 493506 654664 493562 654673
rect 493506 654599 493562 654608
rect 488446 654528 488502 654537
rect 488446 654463 488502 654472
rect 500406 654528 500462 654537
rect 523512 654498 523894 654514
rect 500406 654463 500462 654472
rect 523500 654492 523894 654498
rect 488080 644564 488132 644570
rect 488080 644506 488132 644512
rect 487526 640656 487582 640665
rect 487526 640591 487582 640600
rect 487252 639056 487304 639062
rect 487252 638998 487304 639004
rect 487160 638240 487212 638246
rect 487160 638182 487212 638188
rect 487172 637673 487200 638182
rect 487158 637664 487214 637673
rect 487158 637599 487214 637608
rect 487158 613728 487214 613737
rect 487158 613663 487214 613672
rect 487172 612814 487200 613663
rect 487160 612808 487212 612814
rect 487160 612750 487212 612756
rect 487068 599752 487120 599758
rect 487068 599694 487120 599700
rect 487160 559564 487212 559570
rect 487160 559506 487212 559512
rect 487172 559065 487200 559506
rect 487158 559056 487214 559065
rect 487158 558991 487214 559000
rect 486700 470484 486752 470490
rect 486700 470426 486752 470432
rect 487264 467838 487292 638998
rect 487436 637764 487488 637770
rect 487436 637706 487488 637712
rect 487344 635112 487396 635118
rect 487344 635054 487396 635060
rect 487252 467832 487304 467838
rect 487252 467774 487304 467780
rect 487356 467770 487384 635054
rect 487448 471918 487476 637706
rect 487540 475153 487568 640591
rect 487710 551304 487766 551313
rect 487710 551239 487766 551248
rect 487620 549296 487672 549302
rect 487620 549238 487672 549244
rect 487526 475144 487582 475153
rect 487526 475079 487582 475088
rect 487436 471912 487488 471918
rect 487436 471854 487488 471860
rect 487344 467764 487396 467770
rect 487344 467706 487396 467712
rect 486606 433800 486662 433809
rect 486606 433735 486662 433744
rect 486514 431624 486570 431633
rect 486514 431559 486570 431568
rect 486238 422104 486294 422113
rect 486238 422039 486294 422048
rect 486056 411188 486108 411194
rect 486056 411130 486108 411136
rect 487632 408406 487660 549238
rect 487724 408785 487752 551239
rect 487804 540456 487856 540462
rect 487804 540398 487856 540404
rect 487816 410990 487844 540398
rect 487896 535628 487948 535634
rect 487896 535570 487948 535576
rect 487804 410984 487856 410990
rect 487804 410926 487856 410932
rect 487908 409834 487936 535570
rect 487988 534336 488040 534342
rect 487988 534278 488040 534284
rect 488000 412554 488028 534278
rect 488092 463350 488120 644506
rect 488460 600137 488488 654463
rect 523552 654486 523894 654492
rect 523500 654434 523552 654440
rect 490737 654200 490746 654256
rect 490802 654200 490811 654256
rect 540242 652896 540298 652905
rect 540242 652831 540298 652840
rect 489368 644632 489420 644638
rect 489368 644574 489420 644580
rect 488540 641912 488592 641918
rect 488540 641854 488592 641860
rect 488998 641880 489054 641889
rect 488552 641753 488580 641854
rect 488998 641815 489054 641824
rect 488538 641744 488594 641753
rect 488538 641679 488594 641688
rect 488816 640552 488868 640558
rect 488816 640494 488868 640500
rect 488722 639976 488778 639985
rect 488722 639911 488778 639920
rect 488632 638988 488684 638994
rect 488632 638930 488684 638936
rect 488540 637900 488592 637906
rect 488540 637842 488592 637848
rect 488552 637673 488580 637842
rect 488538 637664 488594 637673
rect 488538 637599 488594 637608
rect 488446 600128 488502 600137
rect 488446 600063 488502 600072
rect 488080 463344 488132 463350
rect 488080 463286 488132 463292
rect 488644 460834 488672 638930
rect 488736 469713 488764 639911
rect 488828 473346 488856 640494
rect 488906 639160 488962 639169
rect 488906 639095 488962 639104
rect 488816 473340 488868 473346
rect 488816 473282 488868 473288
rect 488920 472977 488948 639095
rect 489012 476785 489040 641815
rect 489092 553512 489144 553518
rect 489092 553454 489144 553460
rect 488998 476776 489054 476785
rect 488998 476711 489054 476720
rect 488906 472968 488962 472977
rect 488906 472903 488962 472912
rect 488722 469704 488778 469713
rect 488722 469639 488778 469648
rect 488632 460828 488684 460834
rect 488632 460770 488684 460776
rect 487988 412548 488040 412554
rect 487988 412490 488040 412496
rect 487896 409828 487948 409834
rect 487896 409770 487948 409776
rect 487710 408776 487766 408785
rect 487710 408711 487766 408720
rect 487620 408400 487672 408406
rect 487620 408342 487672 408348
rect 489104 401334 489132 553454
rect 489276 530596 489328 530602
rect 489276 530538 489328 530544
rect 489182 525192 489238 525201
rect 489182 525127 489238 525136
rect 489196 425649 489224 525127
rect 489288 452470 489316 530538
rect 489380 464846 489408 644574
rect 490104 644496 490156 644502
rect 490104 644438 490156 644444
rect 489920 643204 489972 643210
rect 489920 643146 489972 643152
rect 489368 464840 489420 464846
rect 489368 464782 489420 464788
rect 489932 455326 489960 643146
rect 490012 641844 490064 641850
rect 490012 641786 490064 641792
rect 490024 458114 490052 641786
rect 490116 462194 490144 644438
rect 490196 640416 490248 640422
rect 490196 640358 490248 640364
rect 490208 463690 490236 640358
rect 539782 630592 539838 630601
rect 539782 630527 539838 630536
rect 539598 627872 539654 627881
rect 539598 627807 539654 627816
rect 539506 612776 539562 612785
rect 539506 612711 539562 612720
rect 539414 610736 539470 610745
rect 539414 610671 539470 610680
rect 539322 604480 539378 604489
rect 539322 604415 539378 604424
rect 539336 600642 539364 604415
rect 539428 601905 539456 610671
rect 539414 601896 539470 601905
rect 539414 601831 539470 601840
rect 539520 601769 539548 612711
rect 539506 601760 539562 601769
rect 539506 601695 539562 601704
rect 538588 600636 538640 600642
rect 538588 600578 538640 600584
rect 539324 600636 539376 600642
rect 539324 600578 539376 600584
rect 535736 600296 535788 600302
rect 497370 600264 497426 600273
rect 535736 600238 535788 600244
rect 536010 600264 536066 600273
rect 497370 600199 497426 600208
rect 490378 547224 490434 547233
rect 490378 547159 490434 547168
rect 490286 543144 490342 543153
rect 490286 543079 490342 543088
rect 490196 463684 490248 463690
rect 490196 463626 490248 463632
rect 490104 462188 490156 462194
rect 490104 462130 490156 462136
rect 490012 458108 490064 458114
rect 490012 458050 490064 458056
rect 489920 455320 489972 455326
rect 489920 455262 489972 455268
rect 489276 452464 489328 452470
rect 489276 452406 489328 452412
rect 489182 425640 489238 425649
rect 489182 425575 489238 425584
rect 490300 425241 490328 543079
rect 490392 434489 490420 547159
rect 490470 536344 490526 536353
rect 490470 536279 490526 536288
rect 490484 437753 490512 536279
rect 490564 521756 490616 521762
rect 490564 521698 490616 521704
rect 490576 448458 490604 521698
rect 490656 518492 490708 518498
rect 490656 518434 490708 518440
rect 490668 506394 490696 518434
rect 490656 506388 490708 506394
rect 490656 506330 490708 506336
rect 490564 448452 490616 448458
rect 490564 448394 490616 448400
rect 490470 437744 490526 437753
rect 490470 437679 490526 437688
rect 490378 434480 490434 434489
rect 490378 434415 490434 434424
rect 490286 425232 490342 425241
rect 490286 425167 490342 425176
rect 489092 401328 489144 401334
rect 489092 401270 489144 401276
rect 482940 393230 483060 393258
rect 482834 393207 482890 393216
rect 482928 393168 482980 393174
rect 482928 393110 482980 393116
rect 482940 392873 482968 393110
rect 482926 392864 482982 392873
rect 482926 392799 482982 392808
rect 483032 392714 483060 393230
rect 482940 392686 483060 392714
rect 482940 392034 482968 392686
rect 482940 392006 483060 392034
rect 482836 391944 482888 391950
rect 482836 391886 482888 391892
rect 482848 391241 482876 391886
rect 482928 391876 482980 391882
rect 482928 391818 482980 391824
rect 482940 391649 482968 391818
rect 482926 391640 482982 391649
rect 482926 391575 482982 391584
rect 483032 391490 483060 392006
rect 482940 391462 483060 391490
rect 482834 391232 482890 391241
rect 482834 391167 482890 391176
rect 482940 390674 482968 391462
rect 482848 390646 482968 390674
rect 482848 386345 482876 390646
rect 482928 390516 482980 390522
rect 482928 390458 482980 390464
rect 482940 390425 482968 390458
rect 482926 390416 482982 390425
rect 482926 390351 482982 390360
rect 482834 386336 482890 386345
rect 482834 386271 482890 386280
rect 482742 383344 482798 383353
rect 482742 383279 482798 383288
rect 482466 342952 482522 342961
rect 482466 342887 482522 342896
rect 490760 341630 490788 600100
rect 492140 598233 492168 600100
rect 493520 598233 493548 600100
rect 494900 598233 494928 600100
rect 495714 599584 495770 599593
rect 495714 599519 495770 599528
rect 492126 598224 492182 598233
rect 492126 598159 492182 598168
rect 493506 598224 493562 598233
rect 493506 598159 493562 598168
rect 494886 598224 494942 598233
rect 494886 598159 494942 598168
rect 494610 558784 494666 558793
rect 494610 558719 494666 558728
rect 492772 557660 492824 557666
rect 492772 557602 492824 557608
rect 491300 552220 491352 552226
rect 491300 552162 491352 552168
rect 491312 425066 491340 552162
rect 492126 549944 492182 549953
rect 491668 549908 491720 549914
rect 492126 549879 492182 549888
rect 491668 549850 491720 549856
rect 491484 538348 491536 538354
rect 491484 538290 491536 538296
rect 491392 518560 491444 518566
rect 491392 518502 491444 518508
rect 491404 506462 491432 518502
rect 491392 506456 491444 506462
rect 491392 506398 491444 506404
rect 491300 425060 491352 425066
rect 491300 425002 491352 425008
rect 491496 423638 491524 538290
rect 491574 526552 491630 526561
rect 491574 526487 491630 526496
rect 491484 423632 491536 423638
rect 491484 423574 491536 423580
rect 491588 417625 491616 526487
rect 491680 454034 491708 549850
rect 491942 546408 491998 546417
rect 491942 546343 491998 546352
rect 491760 533384 491812 533390
rect 491760 533326 491812 533332
rect 491668 454028 491720 454034
rect 491668 453970 491720 453976
rect 491772 446962 491800 533326
rect 491852 518220 491904 518226
rect 491852 518162 491904 518168
rect 491864 458182 491892 518162
rect 491956 509561 491984 546343
rect 492034 520160 492090 520169
rect 492034 520095 492090 520104
rect 491942 509552 491998 509561
rect 491942 509487 491998 509496
rect 492048 491609 492076 520095
rect 492034 491600 492090 491609
rect 492034 491535 492090 491544
rect 491852 458176 491904 458182
rect 491852 458118 491904 458124
rect 491760 446956 491812 446962
rect 491760 446898 491812 446904
rect 492140 422521 492168 549879
rect 492680 518424 492732 518430
rect 492680 518366 492732 518372
rect 492692 500886 492720 518366
rect 492680 500880 492732 500886
rect 492680 500822 492732 500828
rect 492784 444378 492812 557602
rect 492864 554804 492916 554810
rect 492864 554746 492916 554752
rect 492772 444372 492824 444378
rect 492772 444314 492824 444320
rect 492876 444310 492904 554746
rect 493048 553444 493100 553450
rect 493048 553386 493100 553392
rect 492956 550724 493008 550730
rect 492956 550666 493008 550672
rect 492864 444304 492916 444310
rect 492864 444246 492916 444252
rect 492968 441522 492996 550666
rect 493060 447030 493088 553386
rect 493140 548548 493192 548554
rect 493140 548490 493192 548496
rect 493048 447024 493100 447030
rect 493048 446966 493100 446972
rect 493152 445670 493180 548490
rect 494244 544468 494296 544474
rect 494244 544410 494296 544416
rect 493232 540320 493284 540326
rect 493232 540262 493284 540268
rect 493244 449750 493272 540262
rect 493508 532772 493560 532778
rect 493508 532714 493560 532720
rect 493324 528624 493376 528630
rect 493324 528566 493376 528572
rect 493232 449744 493284 449750
rect 493232 449686 493284 449692
rect 493336 445738 493364 528566
rect 493416 518288 493468 518294
rect 493416 518230 493468 518236
rect 493428 455394 493456 518230
rect 493416 455388 493468 455394
rect 493416 455330 493468 455336
rect 493324 445732 493376 445738
rect 493324 445674 493376 445680
rect 493140 445664 493192 445670
rect 493140 445606 493192 445612
rect 492956 441516 493008 441522
rect 492956 441458 493008 441464
rect 492126 422512 492182 422521
rect 492126 422447 492182 422456
rect 491574 417616 491630 417625
rect 491574 417551 491630 417560
rect 493520 398682 493548 532714
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494060 518968 494112 518974
rect 494060 518910 494112 518916
rect 494072 500954 494100 518910
rect 494060 500948 494112 500954
rect 494060 500890 494112 500896
rect 494164 405686 494192 531286
rect 494256 418130 494284 544410
rect 494428 543040 494480 543046
rect 494428 542982 494480 542988
rect 494336 541000 494388 541006
rect 494336 540942 494388 540948
rect 494244 418124 494296 418130
rect 494244 418066 494296 418072
rect 494348 418062 494376 540942
rect 494440 448526 494468 542982
rect 494520 521688 494572 521694
rect 494520 521630 494572 521636
rect 494532 449818 494560 521630
rect 494624 490521 494652 558719
rect 495440 547188 495492 547194
rect 495440 547130 495492 547136
rect 494888 519988 494940 519994
rect 494888 519930 494940 519936
rect 494704 519920 494756 519926
rect 494704 519862 494756 519868
rect 494610 490512 494666 490521
rect 494610 490447 494666 490456
rect 494716 469130 494744 519862
rect 494796 518152 494848 518158
rect 494796 518094 494848 518100
rect 494808 480214 494836 518094
rect 494796 480208 494848 480214
rect 494796 480150 494848 480156
rect 494704 469124 494756 469130
rect 494704 469066 494756 469072
rect 494520 449812 494572 449818
rect 494520 449754 494572 449760
rect 494428 448520 494480 448526
rect 494428 448462 494480 448468
rect 494336 418056 494388 418062
rect 494336 417998 494388 418004
rect 494152 405680 494204 405686
rect 494152 405622 494204 405628
rect 493508 398676 493560 398682
rect 493508 398618 493560 398624
rect 494900 345014 494928 519930
rect 495452 400110 495480 547130
rect 495532 541680 495584 541686
rect 495532 541622 495584 541628
rect 495440 400104 495492 400110
rect 495440 400046 495492 400052
rect 495544 397390 495572 541622
rect 495622 526416 495678 526425
rect 495622 526351 495678 526360
rect 495636 418713 495664 526351
rect 495728 492017 495756 599519
rect 496082 535120 496138 535129
rect 496082 535055 496138 535064
rect 495990 521384 496046 521393
rect 495990 521319 496046 521328
rect 495806 520160 495862 520169
rect 495806 520095 495862 520104
rect 495714 492008 495770 492017
rect 495714 491943 495770 491952
rect 495622 418704 495678 418713
rect 495622 418639 495678 418648
rect 495820 415449 495848 520095
rect 495900 519852 495952 519858
rect 495900 519794 495952 519800
rect 495912 459474 495940 519794
rect 496004 478553 496032 521319
rect 496096 499225 496124 535055
rect 496082 499216 496138 499225
rect 496082 499151 496138 499160
rect 495990 478544 496046 478553
rect 495990 478479 496046 478488
rect 495900 459468 495952 459474
rect 495900 459410 495952 459416
rect 495806 415440 495862 415449
rect 495806 415375 495862 415384
rect 495532 397384 495584 397390
rect 495532 397326 495584 397332
rect 496280 354113 496308 600100
rect 497004 542496 497056 542502
rect 497004 542438 497056 542444
rect 496912 541748 496964 541754
rect 496912 541690 496964 541696
rect 496818 522336 496874 522345
rect 496818 522271 496874 522280
rect 496832 508473 496860 522271
rect 496818 508464 496874 508473
rect 496818 508399 496874 508408
rect 496924 400178 496952 541690
rect 497016 407046 497044 542438
rect 497188 530120 497240 530126
rect 497188 530062 497240 530068
rect 497096 530052 497148 530058
rect 497096 529994 497148 530000
rect 497108 413914 497136 529994
rect 497200 415410 497228 530062
rect 497280 527264 497332 527270
rect 497280 527206 497332 527212
rect 497188 415404 497240 415410
rect 497188 415346 497240 415352
rect 497292 415342 497320 527206
rect 497384 491881 497412 600199
rect 534724 600160 534776 600166
rect 507858 600128 507914 600137
rect 497660 598233 497688 600100
rect 498200 599752 498252 599758
rect 498200 599694 498252 599700
rect 497646 598224 497702 598233
rect 497646 598159 497702 598168
rect 497464 550656 497516 550662
rect 497464 550598 497516 550604
rect 497370 491872 497426 491881
rect 497370 491807 497426 491816
rect 497476 452606 497504 550598
rect 497556 522436 497608 522442
rect 497556 522378 497608 522384
rect 497568 478854 497596 522378
rect 497646 521656 497702 521665
rect 497646 521591 497702 521600
rect 497556 478848 497608 478854
rect 497556 478790 497608 478796
rect 497464 452600 497516 452606
rect 497464 452542 497516 452548
rect 497280 415336 497332 415342
rect 497280 415278 497332 415284
rect 497096 413908 497148 413914
rect 497096 413850 497148 413856
rect 497004 407040 497056 407046
rect 497004 406982 497056 406988
rect 496912 400172 496964 400178
rect 496912 400114 496964 400120
rect 497660 364334 497688 521591
rect 498212 387598 498240 599694
rect 498382 531992 498438 532001
rect 498382 531927 498438 531936
rect 498292 527876 498344 527882
rect 498292 527818 498344 527824
rect 498304 398750 498332 527818
rect 498396 405113 498424 531927
rect 498566 527912 498622 527921
rect 498566 527847 498622 527856
rect 498476 525904 498528 525910
rect 498476 525846 498528 525852
rect 498488 413982 498516 525846
rect 498580 419801 498608 527847
rect 498750 522064 498806 522073
rect 498750 521999 498806 522008
rect 498660 519784 498712 519790
rect 498660 519726 498712 519732
rect 498672 471986 498700 519726
rect 498764 477465 498792 521999
rect 498750 477456 498806 477465
rect 498750 477391 498806 477400
rect 498660 471980 498712 471986
rect 498660 471922 498712 471928
rect 498566 419792 498622 419801
rect 498566 419727 498622 419736
rect 498476 413976 498528 413982
rect 498476 413918 498528 413924
rect 498382 405104 498438 405113
rect 498382 405039 498438 405048
rect 498292 398744 498344 398750
rect 498292 398686 498344 398692
rect 498200 387592 498252 387598
rect 498200 387534 498252 387540
rect 498844 387592 498896 387598
rect 498844 387534 498896 387540
rect 498212 387122 498240 387534
rect 498200 387116 498252 387122
rect 498200 387058 498252 387064
rect 497476 364306 497688 364334
rect 497476 363633 497504 364306
rect 497462 363624 497518 363633
rect 497462 363559 497518 363568
rect 496266 354104 496322 354113
rect 496266 354039 496322 354048
rect 494716 344986 494928 345014
rect 494716 344350 494744 344986
rect 494704 344344 494756 344350
rect 494704 344286 494756 344292
rect 490748 341624 490800 341630
rect 490748 341566 490800 341572
rect 492586 278080 492642 278089
rect 492586 278015 492642 278024
rect 482374 164792 482430 164801
rect 482374 164727 482430 164736
rect 470876 139392 470928 139398
rect 470876 139334 470928 139340
rect 467288 139324 467340 139330
rect 467288 139266 467340 139272
rect 345664 87372 345716 87378
rect 345664 87314 345716 87320
rect 311438 86184 311494 86193
rect 311438 86119 311494 86128
rect 295984 82816 296036 82822
rect 295984 82758 296036 82764
rect 291844 6860 291896 6866
rect 291844 6802 291896 6808
rect 291752 4072 291804 4078
rect 291752 4014 291804 4020
rect 293682 3496 293738 3505
rect 295996 3466 296024 82758
rect 304354 51912 304410 51921
rect 304354 51847 304410 51856
rect 297270 42256 297326 42265
rect 297270 42191 297326 42200
rect 293682 3431 293738 3440
rect 295984 3460 296036 3466
rect 293696 480 293724 3431
rect 295984 3402 296036 3408
rect 297284 480 297312 42191
rect 300766 3360 300822 3369
rect 300766 3295 300822 3304
rect 300780 480 300808 3295
rect 304368 480 304396 51847
rect 307942 4992 307998 5001
rect 307942 4927 307998 4936
rect 307956 480 307984 4927
rect 311452 480 311480 86119
rect 329194 85640 329250 85649
rect 329194 85575 329250 85584
rect 315026 80744 315082 80753
rect 315026 80679 315082 80688
rect 315040 480 315068 80679
rect 322110 79384 322166 79393
rect 322110 79319 322166 79328
rect 318522 53136 318578 53145
rect 318522 53071 318578 53080
rect 318536 480 318564 53071
rect 322124 480 322152 79319
rect 325606 54632 325662 54641
rect 325606 54567 325662 54576
rect 325620 480 325648 54567
rect 329208 480 329236 85575
rect 343362 84688 343418 84697
rect 343362 84623 343418 84632
rect 336280 83496 336332 83502
rect 336280 83438 336332 83444
rect 334622 58576 334678 58585
rect 334622 58511 334678 58520
rect 334636 7585 334664 58511
rect 332690 7576 332746 7585
rect 332690 7511 332746 7520
rect 334622 7576 334678 7585
rect 334622 7511 334678 7520
rect 332704 480 332732 7511
rect 336292 480 336320 83438
rect 339868 10328 339920 10334
rect 339868 10270 339920 10276
rect 339880 480 339908 10270
rect 343376 480 343404 84623
rect 345676 4214 345704 87314
rect 492600 86193 492628 278015
rect 493968 275324 494020 275330
rect 493968 275266 494020 275272
rect 493980 167006 494008 275266
rect 494716 206990 494744 344286
rect 497476 298761 497504 363559
rect 498856 353258 498884 387534
rect 499040 359417 499068 600100
rect 499578 599720 499634 599729
rect 499578 599655 499634 599664
rect 499026 359408 499082 359417
rect 499026 359343 499082 359352
rect 498844 353252 498896 353258
rect 498844 353194 498896 353200
rect 497462 298752 497518 298761
rect 497462 298687 497518 298696
rect 496728 291848 496780 291854
rect 496728 291790 496780 291796
rect 496740 245614 496768 291790
rect 496728 245608 496780 245614
rect 496728 245550 496780 245556
rect 494704 206984 494756 206990
rect 494704 206926 494756 206932
rect 493968 167000 494020 167006
rect 493968 166942 494020 166948
rect 499592 163985 499620 599655
rect 499762 536208 499818 536217
rect 499762 536143 499818 536152
rect 499672 525972 499724 525978
rect 499672 525914 499724 525920
rect 499684 407114 499712 525914
rect 499776 419257 499804 536143
rect 499946 530904 500002 530913
rect 499946 530839 500002 530848
rect 499856 528692 499908 528698
rect 499856 528634 499908 528640
rect 499762 419248 499818 419257
rect 499762 419183 499818 419192
rect 499868 416770 499896 528634
rect 499960 420345 499988 530839
rect 500040 519716 500092 519722
rect 500040 519658 500092 519664
rect 500052 469198 500080 519658
rect 500132 519648 500184 519654
rect 500132 519590 500184 519596
rect 500144 470558 500172 519590
rect 500132 470552 500184 470558
rect 500132 470494 500184 470500
rect 500040 469192 500092 469198
rect 500040 469134 500092 469140
rect 500222 457464 500278 457473
rect 500222 457399 500278 457408
rect 499946 420336 500002 420345
rect 499946 420271 500002 420280
rect 499856 416764 499908 416770
rect 499856 416706 499908 416712
rect 499672 407108 499724 407114
rect 499672 407050 499724 407056
rect 500236 390153 500264 457399
rect 500222 390144 500278 390153
rect 500222 390079 500278 390088
rect 500420 380089 500448 600100
rect 501144 535492 501196 535498
rect 501144 535434 501196 535440
rect 500960 534132 501012 534138
rect 500960 534074 501012 534080
rect 500972 398818 501000 534074
rect 501052 529236 501104 529242
rect 501052 529178 501104 529184
rect 500960 398812 501012 398818
rect 500960 398754 501012 398760
rect 501064 395962 501092 529178
rect 501156 402966 501184 535434
rect 501234 525056 501290 525065
rect 501234 524991 501290 525000
rect 501248 427417 501276 524991
rect 501326 522744 501382 522753
rect 501326 522679 501382 522688
rect 501340 476377 501368 522679
rect 501418 521248 501474 521257
rect 501418 521183 501474 521192
rect 501432 480729 501460 521183
rect 501510 519752 501566 519761
rect 501510 519687 501566 519696
rect 501524 482361 501552 519687
rect 501510 482352 501566 482361
rect 501510 482287 501566 482296
rect 501418 480720 501474 480729
rect 501418 480655 501474 480664
rect 501326 476368 501382 476377
rect 501326 476303 501382 476312
rect 501234 427408 501290 427417
rect 501234 427343 501290 427352
rect 501144 402960 501196 402966
rect 501144 402902 501196 402908
rect 501052 395956 501104 395962
rect 501052 395898 501104 395904
rect 500406 380080 500462 380089
rect 500406 380015 500462 380024
rect 501800 364993 501828 600100
rect 502984 598256 503036 598262
rect 502984 598198 503036 598204
rect 502524 552152 502576 552158
rect 502524 552094 502576 552100
rect 502340 548616 502392 548622
rect 502340 548558 502392 548564
rect 502352 408474 502380 548558
rect 502432 532840 502484 532846
rect 502432 532782 502484 532788
rect 502340 408468 502392 408474
rect 502340 408410 502392 408416
rect 502444 401606 502472 532782
rect 502536 438802 502564 552094
rect 502706 522608 502762 522617
rect 502706 522543 502762 522552
rect 502616 522368 502668 522374
rect 502616 522310 502668 522316
rect 502628 462262 502656 522310
rect 502720 472569 502748 522543
rect 502706 472560 502762 472569
rect 502706 472495 502762 472504
rect 502616 462256 502668 462262
rect 502616 462198 502668 462204
rect 502524 438796 502576 438802
rect 502524 438738 502576 438744
rect 502432 401600 502484 401606
rect 502432 401542 502484 401548
rect 501786 364984 501842 364993
rect 501786 364919 501842 364928
rect 502996 340338 503024 598198
rect 503074 512000 503130 512009
rect 503074 511935 503130 511944
rect 503088 389065 503116 511935
rect 503074 389056 503130 389065
rect 503074 388991 503130 389000
rect 503180 374649 503208 600100
rect 504086 599992 504142 600001
rect 504086 599927 504142 599936
rect 503810 563000 503866 563009
rect 503810 562935 503866 562944
rect 503720 522640 503772 522646
rect 503720 522582 503772 522588
rect 503166 374640 503222 374649
rect 503166 374575 503222 374584
rect 502984 340332 503036 340338
rect 502984 340274 503036 340280
rect 503732 340202 503760 522582
rect 503824 388929 503852 562935
rect 503996 545760 504048 545766
rect 503996 545702 504048 545708
rect 503904 540252 503956 540258
rect 503904 540194 503956 540200
rect 503916 397458 503944 540194
rect 504008 411262 504036 545702
rect 504100 512009 504128 599927
rect 504178 564360 504234 564369
rect 504178 564295 504234 564304
rect 504192 563009 504220 564295
rect 504178 563000 504234 563009
rect 504178 562935 504234 562944
rect 504180 522572 504232 522578
rect 504180 522514 504232 522520
rect 504086 512000 504142 512009
rect 504086 511935 504142 511944
rect 504100 511329 504128 511935
rect 504086 511320 504142 511329
rect 504086 511255 504142 511264
rect 504192 459542 504220 522514
rect 504362 521520 504418 521529
rect 504362 521455 504418 521464
rect 504272 521280 504324 521286
rect 504272 521222 504324 521228
rect 504284 464982 504312 521222
rect 504376 481817 504404 521455
rect 504362 481808 504418 481817
rect 504362 481743 504418 481752
rect 504272 464976 504324 464982
rect 504272 464918 504324 464924
rect 504180 459536 504232 459542
rect 504180 459478 504232 459484
rect 503996 411256 504048 411262
rect 503996 411198 504048 411204
rect 503904 397452 503956 397458
rect 503904 397394 503956 397400
rect 503810 388920 503866 388929
rect 503810 388855 503866 388864
rect 504560 345681 504588 600100
rect 505100 599684 505152 599690
rect 505100 599626 505152 599632
rect 505112 387666 505140 599626
rect 505466 555928 505522 555937
rect 505466 555863 505522 555872
rect 505192 525836 505244 525842
rect 505192 525778 505244 525784
rect 505204 440230 505232 525778
rect 505376 521212 505428 521218
rect 505376 521154 505428 521160
rect 505284 521076 505336 521082
rect 505284 521018 505336 521024
rect 505296 462330 505324 521018
rect 505388 465050 505416 521154
rect 505480 503033 505508 555863
rect 505558 521112 505614 521121
rect 505558 521047 505614 521056
rect 505466 503024 505522 503033
rect 505466 502959 505522 502968
rect 505572 481273 505600 521047
rect 505558 481264 505614 481273
rect 505558 481199 505614 481208
rect 505376 465044 505428 465050
rect 505376 464986 505428 464992
rect 505284 462324 505336 462330
rect 505284 462266 505336 462272
rect 505192 440224 505244 440230
rect 505192 440166 505244 440172
rect 505100 387660 505152 387666
rect 505100 387602 505152 387608
rect 505940 383081 505968 600100
rect 506480 599616 506532 599622
rect 506480 599558 506532 599564
rect 506492 387734 506520 599558
rect 506664 558476 506716 558482
rect 506664 558418 506716 558424
rect 506572 522504 506624 522510
rect 506572 522446 506624 522452
rect 506480 387728 506532 387734
rect 506480 387670 506532 387676
rect 505926 383072 505982 383081
rect 505926 383007 505982 383016
rect 506584 355366 506612 522446
rect 506676 393174 506704 558418
rect 506938 540560 506994 540569
rect 506938 540495 506994 540504
rect 506756 536104 506808 536110
rect 506756 536046 506808 536052
rect 506768 438870 506796 536046
rect 506848 524476 506900 524482
rect 506848 524418 506900 524424
rect 506860 442950 506888 524418
rect 506952 494873 506980 540495
rect 506938 494864 506994 494873
rect 506938 494799 506994 494808
rect 506848 442944 506900 442950
rect 506848 442886 506900 442892
rect 506756 438864 506808 438870
rect 506756 438806 506808 438812
rect 506664 393168 506716 393174
rect 506664 393110 506716 393116
rect 506572 355360 506624 355366
rect 506572 355302 506624 355308
rect 506584 354674 506612 355302
rect 506492 354646 506612 354674
rect 504546 345672 504602 345681
rect 504546 345607 504602 345616
rect 503720 340196 503772 340202
rect 503720 340138 503772 340144
rect 503732 291854 503760 340138
rect 503720 291848 503772 291854
rect 503720 291790 503772 291796
rect 506492 275330 506520 354646
rect 507320 341562 507348 600100
rect 534724 600102 534776 600108
rect 507858 600063 507914 600072
rect 507872 405249 507900 600063
rect 508042 599856 508098 599865
rect 508042 599791 508098 599800
rect 507950 532128 508006 532137
rect 507950 532063 508006 532072
rect 507858 405240 507914 405249
rect 507858 405175 507914 405184
rect 507964 347041 507992 532063
rect 508056 457473 508084 599791
rect 508136 536852 508188 536858
rect 508136 536794 508188 536800
rect 508042 457464 508098 457473
rect 508042 457399 508098 457408
rect 508148 447098 508176 536794
rect 508228 524544 508280 524550
rect 508228 524486 508280 524492
rect 508136 447092 508188 447098
rect 508136 447034 508188 447040
rect 508240 441590 508268 524486
rect 508228 441584 508280 441590
rect 508228 441526 508280 441532
rect 508700 382945 508728 600100
rect 509424 557592 509476 557598
rect 509424 557534 509476 557540
rect 509332 552424 509384 552430
rect 509332 552366 509384 552372
rect 509240 519580 509292 519586
rect 509240 519522 509292 519528
rect 509252 393242 509280 519522
rect 509344 449886 509372 552366
rect 509436 456754 509464 557534
rect 509424 456748 509476 456754
rect 509424 456690 509476 456696
rect 509332 449880 509384 449886
rect 509332 449822 509384 449828
rect 509240 393236 509292 393242
rect 509240 393178 509292 393184
rect 508686 382936 508742 382945
rect 508686 382871 508742 382880
rect 510080 380905 510108 600100
rect 510620 522300 510672 522306
rect 510620 522242 510672 522248
rect 510632 390522 510660 522242
rect 510620 390516 510672 390522
rect 510620 390458 510672 390464
rect 510066 380896 510122 380905
rect 510066 380831 510122 380840
rect 511460 362273 511488 600100
rect 511906 599040 511962 599049
rect 511906 598975 511962 598984
rect 511920 485897 511948 598975
rect 512000 558272 512052 558278
rect 512000 558214 512052 558220
rect 511906 485888 511962 485897
rect 511906 485823 511962 485832
rect 512012 391950 512040 558214
rect 512092 556912 512144 556918
rect 512092 556854 512144 556860
rect 512104 394602 512132 556854
rect 512184 521144 512236 521150
rect 512184 521086 512236 521092
rect 512092 394596 512144 394602
rect 512092 394538 512144 394544
rect 512000 391944 512052 391950
rect 512000 391886 512052 391892
rect 512196 391882 512224 521086
rect 512184 391876 512236 391882
rect 512184 391818 512236 391824
rect 512840 380769 512868 600100
rect 513380 525088 513432 525094
rect 513380 525030 513432 525036
rect 513392 393310 513420 525030
rect 513380 393304 513432 393310
rect 513380 393246 513432 393252
rect 512826 380760 512882 380769
rect 512826 380695 512882 380704
rect 514220 380361 514248 600100
rect 514760 559632 514812 559638
rect 514760 559574 514812 559580
rect 514772 394670 514800 559574
rect 514852 547936 514904 547942
rect 514852 547878 514904 547884
rect 514864 396030 514892 547878
rect 514852 396024 514904 396030
rect 514852 395966 514904 395972
rect 514760 394664 514812 394670
rect 514760 394606 514812 394612
rect 515600 380633 515628 600100
rect 515586 380624 515642 380633
rect 515586 380559 515642 380568
rect 516980 380497 517008 600100
rect 516966 380488 517022 380497
rect 516966 380423 517022 380432
rect 514206 380352 514262 380361
rect 514206 380287 514262 380296
rect 518360 369209 518388 600100
rect 519740 380225 519768 600100
rect 519726 380216 519782 380225
rect 519726 380151 519782 380160
rect 521120 377505 521148 600100
rect 522500 377777 522528 600100
rect 523682 598360 523738 598369
rect 523682 598295 523738 598304
rect 522486 377768 522542 377777
rect 522486 377703 522542 377712
rect 521106 377496 521162 377505
rect 521106 377431 521162 377440
rect 518346 369200 518402 369209
rect 518346 369135 518402 369144
rect 523696 369073 523724 598295
rect 523880 377641 523908 600100
rect 525260 377913 525288 600100
rect 525246 377904 525302 377913
rect 525246 377839 525302 377848
rect 523866 377632 523922 377641
rect 523866 377567 523922 377576
rect 526640 377369 526668 600100
rect 528020 378729 528048 600100
rect 529202 598088 529258 598097
rect 529202 598023 529258 598032
rect 528006 378720 528062 378729
rect 528006 378655 528062 378664
rect 526626 377360 526682 377369
rect 526626 377295 526682 377304
rect 523682 369064 523738 369073
rect 523682 368999 523738 369008
rect 511446 362264 511502 362273
rect 511446 362199 511502 362208
rect 529216 349897 529244 598023
rect 529400 378146 529428 600100
rect 529388 378140 529440 378146
rect 529388 378082 529440 378088
rect 530780 351257 530808 600100
rect 531962 599856 532018 599865
rect 531962 599791 532018 599800
rect 531976 386209 532004 599791
rect 532160 598369 532188 600100
rect 532146 598360 532202 598369
rect 532146 598295 532202 598304
rect 531962 386200 532018 386209
rect 531962 386135 532018 386144
rect 533540 376009 533568 600100
rect 534736 387802 534764 600102
rect 534724 387796 534776 387802
rect 534724 387738 534776 387744
rect 533526 376000 533582 376009
rect 533526 375935 533582 375944
rect 530766 351248 530822 351257
rect 530766 351183 530822 351192
rect 529202 349888 529258 349897
rect 529202 349823 529258 349832
rect 534920 348401 534948 600100
rect 535748 599185 535776 600238
rect 536010 600199 536066 600208
rect 536840 600228 536892 600234
rect 535734 599176 535790 599185
rect 535734 599111 535790 599120
rect 536024 596174 536052 600199
rect 536840 600170 536892 600176
rect 536024 596146 536144 596174
rect 536116 383489 536144 596146
rect 536102 383480 536158 383489
rect 536102 383415 536158 383424
rect 534906 348392 534962 348401
rect 534906 348327 534962 348336
rect 536300 347177 536328 600100
rect 536852 599049 536880 600170
rect 538600 600137 538628 600578
rect 538586 600128 538642 600137
rect 536838 599040 536894 599049
rect 536838 598975 536894 598984
rect 537680 598097 537708 600100
rect 538586 600063 538642 600072
rect 539060 598262 539088 600100
rect 539048 598256 539100 598262
rect 539048 598198 539100 598204
rect 537666 598088 537722 598097
rect 537666 598023 537722 598032
rect 536286 347168 536342 347177
rect 536286 347103 536342 347112
rect 507950 347032 508006 347041
rect 507950 346967 508006 346976
rect 507308 341556 507360 341562
rect 507308 341498 507360 341504
rect 507964 335354 507992 346967
rect 507872 335326 507992 335354
rect 507872 278089 507900 335326
rect 539612 331809 539640 627807
rect 539690 625152 539746 625161
rect 539690 625087 539746 625096
rect 539598 331800 539654 331809
rect 539598 331735 539654 331744
rect 539704 330449 539732 625087
rect 539796 338881 539824 630527
rect 539966 622432 540022 622441
rect 539966 622367 540022 622376
rect 539874 621072 539930 621081
rect 539874 621007 539930 621016
rect 539888 378078 539916 621007
rect 539980 380866 540008 622367
rect 539968 380860 540020 380866
rect 539968 380802 540020 380808
rect 539876 378072 539928 378078
rect 539876 378014 539928 378020
rect 539782 338872 539838 338881
rect 539782 338807 539838 338816
rect 539690 330440 539746 330449
rect 539690 330375 539746 330384
rect 507858 278080 507914 278089
rect 507858 278015 507914 278024
rect 506480 275324 506532 275330
rect 506480 275266 506532 275272
rect 499578 163976 499634 163985
rect 499578 163911 499634 163920
rect 540256 163169 540284 652831
rect 540348 617574 540376 655658
rect 543476 652905 543504 703520
rect 559668 700369 559696 703520
rect 559654 700360 559710 700369
rect 546500 700324 546552 700330
rect 559654 700295 559710 700304
rect 546500 700266 546552 700272
rect 545118 657384 545174 657393
rect 545118 657319 545174 657328
rect 543738 657248 543794 657257
rect 543738 657183 543794 657192
rect 543462 652896 543518 652905
rect 543462 652831 543518 652840
rect 542358 651264 542414 651273
rect 542358 651199 542414 651208
rect 541162 641744 541218 641753
rect 541162 641679 541218 641688
rect 541070 640384 541126 640393
rect 541070 640319 541126 640328
rect 540978 639024 541034 639033
rect 540978 638959 541034 638968
rect 540336 617568 540388 617574
rect 540336 617510 540388 617516
rect 540348 600166 540376 617510
rect 540336 600160 540388 600166
rect 540336 600102 540388 600108
rect 540992 321473 541020 638959
rect 541084 322289 541112 640319
rect 541176 383217 541204 641679
rect 541254 637664 541310 637673
rect 541254 637599 541310 637608
rect 541162 383208 541218 383217
rect 541162 383143 541218 383152
rect 541268 381041 541296 637599
rect 541346 634944 541402 634953
rect 541346 634879 541402 634888
rect 541360 384441 541388 634879
rect 542372 598369 542400 651199
rect 542818 649904 542874 649913
rect 542818 649839 542874 649848
rect 542450 648544 542506 648553
rect 542450 648479 542506 648488
rect 542358 598360 542414 598369
rect 542358 598295 542414 598304
rect 542464 598233 542492 648479
rect 542634 647184 542690 647193
rect 542634 647119 542690 647128
rect 542542 645824 542598 645833
rect 542542 645759 542598 645768
rect 542450 598224 542506 598233
rect 542450 598159 542506 598168
rect 542556 596873 542584 645759
rect 542648 600302 542676 647119
rect 542726 643104 542782 643113
rect 542726 643039 542782 643048
rect 542636 600296 542688 600302
rect 542636 600238 542688 600244
rect 542740 600234 542768 643039
rect 542832 612785 542860 649839
rect 542910 644464 542966 644473
rect 542910 644399 542966 644408
rect 542818 612776 542874 612785
rect 542818 612711 542874 612720
rect 542924 610745 542952 644399
rect 543370 615904 543426 615913
rect 543370 615839 543426 615848
rect 543002 614544 543058 614553
rect 543002 614479 543058 614488
rect 542910 610736 542966 610745
rect 542910 610671 542966 610680
rect 542728 600228 542780 600234
rect 542728 600170 542780 600176
rect 542542 596864 542598 596873
rect 542542 596799 542598 596808
rect 543016 594833 543044 614479
rect 543186 613184 543242 613193
rect 543186 613119 543242 613128
rect 543094 611824 543150 611833
rect 543094 611759 543150 611768
rect 543108 601089 543136 611759
rect 543094 601080 543150 601089
rect 543094 601015 543150 601024
rect 543200 600273 543228 613119
rect 543186 600264 543242 600273
rect 543186 600199 543242 600208
rect 543002 594824 543058 594833
rect 543002 594759 543058 594768
rect 543384 593473 543412 615839
rect 543370 593464 543426 593473
rect 543370 593399 543426 593408
rect 541346 384432 541402 384441
rect 541346 384367 541402 384376
rect 543752 383625 543780 657183
rect 543832 657076 543884 657082
rect 543832 657018 543884 657024
rect 543844 385014 543872 657018
rect 543922 656976 543978 656985
rect 543922 656911 543978 656920
rect 543936 600273 543964 656911
rect 543922 600264 543978 600273
rect 543922 600199 543978 600208
rect 545132 388657 545160 657319
rect 545210 657112 545266 657121
rect 545210 657047 545266 657056
rect 545224 599865 545252 657047
rect 545210 599856 545266 599865
rect 545210 599791 545266 599800
rect 546512 389162 546540 700266
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 546590 657656 546646 657665
rect 546590 657591 546646 657600
rect 546500 389156 546552 389162
rect 546500 389098 546552 389104
rect 545118 388648 545174 388657
rect 545118 388583 545174 388592
rect 543832 385008 543884 385014
rect 543832 384950 543884 384956
rect 546604 384849 546632 657591
rect 546682 657520 546738 657529
rect 546682 657455 546738 657464
rect 546696 384985 546724 657455
rect 547880 657008 547932 657014
rect 547880 656950 547932 656956
rect 546682 384976 546738 384985
rect 546682 384911 546738 384920
rect 546590 384840 546646 384849
rect 546590 384775 546646 384784
rect 547892 383654 547920 656950
rect 547972 656940 548024 656946
rect 547972 656882 548024 656888
rect 547984 384946 548012 656882
rect 580172 617568 580224 617574
rect 580170 617536 580172 617545
rect 580224 617536 580226 617545
rect 580170 617471 580226 617480
rect 547972 384940 548024 384946
rect 547972 384882 548024 384888
rect 547880 383648 547932 383654
rect 543738 383616 543794 383625
rect 547880 383590 547932 383596
rect 543738 383551 543794 383560
rect 541254 381032 541310 381041
rect 541254 380967 541310 380976
rect 580276 373289 580304 697167
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580262 373280 580318 373289
rect 580262 373215 580318 373224
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580368 340270 580396 643991
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580460 353977 580488 590951
rect 580538 537840 580594 537849
rect 580538 537775 580594 537784
rect 580446 353968 580502 353977
rect 580446 353903 580502 353912
rect 580552 351121 580580 537775
rect 580630 431624 580686 431633
rect 580630 431559 580686 431568
rect 580644 356697 580672 431559
rect 580630 356688 580686 356697
rect 580630 356623 580686 356632
rect 580538 351112 580594 351121
rect 580538 351047 580594 351056
rect 580356 340264 580408 340270
rect 580356 340206 580408 340212
rect 580264 339516 580316 339522
rect 580264 339458 580316 339464
rect 580276 325281 580304 339458
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 541070 322280 541126 322289
rect 541070 322215 541126 322224
rect 540978 321464 541034 321473
rect 540978 321399 541034 321408
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 540242 163160 540298 163169
rect 540242 163095 540298 163104
rect 580276 140554 580304 272167
rect 580354 232384 580410 232393
rect 580354 232319 580410 232328
rect 580368 140622 580396 232319
rect 580446 192536 580502 192545
rect 580446 192471 580502 192480
rect 580460 140690 580488 192471
rect 580538 152688 580594 152697
rect 580538 152623 580594 152632
rect 580448 140684 580500 140690
rect 580448 140626 580500 140632
rect 580356 140616 580408 140622
rect 580356 140558 580408 140564
rect 580264 140548 580316 140554
rect 580264 140490 580316 140496
rect 580552 140486 580580 152623
rect 580540 140480 580592 140486
rect 580540 140422 580592 140428
rect 580262 135960 580318 135969
rect 580262 135895 580318 135904
rect 492586 86184 492642 86193
rect 492586 86119 492642 86128
rect 364614 84960 364670 84969
rect 364614 84895 364670 84904
rect 357530 84824 357586 84833
rect 357530 84759 357586 84768
rect 350448 69692 350500 69698
rect 350448 69634 350500 69640
rect 345664 4208 345716 4214
rect 345664 4150 345716 4156
rect 346952 4208 347004 4214
rect 346952 4150 347004 4156
rect 346964 480 346992 4150
rect 350460 480 350488 69634
rect 355322 55856 355378 55865
rect 355322 55791 355378 55800
rect 355336 4865 355364 55791
rect 355322 4856 355378 4865
rect 354036 4820 354088 4826
rect 355322 4791 355378 4800
rect 354036 4762 354088 4768
rect 354048 480 354076 4762
rect 357544 480 357572 84759
rect 361118 84552 361174 84561
rect 361118 84487 361174 84496
rect 361132 480 361160 84487
rect 364628 480 364656 84895
rect 432602 83056 432658 83065
rect 432602 82991 432658 83000
rect 428554 81696 428610 81705
rect 428554 81631 428610 81640
rect 421562 78976 421618 78985
rect 421562 78911 421618 78920
rect 417422 77616 417478 77625
rect 417422 77551 417478 77560
rect 414662 76256 414718 76265
rect 414662 76191 414718 76200
rect 410522 74896 410578 74905
rect 410522 74831 410578 74840
rect 368204 50380 368256 50386
rect 368204 50322 368256 50328
rect 368216 480 368244 50322
rect 400126 40760 400182 40769
rect 400126 40695 400182 40704
rect 393042 24304 393098 24313
rect 393042 24239 393098 24248
rect 382370 20088 382426 20097
rect 382370 20023 382426 20032
rect 378874 13152 378930 13161
rect 378874 13087 378930 13096
rect 375286 11792 375342 11801
rect 375286 11727 375342 11736
rect 371700 3460 371752 3466
rect 371700 3402 371752 3408
rect 371712 480 371740 3402
rect 375300 480 375328 11727
rect 378888 480 378916 13087
rect 382384 480 382412 20023
rect 389454 16008 389510 16017
rect 389454 15943 389510 15952
rect 385958 14648 386014 14657
rect 385958 14583 386014 14592
rect 385972 480 386000 14583
rect 389468 480 389496 15943
rect 393056 480 393084 24239
rect 396538 17368 396594 17377
rect 396538 17303 396594 17312
rect 396552 480 396580 17303
rect 400140 480 400168 40695
rect 403622 39400 403678 39409
rect 403622 39335 403678 39344
rect 403636 480 403664 39335
rect 407210 18728 407266 18737
rect 407210 18663 407266 18672
rect 407224 480 407252 18663
rect 410536 3641 410564 74831
rect 411902 57216 411958 57225
rect 411902 57151 411958 57160
rect 411916 4865 411944 57151
rect 410798 4856 410854 4865
rect 410798 4791 410854 4800
rect 411902 4856 411958 4865
rect 411902 4791 411958 4800
rect 414294 4856 414350 4865
rect 414294 4791 414350 4800
rect 410522 3632 410578 3641
rect 410522 3567 410578 3576
rect 410812 480 410840 4791
rect 414308 480 414336 4791
rect 414676 3097 414704 76191
rect 417436 3505 417464 77551
rect 418802 59936 418858 59945
rect 418802 59871 418858 59880
rect 417882 7576 417938 7585
rect 417882 7511 417938 7520
rect 417422 3496 417478 3505
rect 417422 3431 417478 3440
rect 414662 3088 414718 3097
rect 414662 3023 414718 3032
rect 417896 480 417924 7511
rect 418816 4185 418844 59871
rect 418802 4176 418858 4185
rect 418802 4111 418858 4120
rect 421378 4176 421434 4185
rect 421378 4111 421434 4120
rect 421392 480 421420 4111
rect 421576 3913 421604 78911
rect 425702 68096 425758 68105
rect 425702 68031 425758 68040
rect 422942 61296 422998 61305
rect 422942 61231 422998 61240
rect 422956 4185 422984 61231
rect 425716 7585 425744 68031
rect 427082 62656 427138 62665
rect 427082 62591 427138 62600
rect 425702 7576 425758 7585
rect 425702 7511 425758 7520
rect 427096 4185 427124 62591
rect 422942 4176 422998 4185
rect 422942 4111 422998 4120
rect 424966 4176 425022 4185
rect 424966 4111 425022 4120
rect 427082 4176 427138 4185
rect 427082 4111 427138 4120
rect 428462 4176 428518 4185
rect 428462 4111 428518 4120
rect 421562 3904 421618 3913
rect 421562 3839 421618 3848
rect 424980 480 425008 4111
rect 428476 480 428504 4111
rect 428568 3777 428596 81631
rect 431222 65376 431278 65385
rect 431222 65311 431278 65320
rect 429842 64016 429898 64025
rect 429842 63951 429898 63960
rect 429856 4865 429884 63951
rect 431236 5001 431264 65311
rect 431222 4992 431278 5001
rect 431222 4927 431278 4936
rect 429842 4856 429898 4865
rect 429842 4791 429898 4800
rect 432050 4856 432106 4865
rect 432050 4791 432106 4800
rect 428554 3768 428610 3777
rect 428554 3703 428610 3712
rect 432064 480 432092 4791
rect 432616 3233 432644 82991
rect 450542 73536 450598 73545
rect 450542 73471 450598 73480
rect 446402 72176 446458 72185
rect 446402 72111 446458 72120
rect 443642 70816 443698 70825
rect 443642 70751 443698 70760
rect 436742 66736 436798 66745
rect 436742 66671 436798 66680
rect 435362 47832 435418 47841
rect 435362 47767 435418 47776
rect 435376 4049 435404 47767
rect 435546 4992 435602 5001
rect 435546 4927 435602 4936
rect 435362 4040 435418 4049
rect 435362 3975 435418 3984
rect 432602 3224 432658 3233
rect 432602 3159 432658 3168
rect 435560 480 435588 4927
rect 436756 4185 436784 66671
rect 439502 47696 439558 47705
rect 439502 47631 439558 47640
rect 436742 4176 436798 4185
rect 436742 4111 436798 4120
rect 439134 4176 439190 4185
rect 439134 4111 439190 4120
rect 438858 4040 438914 4049
rect 438858 3975 438914 3984
rect 438872 2854 438900 3975
rect 438860 2848 438912 2854
rect 438860 2790 438912 2796
rect 439148 480 439176 4111
rect 439516 3369 439544 47631
rect 442262 47560 442318 47569
rect 442262 47495 442318 47504
rect 442276 3466 442304 47495
rect 442630 7576 442686 7585
rect 442630 7511 442686 7520
rect 442264 3460 442316 3466
rect 442264 3402 442316 3408
rect 439502 3360 439558 3369
rect 439502 3295 439558 3304
rect 442644 480 442672 7511
rect 443656 4185 443684 70751
rect 446416 4185 446444 72111
rect 450556 4865 450584 73471
rect 580276 73001 580304 135895
rect 580262 72992 580318 73001
rect 580262 72927 580318 72936
rect 471058 51776 471114 51785
rect 471058 51711 471114 51720
rect 450542 4856 450598 4865
rect 450542 4791 450598 4800
rect 453302 4856 453358 4865
rect 453302 4791 453358 4800
rect 443642 4176 443698 4185
rect 443642 4111 443698 4120
rect 446218 4176 446274 4185
rect 446218 4111 446274 4120
rect 446402 4176 446458 4185
rect 446402 4111 446458 4120
rect 449806 4176 449862 4185
rect 449806 4111 449862 4120
rect 446232 480 446260 4111
rect 449820 480 449848 4111
rect 453316 480 453344 4791
rect 467470 3904 467526 3913
rect 467470 3839 467526 3848
rect 456890 3632 456946 3641
rect 456890 3567 456946 3576
rect 456904 480 456932 3567
rect 463974 3496 464030 3505
rect 463974 3431 464030 3440
rect 460386 3088 460442 3097
rect 460386 3023 460442 3032
rect 460400 480 460428 3023
rect 463988 480 464016 3431
rect 467484 480 467512 3839
rect 471072 480 471100 51711
rect 545486 48920 545542 48929
rect 545486 48855 545542 48864
rect 481730 46200 481786 46209
rect 481730 46135 481786 46144
rect 474554 3768 474610 3777
rect 474554 3703 474610 3712
rect 474568 480 474596 3703
rect 478142 3224 478198 3233
rect 478142 3159 478198 3168
rect 478156 480 478184 3159
rect 481744 480 481772 46135
rect 499394 43480 499450 43489
rect 499394 43415 499450 43424
rect 495898 13016 495954 13025
rect 495898 12951 495954 12960
rect 492310 11656 492366 11665
rect 492310 11591 492366 11600
rect 488814 10296 488870 10305
rect 488814 10231 488870 10240
rect 485226 8936 485282 8945
rect 485226 8871 485282 8880
rect 485240 480 485268 8871
rect 488828 480 488856 10231
rect 492324 480 492352 11591
rect 495912 480 495940 12951
rect 499408 480 499436 43415
rect 506478 42120 506534 42129
rect 506478 42055 506534 42064
rect 502982 19952 503038 19961
rect 502982 19887 503038 19896
rect 502996 480 503024 19887
rect 506492 480 506520 42055
rect 512642 40624 512698 40633
rect 512642 40559 512698 40568
rect 508502 14512 508558 14521
rect 508502 14447 508558 14456
rect 508516 4049 508544 14447
rect 508502 4040 508558 4049
rect 508502 3975 508558 3984
rect 510066 4040 510122 4049
rect 510066 3975 510122 3984
rect 510080 480 510108 3975
rect 512656 3505 512684 40559
rect 520738 39264 520794 39273
rect 520738 39199 520794 39208
rect 517150 17232 517206 17241
rect 517150 17167 517206 17176
rect 512642 3496 512698 3505
rect 512642 3431 512698 3440
rect 513562 3496 513618 3505
rect 513562 3431 513618 3440
rect 513576 480 513604 3431
rect 517164 480 517192 17167
rect 520752 480 520780 39199
rect 524234 37904 524290 37913
rect 524234 37839 524290 37848
rect 524248 480 524276 37839
rect 531318 36544 531374 36553
rect 531318 36479 531374 36488
rect 527822 18592 527878 18601
rect 527822 18527 527878 18536
rect 527836 480 527864 18527
rect 531332 480 531360 36479
rect 534906 35184 534962 35193
rect 534906 35119 534962 35128
rect 534920 480 534948 35119
rect 538402 33824 538458 33833
rect 538402 33759 538458 33768
rect 538416 480 538444 33759
rect 541990 30968 542046 30977
rect 541990 30903 542046 30912
rect 542004 480 542032 30903
rect 545500 480 545528 48855
rect 549074 44840 549130 44849
rect 549074 44775 549130 44784
rect 549088 480 549116 44775
rect 552662 29608 552718 29617
rect 552662 29543 552718 29552
rect 552676 480 552704 29543
rect 559746 28248 559802 28257
rect 559746 28183 559802 28192
rect 556158 24168 556214 24177
rect 556158 24103 556214 24112
rect 556172 480 556200 24103
rect 559760 480 559788 28183
rect 562322 26888 562378 26897
rect 562322 26823 562378 26832
rect 562336 3505 562364 26823
rect 566830 25528 566886 25537
rect 566830 25463 566886 25472
rect 562322 3496 562378 3505
rect 562322 3431 562378 3440
rect 563242 3496 563298 3505
rect 563242 3431 563298 3440
rect 563256 480 563284 3431
rect 566844 480 566872 25463
rect 573914 22672 573970 22681
rect 573914 22607 573970 22616
rect 570326 21312 570382 21321
rect 570326 21247 570382 21256
rect 570340 480 570368 21247
rect 573928 480 573956 22607
rect 576122 15872 576178 15881
rect 576122 15807 576178 15816
rect 576136 4049 576164 15807
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 576122 4040 576178 4049
rect 576122 3975 576178 3984
rect 577410 4040 577466 4049
rect 577410 3975 577466 3984
rect 577424 480 577452 3975
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 581000 2848 581052 2854
rect 581000 2790 581052 2796
rect 581012 480 581040 2790
rect 582208 480 582236 3295
rect 583404 480 583432 3402
rect 50130 326 50384 354
rect 50130 -960 50242 326
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 632032 3478 632088
rect 3422 579944 3478 580000
rect 3422 527856 3478 527912
rect 3422 475632 3478 475688
rect 3422 423544 3478 423600
rect 4066 409944 4122 410000
rect 3974 398112 4030 398168
rect 3974 382880 4030 382936
rect 4066 376080 4122 376136
rect 24306 700304 24362 700360
rect 32402 700304 32458 700360
rect 28906 649984 28962 650040
rect 31666 643592 31722 643648
rect 31574 559680 31630 559736
rect 31482 541048 31538 541104
rect 30286 533296 30342 533352
rect 28906 395256 28962 395312
rect 31390 522008 31446 522064
rect 31390 501880 31446 501936
rect 31574 487192 31630 487248
rect 31482 486648 31538 486704
rect 31666 390360 31722 390416
rect 59266 699760 59322 699816
rect 38566 650120 38622 650176
rect 37186 648624 37242 648680
rect 34426 648352 34482 648408
rect 34334 551112 34390 551168
rect 34242 545672 34298 545728
rect 33046 534112 33102 534168
rect 32862 527312 32918 527368
rect 32954 524456 33010 524512
rect 32862 503512 32918 503568
rect 32954 493720 33010 493776
rect 32402 341808 32458 341864
rect 34150 533024 34206 533080
rect 34058 530576 34114 530632
rect 34058 498072 34114 498128
rect 34242 437144 34298 437200
rect 34334 428440 34390 428496
rect 34150 427352 34206 427408
rect 35806 647400 35862 647456
rect 35714 645496 35770 645552
rect 35622 641688 35678 641744
rect 35438 552472 35494 552528
rect 35346 545400 35402 545456
rect 35530 539824 35586 539880
rect 35438 464344 35494 464400
rect 35346 462168 35402 462224
rect 35714 481208 35770 481264
rect 35622 479576 35678 479632
rect 35530 426264 35586 426320
rect 37002 645904 37058 645960
rect 36910 645088 36966 645144
rect 36818 641280 36874 641336
rect 36634 548120 36690 548176
rect 36726 530168 36782 530224
rect 36634 464888 36690 464944
rect 36818 511128 36874 511184
rect 36910 482296 36966 482352
rect 37094 640464 37150 640520
rect 37002 480664 37058 480720
rect 37094 463256 37150 463312
rect 36726 427896 36782 427952
rect 38474 546488 38530 546544
rect 38198 545128 38254 545184
rect 38106 523232 38162 523288
rect 38382 539960 38438 540016
rect 38290 530304 38346 530360
rect 38198 496440 38254 496496
rect 38106 492768 38162 492824
rect 38290 477400 38346 477456
rect 38382 474680 38438 474736
rect 50802 646720 50858 646776
rect 46846 644136 46902 644192
rect 45282 644000 45338 644056
rect 42614 642640 42670 642696
rect 41326 639920 41382 639976
rect 39854 637744 39910 637800
rect 39762 551384 39818 551440
rect 39670 542408 39726 542464
rect 39394 533568 39450 533624
rect 39578 531528 39634 531584
rect 39486 531256 39542 531312
rect 39394 478488 39450 478544
rect 38566 475768 38622 475824
rect 39486 418648 39542 418704
rect 39578 411032 39634 411088
rect 39670 399064 39726 399120
rect 38474 398520 38530 398576
rect 39854 471960 39910 472016
rect 39762 396888 39818 396944
rect 37186 391992 37242 392048
rect 35806 391448 35862 391504
rect 34426 390904 34482 390960
rect 33046 341672 33102 341728
rect 30286 341536 30342 341592
rect 8114 316648 8170 316704
rect 4802 262248 4858 262304
rect 3422 214920 3478 214976
rect 2870 91704 2926 91760
rect 1674 3440 1730 3496
rect 41050 545264 41106 545320
rect 40774 531664 40830 531720
rect 40590 525952 40646 526008
rect 40498 522688 40554 522744
rect 40498 498888 40554 498944
rect 40682 519424 40738 519480
rect 40590 498752 40646 498808
rect 40682 479032 40738 479088
rect 40958 530984 41014 531040
rect 40866 524728 40922 524784
rect 40774 420280 40830 420336
rect 40866 408856 40922 408912
rect 41234 543904 41290 543960
rect 41142 541184 41198 541240
rect 41050 407768 41106 407824
rect 40958 405592 41014 405648
rect 41142 402872 41198 402928
rect 42430 549752 42486 549808
rect 42154 525136 42210 525192
rect 42062 523504 42118 523560
rect 42062 499704 42118 499760
rect 42246 523776 42302 523832
rect 42154 491136 42210 491192
rect 42338 519288 42394 519344
rect 42246 482840 42302 482896
rect 42338 470328 42394 470384
rect 41326 467064 41382 467120
rect 42522 533432 42578 533488
rect 42430 426808 42486 426864
rect 42706 641416 42762 641472
rect 42614 508952 42670 509008
rect 43994 635704 44050 635760
rect 43534 556144 43590 556200
rect 43442 537648 43498 537704
rect 43350 518880 43406 518936
rect 43442 510448 43498 510504
rect 43810 526088 43866 526144
rect 43718 525272 43774 525328
rect 43626 524864 43682 524920
rect 43534 497392 43590 497448
rect 43350 476312 43406 476368
rect 43626 465976 43682 466032
rect 42706 465432 42762 465488
rect 43718 459448 43774 459504
rect 42522 408312 42578 408368
rect 43902 520376 43958 520432
rect 43810 401784 43866 401840
rect 41234 399608 41290 399664
rect 45006 548392 45062 548448
rect 44086 547848 44142 547904
rect 43994 505144 44050 505200
rect 44638 524592 44694 524648
rect 44178 519424 44234 519480
rect 44914 519968 44970 520024
rect 44822 518064 44878 518120
rect 44638 504328 44694 504384
rect 44822 497664 44878 497720
rect 45190 536968 45246 537024
rect 45098 519696 45154 519752
rect 45006 496304 45062 496360
rect 44914 469784 44970 469840
rect 45098 459992 45154 460048
rect 45190 403416 45246 403472
rect 44086 402328 44142 402384
rect 43902 395800 43958 395856
rect 46754 643456 46810 643512
rect 45466 643184 45522 643240
rect 45374 640736 45430 640792
rect 45282 394712 45338 394768
rect 46662 642096 46718 642152
rect 46478 639376 46534 639432
rect 46386 530032 46442 530088
rect 46294 526360 46350 526416
rect 46110 521872 46166 521928
rect 46018 520784 46074 520840
rect 45926 518880 45982 518936
rect 46018 506232 46074 506288
rect 46110 497800 46166 497856
rect 46570 635296 46626 635352
rect 46478 498208 46534 498264
rect 46754 458904 46810 458960
rect 46662 458360 46718 458416
rect 46570 456864 46626 456920
rect 46386 418104 46442 418160
rect 46294 417016 46350 417072
rect 48226 635024 48282 635080
rect 48134 634480 48190 634536
rect 48042 597352 48098 597408
rect 47398 553696 47454 553752
rect 47858 576680 47914 576736
rect 48042 556960 48098 557016
rect 47950 552336 48006 552392
rect 47858 551248 47914 551304
rect 47766 550976 47822 551032
rect 47674 539688 47730 539744
rect 47582 520512 47638 520568
rect 47490 517792 47546 517848
rect 47490 507320 47546 507376
rect 47582 499160 47638 499216
rect 47398 425176 47454 425232
rect 47674 424632 47730 424688
rect 47766 424088 47822 424144
rect 48042 552200 48098 552256
rect 47950 423544 48006 423600
rect 49606 618024 49662 618080
rect 49422 579944 49478 580000
rect 49514 577768 49570 577824
rect 49422 555464 49478 555520
rect 49514 551928 49570 551984
rect 49514 549888 49570 549944
rect 49422 545536 49478 545592
rect 49146 544040 49202 544096
rect 48870 542680 48926 542736
rect 48226 456728 48282 456784
rect 48134 455640 48190 455696
rect 49054 537240 49110 537296
rect 48962 533704 49018 533760
rect 48962 435512 49018 435568
rect 49238 541320 49294 541376
rect 49146 436600 49202 436656
rect 49054 434424 49110 434480
rect 49330 535880 49386 535936
rect 49238 432792 49294 432848
rect 48870 422456 48926 422512
rect 50710 594088 50766 594144
rect 50526 593000 50582 593056
rect 50434 575592 50490 575648
rect 50066 557640 50122 557696
rect 49606 542272 49662 542328
rect 49514 433336 49570 433392
rect 49422 431704 49478 431760
rect 50526 559000 50582 559056
rect 50710 557368 50766 557424
rect 50434 551520 50490 551576
rect 50710 548256 50766 548312
rect 50526 546760 50582 546816
rect 50342 538464 50398 538520
rect 50250 532208 50306 532264
rect 50158 519288 50214 519344
rect 50434 535744 50490 535800
rect 50342 437688 50398 437744
rect 50250 434968 50306 435024
rect 50066 431160 50122 431216
rect 49330 421912 49386 421968
rect 50526 423000 50582 423056
rect 53746 646584 53802 646640
rect 52182 646448 52238 646504
rect 52090 646176 52146 646232
rect 50986 641960 51042 642016
rect 50894 638968 50950 639024
rect 50802 481752 50858 481808
rect 51998 641144 52054 641200
rect 51906 582120 51962 582176
rect 51814 578856 51870 578912
rect 51722 574504 51778 574560
rect 51722 553968 51778 554024
rect 51906 554104 51962 554160
rect 51906 553560 51962 553616
rect 51814 552744 51870 552800
rect 51814 545944 51870 546000
rect 51722 529488 51778 529544
rect 51538 528672 51594 528728
rect 50986 462712 51042 462768
rect 50894 461624 50950 461680
rect 51630 525000 51686 525056
rect 51538 432248 51594 432304
rect 51630 425720 51686 425776
rect 50710 421368 50766 421424
rect 50434 420824 50490 420880
rect 51722 417560 51778 417616
rect 52090 473592 52146 473648
rect 53654 646312 53710 646368
rect 53470 646040 53526 646096
rect 52366 643320 52422 643376
rect 52274 640872 52330 640928
rect 52182 472504 52238 472560
rect 51998 471416 52054 471472
rect 52274 461080 52330 461136
rect 53286 636248 53342 636304
rect 53194 587560 53250 587616
rect 53102 573416 53158 573472
rect 53194 559544 53250 559600
rect 53102 555328 53158 555384
rect 52458 551112 52514 551168
rect 53102 550840 53158 550896
rect 53010 537104 53066 537160
rect 52918 529896 52974 529952
rect 52366 460536 52422 460592
rect 52918 433880 52974 433936
rect 53010 412120 53066 412176
rect 53194 549616 53250 549672
rect 53102 410488 53158 410544
rect 53378 558456 53434 558512
rect 53378 540368 53434 540424
rect 53286 494128 53342 494184
rect 53194 409400 53250 409456
rect 51906 400696 51962 400752
rect 51814 400152 51870 400208
rect 48042 397976 48098 398032
rect 53562 642776 53618 642832
rect 53470 477944 53526 478000
rect 53654 474136 53710 474192
rect 54298 644816 54354 644872
rect 53838 635296 53894 635352
rect 53746 473048 53802 473104
rect 53562 470872 53618 470928
rect 55034 639240 55090 639296
rect 54850 635976 54906 636032
rect 54666 635296 54722 635352
rect 54758 633392 54814 633448
rect 54666 601704 54722 601760
rect 54942 635432 54998 635488
rect 54850 600616 54906 600672
rect 54758 599528 54814 599584
rect 54942 596264 54998 596320
rect 54850 591912 54906 591968
rect 54758 586336 54814 586392
rect 54666 585384 54722 585440
rect 54482 584296 54538 584352
rect 54574 581032 54630 581088
rect 54482 555600 54538 555656
rect 54942 588648 54998 588704
rect 54850 559408 54906 559464
rect 54942 556824 54998 556880
rect 54758 556688 54814 556744
rect 54666 555736 54722 555792
rect 54574 552880 54630 552936
rect 54758 547984 54814 548040
rect 54666 542544 54722 542600
rect 54574 539552 54630 539608
rect 54482 535608 54538 535664
rect 54390 532752 54446 532808
rect 54298 469240 54354 469296
rect 54482 411576 54538 411632
rect 54390 409944 54446 410000
rect 54850 546624 54906 546680
rect 54758 407224 54814 407280
rect 54942 543768 54998 543824
rect 54850 406136 54906 406192
rect 54666 405048 54722 405104
rect 54574 404504 54630 404560
rect 53378 397432 53434 397488
rect 55126 583208 55182 583264
rect 65246 647672 65302 647728
rect 56506 640736 56562 640792
rect 55494 633256 55550 633312
rect 55218 564304 55274 564360
rect 55126 558320 55182 558376
rect 63958 637200 64014 637256
rect 62670 636656 62726 636712
rect 67822 639648 67878 639704
rect 66534 637880 66590 637936
rect 69110 638016 69166 638072
rect 71686 637336 71742 637392
rect 70398 635840 70454 635896
rect 70582 635704 70638 635760
rect 89166 700304 89222 700360
rect 103886 648080 103942 648136
rect 96158 647944 96214 648000
rect 91006 647808 91062 647864
rect 86866 644136 86922 644192
rect 80058 644000 80114 644056
rect 85854 644000 85910 644056
rect 80702 643728 80758 643784
rect 76838 638152 76894 638208
rect 75550 636928 75606 636984
rect 73158 636520 73214 636576
rect 74262 636384 74318 636440
rect 71870 635160 71926 635216
rect 72974 635160 73030 635216
rect 75826 636792 75882 636848
rect 78126 636928 78182 636984
rect 78586 636248 78642 636304
rect 79414 635704 79470 635760
rect 79322 635024 79378 635080
rect 84566 642368 84622 642424
rect 82818 639920 82874 639976
rect 81438 639240 81494 639296
rect 83278 639240 83334 639296
rect 81990 639104 82046 639160
rect 85486 641688 85542 641744
rect 88430 643864 88486 643920
rect 87142 638560 87198 638616
rect 88982 643184 89038 643240
rect 89718 638288 89774 638344
rect 92478 642504 92534 642560
rect 93582 642504 93638 642560
rect 91098 641144 91154 641200
rect 92294 641144 92350 641200
rect 94870 639920 94926 639976
rect 95146 639784 95202 639840
rect 102598 645360 102654 645416
rect 98734 645224 98790 645280
rect 97906 635568 97962 635624
rect 98090 635568 98146 635624
rect 102138 645088 102194 645144
rect 99378 637472 99434 637528
rect 100022 637064 100078 637120
rect 106186 645496 106242 645552
rect 105174 645088 105230 645144
rect 125598 640056 125654 640112
rect 121918 639512 121974 639568
rect 109038 638696 109094 638752
rect 107750 638424 107806 638480
rect 108302 637744 108358 637800
rect 109498 637608 109554 637664
rect 121366 635704 121422 635760
rect 119986 635568 120042 635624
rect 121090 635024 121146 635080
rect 119342 634888 119398 634944
rect 122746 638968 122802 639024
rect 125782 638968 125838 639024
rect 123206 637744 123262 637800
rect 123482 637608 123538 637664
rect 124218 637064 124274 637120
rect 124494 636248 124550 636304
rect 129738 638444 129794 638480
rect 129738 638424 129740 638444
rect 129740 638424 129792 638444
rect 129792 638424 129794 638444
rect 130934 638424 130990 638480
rect 127070 634616 127126 634672
rect 136086 637336 136142 637392
rect 131118 636928 131174 636984
rect 134614 636792 134670 636848
rect 132222 636520 132278 636576
rect 129830 634480 129886 634536
rect 130934 634480 130990 634536
rect 118054 634344 118110 634400
rect 116766 634208 116822 634264
rect 128358 634208 128414 634264
rect 55586 632732 55642 632768
rect 55586 632712 55588 632732
rect 55588 632712 55640 632732
rect 55640 632712 55642 632732
rect 58622 632712 58678 632768
rect 55586 632032 55642 632088
rect 56322 629856 56378 629912
rect 56138 609320 56194 609376
rect 55954 570152 56010 570208
rect 55678 563488 55734 563544
rect 55770 558864 55826 558920
rect 55678 554512 55734 554568
rect 55494 534928 55550 534984
rect 55678 529760 55734 529816
rect 55126 519560 55182 519616
rect 55126 518880 55182 518936
rect 55034 468152 55090 468208
rect 54942 396344 54998 396400
rect 46846 394168 46902 394224
rect 45466 393624 45522 393680
rect 45374 393080 45430 393136
rect 55862 556552 55918 556608
rect 56046 567976 56102 568032
rect 55954 552608 56010 552664
rect 56046 547440 56102 547496
rect 56230 598440 56286 598496
rect 56230 557232 56286 557288
rect 56230 554784 56286 554840
rect 56138 539144 56194 539200
rect 55954 538328 56010 538384
rect 55862 532888 55918 532944
rect 55770 522960 55826 523016
rect 55770 467608 55826 467664
rect 55862 419192 55918 419248
rect 56046 534112 56102 534168
rect 55954 412664 56010 412720
rect 56046 406680 56102 406736
rect 56414 628768 56470 628824
rect 56322 542000 56378 542056
rect 59174 625640 59230 625696
rect 57610 624552 57666 624608
rect 57518 615848 57574 615904
rect 57334 612584 57390 612640
rect 57242 607144 57298 607200
rect 57058 604968 57114 605024
rect 56966 595176 57022 595232
rect 56966 590824 57022 590880
rect 56966 589736 57022 589792
rect 57150 602792 57206 602848
rect 57058 559816 57114 559872
rect 57058 558592 57114 558648
rect 56506 557640 56562 557696
rect 56506 556144 56562 556200
rect 57426 603880 57482 603936
rect 57242 559952 57298 560008
rect 57334 559272 57390 559328
rect 57150 555872 57206 555928
rect 56414 540776 56470 540832
rect 56414 538192 56470 538248
rect 56322 535472 56378 535528
rect 56230 419736 56286 419792
rect 56874 528536 56930 528592
rect 56506 522552 56562 522608
rect 56966 524184 57022 524240
rect 56874 515480 56930 515536
rect 56966 514392 57022 514448
rect 59082 622376 59138 622432
rect 57794 621288 57850 621344
rect 57702 613672 57758 613728
rect 57518 560224 57574 560280
rect 57610 559680 57666 559736
rect 57518 559136 57574 559192
rect 57610 557912 57666 557968
rect 58438 620200 58494 620256
rect 57886 616936 57942 616992
rect 57610 554920 57666 554976
rect 57518 550432 57574 550488
rect 57426 547168 57482 547224
rect 57334 546896 57390 546952
rect 57150 513304 57206 513360
rect 56414 403960 56470 404016
rect 56322 401240 56378 401296
rect 55678 387096 55734 387152
rect 57058 496304 57114 496360
rect 57150 495488 57206 495544
rect 57150 492632 57206 492688
rect 57150 480120 57206 480176
rect 57426 529080 57482 529136
rect 57518 527584 57574 527640
rect 57426 517112 57482 517168
rect 57334 516024 57390 516080
rect 57518 513848 57574 513904
rect 57794 552472 57850 552528
rect 57702 543632 57758 543688
rect 58346 565800 58402 565856
rect 58070 559272 58126 559328
rect 58346 549072 58402 549128
rect 58990 619112 59046 619168
rect 58898 614760 58954 614816
rect 58806 610408 58862 610464
rect 58714 608232 58770 608288
rect 58622 571240 58678 571296
rect 58530 551792 58586 551848
rect 58438 543360 58494 543416
rect 58714 544720 58770 544776
rect 58622 541456 58678 541512
rect 57886 539416 57942 539472
rect 59082 536424 59138 536480
rect 59818 623464 59874 623520
rect 59726 611496 59782 611552
rect 59542 569064 59598 569120
rect 59266 566752 59322 566808
rect 59542 557096 59598 557152
rect 59266 554648 59322 554704
rect 59266 550976 59322 551032
rect 59266 548392 59322 548448
rect 59082 533840 59138 533896
rect 59174 533568 59230 533624
rect 58990 532480 59046 532536
rect 58898 530440 58954 530496
rect 59174 530304 59230 530360
rect 59082 529216 59138 529272
rect 57794 528808 57850 528864
rect 57702 519988 57758 520024
rect 57702 519968 57704 519988
rect 57704 519968 57756 519988
rect 57756 519968 57758 519988
rect 57610 512760 57666 512816
rect 57518 506368 57574 506424
rect 57334 504464 57390 504520
rect 57610 504328 57666 504384
rect 57518 500248 57574 500304
rect 57886 527448 57942 527504
rect 57794 516568 57850 516624
rect 57978 523776 58034 523832
rect 57886 512216 57942 512272
rect 57794 509904 57850 509960
rect 57610 499296 57666 499352
rect 57518 499160 57574 499216
rect 57426 497800 57482 497856
rect 57334 497664 57390 497720
rect 57610 498888 57666 498944
rect 57702 498752 57758 498808
rect 57610 497528 57666 497584
rect 57610 497392 57666 497448
rect 57518 496984 57574 497040
rect 57702 495352 57758 495408
rect 57610 494264 57666 494320
rect 57518 494128 57574 494184
rect 57426 493176 57482 493232
rect 57334 491544 57390 491600
rect 57702 492904 57758 492960
rect 57518 491272 57574 491328
rect 57610 489776 57666 489832
rect 57518 475224 57574 475280
rect 57426 468696 57482 468752
rect 57610 463800 57666 463856
rect 57702 430616 57758 430672
rect 57334 392536 57390 392592
rect 57886 509088 57942 509144
rect 57886 502968 57942 503024
rect 58070 517520 58126 517576
rect 57978 491272 58034 491328
rect 58530 518744 58586 518800
rect 58530 506368 58586 506424
rect 58070 489776 58126 489832
rect 57794 386416 57850 386472
rect 59174 528672 59230 528728
rect 59174 523912 59230 523968
rect 59082 521600 59138 521656
rect 58990 517928 59046 517984
rect 58898 517792 58954 517848
rect 58898 511672 58954 511728
rect 58990 509088 59046 509144
rect 58990 504464 59046 504520
rect 58898 495488 58954 495544
rect 58990 492632 59046 492688
rect 59174 502424 59230 502480
rect 59174 489776 59230 489832
rect 59082 466520 59138 466576
rect 58898 428984 58954 429040
rect 59174 389136 59230 389192
rect 59542 530712 59598 530768
rect 59450 529080 59506 529136
rect 59542 522960 59598 523016
rect 59542 509904 59598 509960
rect 59818 606056 59874 606112
rect 59726 538056 59782 538112
rect 59818 531800 59874 531856
rect 60738 560360 60794 560416
rect 60002 560224 60058 560280
rect 59910 529896 59966 529952
rect 59910 529760 59966 529816
rect 59910 522008 59966 522064
rect 59634 492904 59690 492960
rect 59450 492632 59506 492688
rect 59450 489776 59506 489832
rect 60094 556280 60150 556336
rect 60370 545808 60426 545864
rect 60186 545672 60242 545728
rect 60186 537376 60242 537432
rect 60278 534248 60334 534304
rect 60186 436328 60242 436384
rect 60094 430344 60150 430400
rect 60278 429800 60334 429856
rect 59266 387232 59322 387288
rect 96526 560224 96582 560280
rect 60830 537648 60886 537704
rect 61566 538736 61622 538792
rect 61474 537512 61530 537568
rect 60738 533704 60794 533760
rect 60738 533160 60794 533216
rect 62118 522144 62174 522200
rect 63774 560088 63830 560144
rect 64326 559680 64382 559736
rect 62486 522960 62542 523016
rect 63498 524184 63554 524240
rect 63682 522824 63738 522880
rect 63498 522688 63554 522744
rect 64510 523912 64566 523968
rect 65890 558184 65946 558240
rect 65522 523776 65578 523832
rect 67454 555328 67510 555384
rect 66534 536560 66590 536616
rect 66166 524048 66222 524104
rect 67638 531120 67694 531176
rect 67546 530168 67602 530224
rect 68926 553968 68982 554024
rect 68558 532072 68614 532128
rect 70582 551520 70638 551576
rect 70398 533024 70454 533080
rect 69570 524048 69626 524104
rect 69662 523504 69718 523560
rect 70674 533568 70730 533624
rect 71778 551656 71834 551712
rect 71778 551248 71834 551304
rect 71594 538600 71650 538656
rect 73618 554376 73674 554432
rect 73158 553696 73214 553752
rect 73710 551928 73766 551984
rect 72606 543496 72662 543552
rect 75274 552744 75330 552800
rect 74630 540232 74686 540288
rect 75642 549208 75698 549264
rect 75826 548120 75882 548176
rect 76838 555464 76894 555520
rect 76654 541592 76710 541648
rect 75826 539960 75882 540016
rect 78402 553016 78458 553072
rect 77666 547304 77722 547360
rect 78586 546896 78642 546952
rect 78678 545672 78734 545728
rect 79322 545536 79378 545592
rect 79966 554104 80022 554160
rect 79690 544856 79746 544912
rect 81530 558320 81586 558376
rect 81438 552336 81494 552392
rect 81438 550840 81494 550896
rect 80702 522688 80758 522744
rect 80058 521872 80114 521928
rect 81714 553152 81770 553208
rect 83094 555600 83150 555656
rect 82726 551112 82782 551168
rect 82818 537376 82874 537432
rect 84658 555736 84714 555792
rect 83738 537376 83794 537432
rect 84750 550024 84806 550080
rect 85486 549888 85542 549944
rect 86222 556688 86278 556744
rect 85762 548528 85818 548584
rect 87786 559544 87842 559600
rect 86866 548256 86922 548312
rect 86774 539280 86830 539336
rect 86866 538464 86922 538520
rect 89350 556824 89406 556880
rect 88798 554104 88854 554160
rect 88982 553560 89038 553616
rect 87878 542952 87934 543008
rect 89810 547032 89866 547088
rect 89718 546760 89774 546816
rect 91006 558456 91062 558512
rect 91006 557640 91062 557696
rect 90822 545808 90878 545864
rect 89718 545400 89774 545456
rect 91834 540912 91890 540968
rect 91098 539824 91154 539880
rect 61566 517928 61622 517984
rect 94594 560088 94650 560144
rect 94226 559408 94282 559464
rect 94594 559408 94650 559464
rect 94134 556552 94190 556608
rect 92846 544448 92902 544504
rect 92478 544176 92534 544232
rect 95606 559000 95662 559056
rect 95146 556416 95202 556472
rect 94870 543088 94926 543144
rect 95146 542680 95202 542736
rect 96526 559000 96582 559056
rect 97722 559408 97778 559464
rect 97814 559272 97870 559328
rect 97170 557368 97226 557424
rect 96894 535336 96950 535392
rect 96526 532208 96582 532264
rect 95882 531936 95938 531992
rect 98642 552200 98698 552256
rect 97814 536152 97870 536208
rect 97906 535880 97962 535936
rect 97906 534248 97962 534304
rect 98918 552880 98974 552936
rect 100850 556960 100906 557016
rect 100850 556008 100906 556064
rect 100758 554920 100814 554976
rect 99930 551248 99986 551304
rect 99378 550704 99434 550760
rect 101862 556008 101918 556064
rect 100942 549888 100998 549944
rect 100758 549752 100814 549808
rect 100758 525136 100814 525192
rect 100298 521464 100354 521520
rect 99378 520784 99434 520840
rect 102138 557232 102194 557288
rect 102138 556960 102194 557016
rect 101954 525544 102010 525600
rect 103426 556960 103482 557016
rect 102138 525272 102194 525328
rect 102966 525272 103022 525328
rect 104990 557232 105046 557288
rect 103978 527040 104034 527096
rect 106554 553832 106610 553888
rect 106002 526904 106058 526960
rect 105082 526224 105138 526280
rect 107566 553424 107622 553480
rect 107014 526768 107070 526824
rect 108302 554512 108358 554568
rect 108118 553696 108174 553752
rect 108026 526632 108082 526688
rect 107566 526360 107622 526416
rect 109682 558456 109738 558512
rect 109130 557504 109186 557560
rect 109038 526088 109094 526144
rect 108302 525952 108358 526008
rect 109314 526496 109370 526552
rect 109130 525816 109186 525872
rect 111798 541320 111854 541376
rect 112810 557368 112866 557424
rect 112074 530848 112130 530904
rect 111798 530032 111854 530088
rect 110050 526360 110106 526416
rect 111246 521600 111302 521656
rect 110418 520648 110474 520704
rect 113086 541728 113142 541784
rect 114098 522144 114154 522200
rect 114466 521736 114522 521792
rect 114374 520784 114430 520840
rect 115846 554648 115902 554704
rect 115754 554512 115810 554568
rect 115110 521328 115166 521384
rect 114466 520512 114522 520568
rect 115754 520240 115810 520296
rect 117778 558728 117834 558784
rect 117502 558048 117558 558104
rect 117134 532208 117190 532264
rect 117226 531664 117282 531720
rect 116122 521192 116178 521248
rect 117226 520376 117282 520432
rect 117962 558592 118018 558648
rect 119066 558864 119122 558920
rect 118146 557912 118202 557968
rect 118698 538328 118754 538384
rect 118698 524864 118754 524920
rect 120170 558728 120226 558784
rect 119342 557912 119398 557968
rect 120170 558592 120226 558648
rect 120814 558592 120870 558648
rect 120078 557640 120134 557696
rect 119342 538872 119398 538928
rect 119158 525136 119214 525192
rect 120078 525000 120134 525056
rect 122102 558728 122158 558784
rect 121458 554784 121514 554840
rect 121458 545264 121514 545320
rect 122194 555192 122250 555248
rect 122102 540640 122158 540696
rect 121458 539688 121514 539744
rect 121182 525000 121238 525056
rect 122286 545536 122342 545592
rect 124218 558864 124274 558920
rect 123206 537784 123262 537840
rect 124126 555872 124182 555928
rect 124402 555872 124458 555928
rect 124126 537240 124182 537296
rect 126334 558864 126390 558920
rect 126334 548664 126390 548720
rect 126886 547984 126942 548040
rect 126242 546896 126298 546952
rect 126886 546624 126942 546680
rect 125230 543224 125286 543280
rect 125506 542544 125562 542600
rect 125322 537512 125378 537568
rect 128174 544584 128230 544640
rect 127622 544040 127678 544096
rect 129278 536288 129334 536344
rect 128358 535744 128414 535800
rect 127254 529624 127310 529680
rect 127622 528808 127678 528864
rect 131302 539008 131358 539064
rect 131118 538192 131174 538248
rect 133142 536560 133198 536616
rect 132314 532344 132370 532400
rect 131118 531528 131174 531584
rect 130014 523912 130070 523968
rect 130290 523912 130346 523968
rect 126886 522960 126942 523016
rect 128450 522824 128506 522880
rect 131578 523776 131634 523832
rect 135258 636248 135314 636304
rect 134798 604424 134854 604480
rect 134706 531120 134762 531176
rect 134522 528944 134578 529000
rect 133326 524864 133382 524920
rect 133786 524728 133842 524784
rect 135166 561584 135222 561640
rect 135350 634888 135406 634944
rect 135258 558728 135314 558784
rect 135350 557368 135406 557424
rect 134982 556552 135038 556608
rect 136914 635432 136970 635488
rect 136638 635024 136694 635080
rect 136270 532072 136326 532128
rect 135166 528672 135222 528728
rect 134798 521464 134854 521520
rect 134982 521464 135038 521520
rect 136822 633936 136878 633992
rect 136730 633800 136786 633856
rect 137282 619656 137338 619712
rect 136914 605104 136970 605160
rect 136914 604424 136970 604480
rect 136822 558456 136878 558512
rect 137466 598304 137522 598360
rect 137374 576816 137430 576872
rect 137650 597624 137706 597680
rect 137558 572872 137614 572928
rect 137466 556960 137522 557016
rect 137650 560904 137706 560960
rect 137558 524320 137614 524376
rect 137742 524048 137798 524104
rect 137374 523776 137430 523832
rect 136730 521600 136786 521656
rect 136638 520784 136694 520840
rect 141422 699760 141478 699816
rect 153198 681808 153254 681864
rect 150530 660864 150586 660920
rect 152462 660864 152518 660920
rect 140778 639512 140834 639568
rect 138110 638968 138166 639024
rect 138110 558592 138166 558648
rect 138846 635296 138902 635352
rect 138938 633392 138994 633448
rect 139398 637744 139454 637800
rect 138846 602928 138902 602984
rect 138938 600208 138994 600264
rect 140042 635976 140098 636032
rect 139490 634208 139546 634264
rect 140042 601568 140098 601624
rect 139582 565800 139638 565856
rect 139490 558048 139546 558104
rect 138938 557232 138994 557288
rect 139674 555872 139730 555928
rect 140870 634616 140926 634672
rect 140962 634480 141018 634536
rect 144182 633392 144238 633448
rect 149702 649848 149758 649904
rect 142802 625096 142858 625152
rect 141422 590552 141478 590608
rect 142158 569880 142214 569936
rect 141422 565800 141478 565856
rect 142158 561720 142214 561776
rect 140962 559680 141018 559736
rect 140870 555192 140926 555248
rect 140778 554512 140834 554568
rect 149794 633392 149850 633448
rect 148414 629176 148470 629232
rect 149702 629176 149758 629232
rect 148322 623328 148378 623384
rect 146942 621152 146998 621208
rect 146298 603200 146354 603256
rect 144182 590552 144238 590608
rect 144182 585248 144238 585304
rect 145562 585248 145618 585304
rect 144182 569880 144238 569936
rect 146942 561040 146998 561096
rect 144090 554376 144146 554432
rect 140042 553832 140098 553888
rect 142802 553832 142858 553888
rect 138846 553696 138902 553752
rect 142526 543496 142582 543552
rect 140962 538600 141018 538656
rect 139306 533568 139362 533624
rect 147218 549208 147274 549264
rect 145654 540232 145710 540288
rect 148414 603200 148470 603256
rect 153566 652840 153622 652896
rect 153566 649848 153622 649904
rect 152554 639784 152610 639840
rect 152462 637200 152518 637256
rect 150346 547304 150402 547360
rect 148782 541592 148838 541648
rect 148322 532072 148378 532128
rect 151910 545672 151966 545728
rect 152646 622648 152702 622704
rect 152646 561176 152702 561232
rect 152554 544176 152610 544232
rect 153474 544856 153530 544912
rect 153106 543904 153162 543960
rect 152462 538600 152518 538656
rect 160098 700304 160154 700360
rect 156602 698264 156658 698320
rect 160098 698264 160154 698320
rect 167642 687112 167698 687168
rect 156602 681808 156658 681864
rect 167642 678952 167698 679008
rect 158902 678136 158958 678192
rect 157982 675824 158038 675880
rect 158902 675824 158958 675880
rect 155314 666440 155370 666496
rect 157982 666440 158038 666496
rect 176934 700440 176990 700496
rect 218978 700440 219034 700496
rect 202786 700304 202842 700360
rect 173162 698264 173218 698320
rect 176934 698264 176990 698320
rect 173162 687248 173218 687304
rect 155314 652840 155370 652896
rect 155314 639240 155370 639296
rect 155498 639104 155554 639160
rect 155406 638560 155462 638616
rect 155406 542816 155462 542872
rect 157982 581168 158038 581224
rect 158166 579672 158222 579728
rect 158074 578312 158130 578368
rect 157982 554240 158038 554296
rect 156602 553152 156658 553208
rect 155498 534520 155554 534576
rect 155866 534112 155922 534168
rect 155314 528400 155370 528456
rect 155038 522688 155094 522744
rect 158350 576816 158406 576872
rect 158166 555464 158222 555520
rect 158074 552744 158130 552800
rect 158534 575456 158590 575512
rect 158350 551928 158406 551984
rect 158534 551656 158590 551712
rect 158166 551112 158222 551168
rect 159454 636384 159510 636440
rect 160834 594768 160890 594824
rect 160742 593408 160798 593464
rect 159546 581032 159602 581088
rect 160926 592048 160982 592104
rect 161110 590688 161166 590744
rect 161018 575592 161074 575648
rect 160926 560224 160982 560280
rect 160742 559408 160798 559464
rect 159546 553016 159602 553072
rect 161202 570424 161258 570480
rect 161110 560088 161166 560144
rect 161018 551520 161074 551576
rect 161294 550024 161350 550080
rect 161202 546624 161258 546680
rect 159454 544992 159510 545048
rect 159730 537376 159786 537432
rect 163594 636520 163650 636576
rect 162214 624280 162270 624336
rect 163502 625912 163558 625968
rect 162766 548528 162822 548584
rect 162214 533704 162270 533760
rect 164882 619384 164938 619440
rect 163778 590960 163834 591016
rect 163686 568792 163742 568848
rect 163594 552336 163650 552392
rect 163502 534384 163558 534440
rect 163870 589328 163926 589384
rect 163962 588240 164018 588296
rect 164054 574504 164110 574560
rect 163962 556824 164018 556880
rect 164054 553968 164110 554024
rect 164422 539280 164478 539336
rect 164146 535336 164202 535392
rect 164146 519696 164202 519752
rect 164330 519696 164386 519752
rect 169022 618568 169078 618624
rect 166354 616936 166410 616992
rect 166262 612856 166318 612912
rect 164974 601432 165030 601488
rect 165986 542952 166042 543008
rect 164974 537512 165030 537568
rect 164882 527856 164938 527912
rect 167642 616120 167698 616176
rect 166446 596536 166502 596592
rect 166354 555464 166410 555520
rect 166538 585384 166594 585440
rect 166998 582120 167054 582176
rect 166998 581168 167054 581224
rect 166906 575320 166962 575376
rect 166722 573416 166778 573472
rect 166630 556688 166686 556744
rect 166538 555736 166594 555792
rect 166814 559544 166870 559600
rect 166906 556688 166962 556744
rect 166722 555328 166778 555384
rect 167550 554104 167606 554160
rect 166446 541592 166502 541648
rect 166998 532888 167054 532944
rect 166262 529352 166318 529408
rect 166262 528672 166318 528728
rect 167734 603880 167790 603936
rect 167642 542952 167698 543008
rect 167918 597352 167974 597408
rect 167826 595720 167882 595776
rect 167734 540232 167790 540288
rect 168286 582120 168342 582176
rect 168194 579672 168250 579728
rect 168010 574368 168066 574424
rect 168010 556824 168066 556880
rect 168194 553016 168250 553072
rect 168286 550568 168342 550624
rect 167918 548528 167974 548584
rect 169298 608776 169354 608832
rect 169206 603064 169262 603120
rect 169114 583752 169170 583808
rect 169114 555600 169170 555656
rect 169114 547032 169170 547088
rect 167826 533568 167882 533624
rect 170494 605512 170550 605568
rect 170402 594904 170458 594960
rect 169758 593000 169814 593056
rect 169758 592048 169814 592104
rect 169390 582392 169446 582448
rect 169758 578856 169814 578912
rect 170310 578856 170366 578912
rect 169758 578312 169814 578368
rect 170218 575592 170274 575648
rect 169482 572872 169538 572928
rect 169390 558320 169446 558376
rect 169482 556960 169538 557016
rect 169758 553152 169814 553208
rect 170218 551928 170274 551984
rect 169758 549616 169814 549672
rect 170310 549208 170366 549264
rect 169298 545672 169354 545728
rect 170586 599800 170642 599856
rect 170678 597352 170734 597408
rect 170954 593272 171010 593328
rect 170862 589192 170918 589248
rect 170770 569608 170826 569664
rect 170678 556008 170734 556064
rect 170586 550024 170642 550080
rect 170678 545808 170734 545864
rect 170494 537240 170550 537296
rect 170402 528128 170458 528184
rect 169206 527992 169262 528048
rect 169758 527856 169814 527912
rect 169758 523368 169814 523424
rect 171046 593000 171102 593056
rect 171046 558728 171102 558784
rect 170954 556552 171010 556608
rect 170862 546216 170918 546272
rect 171046 537376 171102 537432
rect 170770 524184 170826 524240
rect 204902 648352 204958 648408
rect 193034 648216 193090 648272
rect 176658 643612 176714 643648
rect 176658 643592 176660 643612
rect 176660 643592 176712 643612
rect 176712 643592 176714 643612
rect 177670 643592 177726 643648
rect 177578 637064 177634 637120
rect 176566 636792 176622 636848
rect 174542 621832 174598 621888
rect 173254 617752 173310 617808
rect 171782 614488 171838 614544
rect 173162 607144 173218 607200
rect 171874 606328 171930 606384
rect 171966 600616 172022 600672
rect 172334 595176 172390 595232
rect 172058 591640 172114 591696
rect 171966 544856 172022 544912
rect 172242 586336 172298 586392
rect 172150 572056 172206 572112
rect 172150 557232 172206 557288
rect 172426 586744 172482 586800
rect 172334 561584 172390 561640
rect 172242 554512 172298 554568
rect 172518 577768 172574 577824
rect 172518 576816 172574 576872
rect 173070 557368 173126 557424
rect 172978 554376 173034 554432
rect 172426 543768 172482 543824
rect 172518 542952 172574 543008
rect 172518 541184 172574 541240
rect 172150 540912 172206 540968
rect 172058 537648 172114 537704
rect 171782 537104 171838 537160
rect 171782 536696 171838 536752
rect 172334 540912 172390 540968
rect 174358 593408 174414 593464
rect 173806 591912 173862 591968
rect 173438 590008 173494 590064
rect 173346 588376 173402 588432
rect 173254 551112 173310 551168
rect 173530 581848 173586 581904
rect 173438 547304 173494 547360
rect 173622 576136 173678 576192
rect 173530 543496 173586 543552
rect 173346 542136 173402 542192
rect 173806 590688 173862 590744
rect 173806 587560 173862 587616
rect 173714 560088 173770 560144
rect 174450 583752 174506 583808
rect 174358 559408 174414 559464
rect 174450 557640 174506 557696
rect 173806 556008 173862 556064
rect 173806 552744 173862 552800
rect 173806 547712 173862 547768
rect 173714 544448 173770 544504
rect 173622 539280 173678 539336
rect 173162 531120 173218 531176
rect 172426 526088 172482 526144
rect 174634 610408 174690 610464
rect 173990 536696 174046 536752
rect 174818 609592 174874 609648
rect 174726 587424 174782 587480
rect 177578 626728 177634 626784
rect 179326 643184 179382 643240
rect 177762 633256 177818 633312
rect 177946 641688 178002 641744
rect 179326 641688 179382 641744
rect 184294 639104 184350 639160
rect 179050 635568 179106 635624
rect 177946 634616 178002 634672
rect 177854 631080 177910 631136
rect 178958 633528 179014 633584
rect 177946 627816 178002 627872
rect 177670 625640 177726 625696
rect 177302 612720 177358 612776
rect 177210 610680 177266 610736
rect 176566 602928 176622 602984
rect 176198 602248 176254 602304
rect 175922 598984 175978 599040
rect 175094 593952 175150 594008
rect 174910 590824 174966 590880
rect 174818 555600 174874 555656
rect 175002 581304 175058 581360
rect 174910 544448 174966 544504
rect 175830 585384 175886 585440
rect 175738 576680 175794 576736
rect 175738 575456 175794 575512
rect 175462 571240 175518 571296
rect 175370 561040 175426 561096
rect 175186 560224 175242 560280
rect 175002 536560 175058 536616
rect 175278 544856 175334 544912
rect 175278 542408 175334 542464
rect 174726 528264 174782 528320
rect 175186 527584 175242 527640
rect 175186 525680 175242 525736
rect 174542 522960 174598 523016
rect 175830 559136 175886 559192
rect 175830 553152 175886 553208
rect 175738 544856 175794 544912
rect 175830 532752 175886 532808
rect 175830 527448 175886 527504
rect 176014 584160 176070 584216
rect 175922 524592 175978 524648
rect 176106 582664 176162 582720
rect 176566 601840 176622 601896
rect 176566 589736 176622 589792
rect 176566 589328 176622 589384
rect 176474 585928 176530 585984
rect 176290 579400 176346 579456
rect 176198 553152 176254 553208
rect 176382 575456 176438 575512
rect 176382 560496 176438 560552
rect 176474 559680 176530 559736
rect 177118 569880 177174 569936
rect 176566 558592 176622 558648
rect 177946 611632 178002 611688
rect 177670 611360 177726 611416
rect 177394 607008 177450 607064
rect 177578 607008 177634 607064
rect 177578 601704 177634 601760
rect 176290 533976 176346 534032
rect 177854 609728 177910 609784
rect 177762 604424 177818 604480
rect 177486 529352 177542 529408
rect 176106 525408 176162 525464
rect 176934 522960 176990 523016
rect 177578 522960 177634 523016
rect 176014 522688 176070 522744
rect 175922 522144 175978 522200
rect 175922 520784 175978 520840
rect 177670 522144 177726 522200
rect 178682 607960 178738 608016
rect 178038 601568 178094 601624
rect 178038 600616 178094 600672
rect 178590 590824 178646 590880
rect 178406 572328 178462 572384
rect 178498 561176 178554 561232
rect 178406 558184 178462 558240
rect 178038 556552 178094 556608
rect 178406 555872 178462 555928
rect 178038 550976 178094 551032
rect 178038 535608 178094 535664
rect 178038 531392 178094 531448
rect 178038 523232 178094 523288
rect 179234 635432 179290 635488
rect 179142 634480 179198 634536
rect 179050 600616 179106 600672
rect 178958 599528 179014 599584
rect 179142 598440 179198 598496
rect 179326 635296 179382 635352
rect 183190 637744 183246 637800
rect 202050 647536 202106 647592
rect 199750 640056 199806 640112
rect 197266 638968 197322 639024
rect 195886 637608 195942 637664
rect 198646 639512 198702 639568
rect 201130 635704 201186 635760
rect 208398 648216 208454 648272
rect 202786 647420 202842 647456
rect 202786 647400 202788 647420
rect 202788 647400 202840 647420
rect 202840 647400 202842 647420
rect 204626 647264 204682 647320
rect 208490 647400 208546 647456
rect 204166 643592 204222 643648
rect 203798 643184 203854 643240
rect 207478 643592 207534 643648
rect 207018 643184 207074 643240
rect 206374 639920 206430 639976
rect 212354 646856 212410 646912
rect 210146 638560 210202 638616
rect 211066 637744 211122 637800
rect 212446 646720 212502 646776
rect 283838 681672 283894 681728
rect 288346 681672 288402 681728
rect 288346 678680 288402 678736
rect 290462 678680 290518 678736
rect 290462 657736 290518 657792
rect 309782 657736 309838 657792
rect 235170 657464 235226 657520
rect 280802 648080 280858 648136
rect 275282 647672 275338 647728
rect 233146 647536 233202 647592
rect 233422 647536 233478 647592
rect 216218 645496 216274 645552
rect 215298 644816 215354 644872
rect 214562 640328 214618 640384
rect 215206 640328 215262 640384
rect 213826 639240 213882 639296
rect 213826 639104 213882 639160
rect 218058 641416 218114 641472
rect 216770 640328 216826 640384
rect 217966 640736 218022 640792
rect 219070 640600 219126 640656
rect 220358 639240 220414 639296
rect 220726 638968 220782 639024
rect 221830 636520 221886 636576
rect 227718 645496 227774 645552
rect 231766 644952 231822 645008
rect 227810 644816 227866 644872
rect 223486 642776 223542 642832
rect 222934 641824 222990 641880
rect 224314 637744 224370 637800
rect 224222 637608 224278 637664
rect 225694 636248 225750 636304
rect 232042 644952 232098 645008
rect 230386 640736 230442 640792
rect 230662 640736 230718 640792
rect 226338 635044 226394 635080
rect 226338 635024 226340 635044
rect 226340 635024 226392 635044
rect 226392 635024 226394 635044
rect 226476 634888 226532 634944
rect 229558 637608 229614 637664
rect 230386 638560 230442 638616
rect 233882 643592 233938 643648
rect 234526 643592 234582 643648
rect 234618 639512 234674 639568
rect 235906 639512 235962 639568
rect 244278 635704 244334 635760
rect 245014 637200 245070 637256
rect 249614 637200 249670 637256
rect 248786 636248 248842 636304
rect 251086 640056 251142 640112
rect 250994 639784 251050 639840
rect 250994 638424 251050 638480
rect 254582 636656 254638 636712
rect 252466 636112 252522 636168
rect 252466 635024 252522 635080
rect 241932 634208 241988 634264
rect 179326 605104 179382 605160
rect 179234 597352 179290 597408
rect 179326 596264 179382 596320
rect 179234 592456 179290 592512
rect 179142 585112 179198 585168
rect 178866 583480 178922 583536
rect 178774 577632 178830 577688
rect 179050 580216 179106 580272
rect 178958 578584 179014 578640
rect 179326 588648 179382 588704
rect 179234 560224 179290 560280
rect 179142 551656 179198 551712
rect 179050 536696 179106 536752
rect 179878 581032 179934 581088
rect 179878 574504 179934 574560
rect 179786 573416 179842 573472
rect 179602 562128 179658 562184
rect 179418 561584 179474 561640
rect 179510 559544 179566 559600
rect 179326 556552 179382 556608
rect 179418 552064 179474 552120
rect 179418 549480 179474 549536
rect 179694 560904 179750 560960
rect 178958 532616 179014 532672
rect 178774 524048 178830 524104
rect 179786 552744 179842 552800
rect 262862 636248 262918 636304
rect 256146 635840 256202 635896
rect 255962 635160 256018 635216
rect 254582 561584 254638 561640
rect 229742 560496 229798 560552
rect 179970 555736 180026 555792
rect 179878 549752 179934 549808
rect 180062 532072 180118 532128
rect 179694 521600 179750 521656
rect 183190 553832 183246 553888
rect 181626 533704 181682 533760
rect 180246 525680 180302 525736
rect 184754 534384 184810 534440
rect 185582 534384 185638 534440
rect 184570 533704 184626 533760
rect 190918 553832 190974 553888
rect 187882 543088 187938 543144
rect 186226 521464 186282 521520
rect 191010 536152 191066 536208
rect 189446 531936 189502 531992
rect 192574 552880 192630 552936
rect 191746 533704 191802 533760
rect 191930 533704 191986 533760
rect 192666 536152 192722 536208
rect 194138 551248 194194 551304
rect 193678 535336 193734 535392
rect 195702 549888 195758 549944
rect 194506 534384 194562 534440
rect 200762 543088 200818 543144
rect 198738 531936 198794 531992
rect 197726 531664 197782 531720
rect 200394 527040 200450 527096
rect 197266 525544 197322 525600
rect 198830 525272 198886 525328
rect 206098 551248 206154 551304
rect 204810 550160 204866 550216
rect 205638 536152 205694 536208
rect 206834 536152 206890 536208
rect 212446 535336 212502 535392
rect 211894 534384 211950 534440
rect 214470 541728 214526 541784
rect 213918 541320 213974 541376
rect 212906 532072 212962 532128
rect 213826 531664 213882 531720
rect 211066 531392 211122 531448
rect 211066 531256 211122 531312
rect 212906 530848 212962 530904
rect 203522 526904 203578 526960
rect 201958 526224 202014 526280
rect 201774 526088 201830 526144
rect 205086 526768 205142 526824
rect 206650 526632 206706 526688
rect 208214 526496 208270 526552
rect 209686 526360 209742 526416
rect 211066 524864 211122 524920
rect 211066 521464 211122 521520
rect 214930 526496 214986 526552
rect 216954 547032 217010 547088
rect 216678 546488 216734 546544
rect 218058 536152 218114 536208
rect 218978 536152 219034 536208
rect 218702 532344 218758 532400
rect 217966 526360 218022 526416
rect 220726 532208 220782 532264
rect 219990 527856 220046 527912
rect 220634 527312 220690 527368
rect 217506 521328 217562 521384
rect 218702 521328 218758 521384
rect 215942 520784 215998 520840
rect 219070 521192 219126 521248
rect 221002 530848 221058 530904
rect 223026 545808 223082 545864
rect 223486 545128 223542 545184
rect 224958 550160 225014 550216
rect 225050 549888 225106 549944
rect 224038 541728 224094 541784
rect 224222 541048 224278 541104
rect 225418 540640 225474 540696
rect 222290 538872 222346 538928
rect 222014 526632 222070 526688
rect 223854 525136 223910 525192
rect 228362 558456 228418 558512
rect 229374 552472 229430 552528
rect 229742 546760 229798 546816
rect 228546 545536 228602 545592
rect 227074 538464 227130 538520
rect 226982 525000 227038 525056
rect 230386 547576 230442 547632
rect 230386 543088 230442 543144
rect 230662 543088 230718 543144
rect 230110 537784 230166 537840
rect 231674 548664 231730 548720
rect 231214 543224 231270 543280
rect 231122 525136 231178 525192
rect 231214 521192 231270 521248
rect 233054 550160 233110 550216
rect 233146 549344 233202 549400
rect 233882 546896 233938 546952
rect 232134 541864 232190 541920
rect 233146 541320 233202 541376
rect 238206 548664 238262 548720
rect 237930 544584 237986 544640
rect 237194 543224 237250 543280
rect 236182 537784 236238 537840
rect 236366 529624 236422 529680
rect 235170 526768 235226 526824
rect 234158 525000 234214 525056
rect 233146 521192 233202 521248
rect 233882 521192 233938 521248
rect 234710 521192 234766 521248
rect 239218 540640 239274 540696
rect 241426 551520 241482 551576
rect 241610 551520 241666 551576
rect 240782 539008 240838 539064
rect 240230 538872 240286 538928
rect 239494 536288 239550 536344
rect 238758 521328 238814 521384
rect 238758 520784 238814 520840
rect 243266 535336 243322 535392
rect 243542 534384 243598 534440
rect 242254 529624 242310 529680
rect 244370 533704 244426 533760
rect 245290 533704 245346 533760
rect 246394 547168 246450 547224
rect 246302 526904 246358 526960
rect 244278 525272 244334 525328
rect 241058 523912 241114 523968
rect 240782 521464 240838 521520
rect 242530 521464 242586 521520
rect 246394 521464 246450 521520
rect 245658 521192 245714 521248
rect 244094 520784 244150 520840
rect 247406 547168 247462 547224
rect 248878 547440 248934 547496
rect 248326 532208 248382 532264
rect 249338 544584 249394 544640
rect 250442 557096 250498 557152
rect 250350 530304 250406 530360
rect 253202 559952 253258 560008
rect 252466 554104 252522 554160
rect 252006 552608 252062 552664
rect 251362 537920 251418 537976
rect 251086 531256 251142 531312
rect 252466 536968 252522 537024
rect 253570 541456 253626 541512
rect 253386 536288 253442 536344
rect 253202 520784 253258 520840
rect 255134 533160 255190 533216
rect 257986 594768 258042 594824
rect 257894 574096 257950 574152
rect 257894 539008 257950 539064
rect 256698 538464 256754 538520
rect 258722 559816 258778 559872
rect 257986 523912 258042 523968
rect 256146 521328 256202 521384
rect 255962 521192 256018 521248
rect 258446 521600 258502 521656
rect 258722 521600 258778 521656
rect 261390 549072 261446 549128
rect 262862 549072 262918 549128
rect 270774 551792 270830 551848
rect 269118 551112 269174 551168
rect 269762 543632 269818 543688
rect 264334 539416 264390 539472
rect 267646 531800 267702 531856
rect 265990 521600 266046 521656
rect 264426 521464 264482 521520
rect 264610 521464 264666 521520
rect 269210 520784 269266 520840
rect 269026 518764 269082 518800
rect 269026 518744 269028 518764
rect 269028 518744 269080 518764
rect 269080 518744 269082 518764
rect 269762 520648 269818 520704
rect 270406 519288 270462 519344
rect 273902 544720 273958 544776
rect 272522 539552 272578 539608
rect 272338 539144 272394 539200
rect 278318 645360 278374 645416
rect 275466 645224 275522 645280
rect 275190 523504 275246 523560
rect 274638 523096 274694 523152
rect 276662 644000 276718 644056
rect 275926 555192 275982 555248
rect 275466 553560 275522 553616
rect 275558 550432 275614 550488
rect 275466 538056 275522 538112
rect 278226 642504 278282 642560
rect 276754 641144 276810 641200
rect 278042 638016 278098 638072
rect 276754 544720 276810 544776
rect 277306 571240 277362 571296
rect 277306 560360 277362 560416
rect 276662 539144 276718 539200
rect 279514 642368 279570 642424
rect 279422 638152 279478 638208
rect 278686 552472 278742 552528
rect 278318 552200 278374 552256
rect 278686 549072 278742 549128
rect 278226 548392 278282 548448
rect 279606 638288 279662 638344
rect 279790 633936 279846 633992
rect 279882 582120 279938 582176
rect 280158 558048 280214 558104
rect 279882 550568 279938 550624
rect 279606 548256 279662 548312
rect 280066 547848 280122 547904
rect 286322 647944 286378 648000
rect 282182 645088 282238 645144
rect 280802 537240 280858 537296
rect 279514 535200 279570 535256
rect 281446 615848 281502 615904
rect 281446 558048 281502 558104
rect 282550 581032 282606 581088
rect 282458 579944 282514 580000
rect 282274 578856 282330 578912
rect 282182 553696 282238 553752
rect 282366 576680 282422 576736
rect 282274 549208 282330 549264
rect 282734 577768 282790 577824
rect 282642 575592 282698 575648
rect 282550 555736 282606 555792
rect 282458 553016 282514 553072
rect 282734 554376 282790 554432
rect 282642 551928 282698 551984
rect 282366 546760 282422 546816
rect 280066 530440 280122 530496
rect 279422 527448 279478 527504
rect 279974 527176 280030 527232
rect 278042 521464 278098 521520
rect 275558 520784 275614 520840
rect 278502 520648 278558 520704
rect 283194 521600 283250 521656
rect 282918 519152 282974 519208
rect 284206 558864 284262 558920
rect 285218 594088 285274 594144
rect 285126 593000 285182 593056
rect 284850 542272 284906 542328
rect 285402 591912 285458 591968
rect 285494 589736 285550 589792
rect 285402 560088 285458 560144
rect 285218 559408 285274 559464
rect 285126 558728 285182 558784
rect 285586 574504 285642 574560
rect 285494 558592 285550 558648
rect 289266 647808 289322 647864
rect 287794 643864 287850 643920
rect 287702 639648 287758 639704
rect 286966 583752 287022 583808
rect 286322 551792 286378 551848
rect 285586 549752 285642 549808
rect 286414 532480 286470 532536
rect 286322 527584 286378 527640
rect 286874 527040 286930 527096
rect 287978 588648 288034 588704
rect 287886 586336 287942 586392
rect 288070 587560 288126 587616
rect 287978 556552 288034 556608
rect 288254 585384 288310 585440
rect 288346 573416 288402 573472
rect 288254 559136 288310 559192
rect 288070 556008 288126 556064
rect 287886 554512 287942 554568
rect 288346 552744 288402 552800
rect 287978 543360 288034 543416
rect 287794 541456 287850 541512
rect 287702 521056 287758 521112
rect 298006 644544 298062 644600
rect 291842 643728 291898 643784
rect 289266 544040 289322 544096
rect 290554 584296 290610 584352
rect 290646 583208 290702 583264
rect 290554 557640 290610 557696
rect 291014 578176 291070 578232
rect 290738 572328 290794 572384
rect 290646 557368 290702 557424
rect 290738 555872 290794 555928
rect 289726 530440 289782 530496
rect 289726 529352 289782 529408
rect 291750 553152 291806 553208
rect 297454 643456 297510 643512
rect 297362 641008 297418 641064
rect 294602 637880 294658 637936
rect 291934 635568 291990 635624
rect 293866 617752 293922 617808
rect 293774 612720 293830 612776
rect 291934 600616 291990 600672
rect 292394 579536 292450 579592
rect 292302 572872 292358 572928
rect 292210 572736 292266 572792
rect 291106 536424 291162 536480
rect 289726 527040 289782 527096
rect 289450 520784 289506 520840
rect 290922 520104 290978 520160
rect 291014 519016 291070 519072
rect 291842 536832 291898 536888
rect 291842 535880 291898 535936
rect 292210 558728 292266 558784
rect 292302 540504 292358 540560
rect 292486 578176 292542 578232
rect 292394 538056 292450 538112
rect 293682 574096 293738 574152
rect 293682 542272 293738 542328
rect 293774 536424 293830 536480
rect 292578 535472 292634 535528
rect 292670 529760 292726 529816
rect 292578 523504 292634 523560
rect 292486 523368 292542 523424
rect 291934 519832 291990 519888
rect 291842 518916 291844 518936
rect 291844 518916 291896 518936
rect 291896 518916 291898 518936
rect 291842 518880 291898 518916
rect 293958 554648 294014 554704
rect 293958 544176 294014 544232
rect 293866 523640 293922 523696
rect 293958 522144 294014 522200
rect 295062 636792 295118 636848
rect 294694 635432 294750 635488
rect 294878 635296 294934 635352
rect 294786 634480 294842 634536
rect 294786 598440 294842 598496
rect 294694 597352 294750 597408
rect 294970 633528 295026 633584
rect 295062 601704 295118 601760
rect 294970 599528 295026 599584
rect 295062 597488 295118 597544
rect 294878 596264 294934 596320
rect 295246 592048 295302 592104
rect 295154 571376 295210 571432
rect 295062 550432 295118 550488
rect 295154 522280 295210 522336
rect 295338 552200 295394 552256
rect 295798 533840 295854 533896
rect 295338 531256 295394 531312
rect 295246 522144 295302 522200
rect 294602 521600 294658 521656
rect 296718 628904 296774 628960
rect 297638 642096 297694 642152
rect 297454 633256 297510 633312
rect 297362 627816 297418 627872
rect 297178 626728 297234 626784
rect 297730 639376 297786 639432
rect 297638 632168 297694 632224
rect 297914 634752 297970 634808
rect 297730 631080 297786 631136
rect 297546 625640 297602 625696
rect 297546 624552 297602 624608
rect 297454 620200 297510 620256
rect 297362 618024 297418 618080
rect 296626 590552 296682 590608
rect 296534 585112 296590 585168
rect 296350 575456 296406 575512
rect 296442 568656 296498 568712
rect 296350 555872 296406 555928
rect 296442 535064 296498 535120
rect 296534 533840 296590 533896
rect 296718 567976 296774 568032
rect 296626 530440 296682 530496
rect 298006 629992 298062 630048
rect 297914 622376 297970 622432
rect 297638 619112 297694 619168
rect 298006 614760 298062 614816
rect 298006 612584 298062 612640
rect 298006 610408 298062 610464
rect 297822 608232 297878 608288
rect 297730 606056 297786 606112
rect 298006 595176 298062 595232
rect 298006 590824 298062 590880
rect 297914 569064 297970 569120
rect 298006 561312 298062 561368
rect 300122 657600 300178 657656
rect 413650 700440 413706 700496
rect 397458 700304 397514 700360
rect 309782 650256 309838 650312
rect 312910 650256 312966 650312
rect 340050 650120 340106 650176
rect 333610 646584 333666 646640
rect 332322 646448 332378 646504
rect 312910 645088 312966 645144
rect 331862 645088 331918 645144
rect 303986 643320 304042 643376
rect 309138 641960 309194 642016
rect 305274 640872 305330 640928
rect 310426 640464 310482 640520
rect 331862 636112 331918 636168
rect 336186 646312 336242 646368
rect 334898 646176 334954 646232
rect 335174 636112 335230 636168
rect 368386 649984 368442 650040
rect 360658 648624 360714 648680
rect 345202 646040 345258 646096
rect 351642 645904 351698 645960
rect 358726 639784 358782 639840
rect 358726 636792 358782 636848
rect 370962 636792 371018 636848
rect 335174 634480 335230 634536
rect 375378 619384 375434 619440
rect 374550 616664 374606 616720
rect 299294 608504 299350 608560
rect 299202 591368 299258 591424
rect 299110 570016 299166 570072
rect 299202 554512 299258 554568
rect 299386 604424 299442 604480
rect 299294 553832 299350 553888
rect 299294 553308 299350 553344
rect 299294 553288 299296 553308
rect 299296 553288 299348 553308
rect 299348 553288 299350 553308
rect 299294 553152 299350 553208
rect 298926 546352 298982 546408
rect 299110 546352 299166 546408
rect 297362 522552 297418 522608
rect 299846 570016 299902 570072
rect 299754 561584 299810 561640
rect 299386 524456 299442 524512
rect 299294 523504 299350 523560
rect 299386 523368 299442 523424
rect 300490 540776 300546 540832
rect 299846 520920 299902 520976
rect 300766 526088 300822 526144
rect 303250 551384 303306 551440
rect 302054 542000 302110 542056
rect 304538 540368 304594 540424
rect 308310 552336 308366 552392
rect 306746 534928 306802 534984
rect 309598 545944 309654 546000
rect 311438 538600 311494 538656
rect 319718 530984 319774 531040
rect 314474 521600 314530 521656
rect 317602 521464 317658 521520
rect 316038 521056 316094 521112
rect 319166 521328 319222 521384
rect 323950 544992 324006 545048
rect 322294 521192 322350 521248
rect 324778 533432 324834 533488
rect 325514 528944 325570 529000
rect 324318 524320 324374 524376
rect 324318 521056 324374 521112
rect 326986 527584 327042 527640
rect 331770 535880 331826 535936
rect 333334 534520 333390 534576
rect 336922 538736 336978 538792
rect 336462 535200 336518 535256
rect 334898 529488 334954 529544
rect 334898 528400 334954 528456
rect 338026 539144 338082 539200
rect 339590 542816 339646 542872
rect 341154 541456 341210 541512
rect 342718 548256 342774 548312
rect 344282 544040 344338 544096
rect 347410 548392 347466 548448
rect 345846 544720 345902 544776
rect 350446 551792 350502 551848
rect 353666 553560 353722 553616
rect 359922 537240 359978 537296
rect 361486 553696 361542 553752
rect 367006 523776 367062 523832
rect 367006 521192 367062 521248
rect 372250 546624 372306 546680
rect 372250 521328 372306 521384
rect 374734 614760 374790 614816
rect 374642 599120 374698 599176
rect 461674 647536 461730 647592
rect 461582 644816 461638 644872
rect 376758 642640 376814 642696
rect 375470 610408 375526 610464
rect 376022 634480 376078 634536
rect 376022 622920 376078 622976
rect 375654 618568 375710 618624
rect 375562 609592 375618 609648
rect 375470 600616 375526 600672
rect 375562 597352 375618 597408
rect 375930 614488 375986 614544
rect 375838 596536 375894 596592
rect 375746 594088 375802 594144
rect 376942 641280 376998 641336
rect 376758 607960 376814 608016
rect 377126 625096 377182 625152
rect 377678 625912 377734 625968
rect 377678 624280 377734 624336
rect 377770 623464 377826 623520
rect 377218 622648 377274 622704
rect 377034 621832 377090 621888
rect 377034 621036 377090 621072
rect 377034 621016 377036 621036
rect 377036 621016 377088 621036
rect 377088 621016 377090 621036
rect 378046 619656 378102 619712
rect 378046 616120 378102 616176
rect 377126 612040 377182 612096
rect 376942 611224 376998 611280
rect 376850 607144 376906 607200
rect 376758 601432 376814 601488
rect 376114 575320 376170 575376
rect 376022 573688 376078 573744
rect 376850 598168 376906 598224
rect 376758 530712 376814 530768
rect 377034 588376 377090 588432
rect 377034 585928 377090 585984
rect 377034 579400 377090 579456
rect 377034 576136 377090 576192
rect 378046 606328 378102 606384
rect 377954 605512 378010 605568
rect 378046 604696 378102 604752
rect 378046 603880 378102 603936
rect 378046 603100 378048 603120
rect 378048 603100 378100 603120
rect 378100 603100 378102 603120
rect 378046 603064 378102 603100
rect 378046 594904 378102 594960
rect 377954 593272 378010 593328
rect 378046 592456 378102 592512
rect 378046 590824 378102 590880
rect 378046 590008 378102 590064
rect 378046 589192 378102 589248
rect 377862 587560 377918 587616
rect 377862 586744 377918 586800
rect 377218 585112 377274 585168
rect 377770 584296 377826 584352
rect 378046 583480 378102 583536
rect 378046 582664 378102 582720
rect 378046 581052 378102 581088
rect 378046 581032 378048 581052
rect 378048 581032 378100 581052
rect 378100 581032 378102 581052
rect 378046 580216 378102 580272
rect 378046 578584 378102 578640
rect 378046 574504 378102 574560
rect 377586 572872 377642 572928
rect 377954 569608 378010 569664
rect 376850 529216 376906 529272
rect 378322 617752 378378 617808
rect 378690 613672 378746 613728
rect 378414 612856 378470 612912
rect 378598 599800 378654 599856
rect 378506 595720 378562 595776
rect 377126 524184 377182 524240
rect 375470 519696 375526 519752
rect 379610 577768 379666 577824
rect 380254 544856 380310 544912
rect 379610 534112 379666 534168
rect 378598 521328 378654 521384
rect 384302 622920 384358 622976
rect 384302 611360 384358 611416
rect 391202 611360 391258 611416
rect 382278 581848 382334 581904
rect 381818 557232 381874 557288
rect 383382 556960 383438 557016
rect 382278 518064 382334 518120
rect 383842 591640 383898 591696
rect 383842 530576 383898 530632
rect 384854 521056 384910 521112
rect 386510 556824 386566 556880
rect 388074 556688 388130 556744
rect 391202 599528 391258 599584
rect 403622 599528 403678 599584
rect 403622 582936 403678 582992
rect 427082 582936 427138 582992
rect 427082 578312 427138 578368
rect 431958 578312 432014 578368
rect 431958 572736 432014 572792
rect 408406 559680 408462 559736
rect 406842 551656 406898 551712
rect 400586 543496 400642 543552
rect 389638 539280 389694 539336
rect 397366 536696 397422 536752
rect 395894 533976 395950 534032
rect 394330 532616 394386 532672
rect 392766 524048 392822 524104
rect 391110 521192 391166 521248
rect 399022 536560 399078 536616
rect 402150 525408 402206 525464
rect 405278 522688 405334 522744
rect 420826 559544 420882 559600
rect 416226 547304 416282 547360
rect 414662 546216 414718 546272
rect 413098 542136 413154 542192
rect 409970 540912 410026 540968
rect 411534 528264 411590 528320
rect 417790 544448 417846 544504
rect 419354 537648 419410 537704
rect 435362 572736 435418 572792
rect 435362 560224 435418 560280
rect 437662 560224 437718 560280
rect 453762 555600 453818 555656
rect 437662 553288 437718 553344
rect 434994 550024 435050 550080
rect 430302 548528 430358 548584
rect 428738 541592 428794 541648
rect 425610 528128 425666 528184
rect 427174 533568 427230 533624
rect 438122 537512 438178 537568
rect 452198 545672 452254 545728
rect 444286 542952 444342 543008
rect 442814 540232 442870 540288
rect 441250 527992 441306 528048
rect 445942 537376 445998 537432
rect 449070 531120 449126 531176
rect 460018 528672 460074 528728
rect 458454 527720 458510 527776
rect 461674 521056 461730 521112
rect 461858 644952 461914 645008
rect 473266 655968 473322 656024
rect 467286 647400 467342 647456
rect 467102 647264 467158 647320
rect 464342 646720 464398 646776
rect 462962 639512 463018 639568
rect 462318 599528 462374 599584
rect 462226 553288 462282 553344
rect 462226 550024 462282 550080
rect 461858 521192 461914 521248
rect 462962 519696 463018 519752
rect 461582 518336 461638 518392
rect 464342 522552 464398 522608
rect 464618 636520 464674 636576
rect 464526 634888 464582 634944
rect 464618 522688 464674 522744
rect 464526 521328 464582 521384
rect 467746 555464 467802 555520
rect 472622 643592 472678 643648
rect 471518 637744 471574 637800
rect 471426 635024 471482 635080
rect 471610 550024 471666 550080
rect 471610 524320 471666 524376
rect 471886 522960 471942 523016
rect 471518 522008 471574 522064
rect 476026 655832 476082 655888
rect 475934 654608 475990 654664
rect 473358 524320 473414 524376
rect 473266 521600 473322 521656
rect 472622 521464 472678 521520
rect 473358 520784 473414 520840
rect 477406 655696 477462 655752
rect 476118 518336 476174 518392
rect 476946 547032 477002 547088
rect 486974 657736 487030 657792
rect 508502 700304 508558 700360
rect 484030 657328 484086 657384
rect 479246 639240 479302 639296
rect 478510 599664 478566 599720
rect 477406 518744 477462 518800
rect 478786 518744 478842 518800
rect 476946 518200 477002 518256
rect 478510 518200 478566 518256
rect 477314 518064 477370 518120
rect 478786 518084 478842 518120
rect 478786 518064 478788 518084
rect 478788 518064 478840 518084
rect 478840 518064 478842 518084
rect 478510 517792 478566 517848
rect 479338 467336 479394 467392
rect 479982 637608 480038 637664
rect 479890 539008 479946 539064
rect 479522 476040 479578 476096
rect 479430 453192 479486 453248
rect 479522 449928 479578 449984
rect 60738 389000 60794 389056
rect 60646 387640 60702 387696
rect 60462 387368 60518 387424
rect 62118 387368 62174 387424
rect 62578 386960 62634 387016
rect 60922 386824 60978 386880
rect 60738 383696 60794 383752
rect 59266 298696 59322 298752
rect 50986 262928 51042 262984
rect 47582 261160 47638 261216
rect 40682 261024 40738 261080
rect 35162 260888 35218 260944
rect 15842 193840 15898 193896
rect 14738 127608 14794 127664
rect 11702 126248 11758 126304
rect 8758 98640 8814 98696
rect 4894 32816 4950 32872
rect 4802 32408 4858 32464
rect 4066 26968 4122 27024
rect 7654 4800 7710 4856
rect 4894 3440 4950 3496
rect 6458 3440 6514 3496
rect 5262 3304 5318 3360
rect 13542 100000 13598 100056
rect 12346 6160 12402 6216
rect 9954 3440 10010 3496
rect 11702 3440 11758 3496
rect 31298 181328 31354 181384
rect 23018 144064 23074 144120
rect 17038 137672 17094 137728
rect 15842 3712 15898 3768
rect 21822 137536 21878 137592
rect 18234 122168 18290 122224
rect 19430 116456 19486 116512
rect 26514 137808 26570 137864
rect 24214 115096 24270 115152
rect 30102 137128 30158 137184
rect 28906 134408 28962 134464
rect 27710 3440 27766 3496
rect 33598 136992 33654 137048
rect 32402 101360 32458 101416
rect 34794 109656 34850 109712
rect 40682 162832 40738 162888
rect 44178 137672 44234 137728
rect 44270 137264 44326 137320
rect 37186 136856 37242 136912
rect 35990 120672 36046 120728
rect 35254 112376 35310 112432
rect 35162 71576 35218 71632
rect 35254 3440 35310 3496
rect 40682 136720 40738 136776
rect 38382 113736 38438 113792
rect 39578 104080 39634 104136
rect 43074 122032 43130 122088
rect 41878 111016 41934 111072
rect 45466 124888 45522 124944
rect 52918 262792 52974 262848
rect 63498 383560 63554 383616
rect 63498 375400 63554 375456
rect 65062 375400 65118 375456
rect 65062 369688 65118 369744
rect 67546 385600 67602 385656
rect 65890 373224 65946 373280
rect 65430 338680 65486 338736
rect 64510 265512 64566 265568
rect 65522 262928 65578 262984
rect 70306 369688 70362 369744
rect 70398 366288 70454 366344
rect 77942 366288 77998 366344
rect 69018 346976 69074 347032
rect 69662 262792 69718 262848
rect 77942 347656 77998 347712
rect 78862 347656 78918 347712
rect 78862 344664 78918 344720
rect 72514 272584 72570 272640
rect 94134 390088 94190 390144
rect 90546 388728 90602 388784
rect 90546 386960 90602 387016
rect 86958 386824 87014 386880
rect 83462 363568 83518 363624
rect 79138 301416 79194 301472
rect 83462 298696 83518 298752
rect 86866 344664 86922 344720
rect 86866 341944 86922 342000
rect 90362 341944 90418 342000
rect 90362 332560 90418 332616
rect 91742 332560 91798 332616
rect 91742 323584 91798 323640
rect 97262 389000 97318 389056
rect 95698 386552 95754 386608
rect 94134 265512 94190 265568
rect 101310 388864 101366 388920
rect 106186 387096 106242 387152
rect 105634 386688 105690 386744
rect 101310 385600 101366 385656
rect 97262 373224 97318 373280
rect 97354 371864 97410 371920
rect 95882 323584 95938 323640
rect 95882 311888 95938 311944
rect 99010 319232 99066 319288
rect 99378 311888 99434 311944
rect 99378 307672 99434 307728
rect 102046 307672 102102 307728
rect 102046 304544 102102 304600
rect 104806 304544 104862 304600
rect 104806 300600 104862 300656
rect 100574 267144 100630 267200
rect 108394 386960 108450 387016
rect 108302 386552 108358 386608
rect 115294 387096 115350 387152
rect 112074 386280 112130 386336
rect 112442 386280 112498 386336
rect 109682 300600 109738 300656
rect 109682 295296 109738 295352
rect 115846 386824 115902 386880
rect 119342 387232 119398 387288
rect 118698 386688 118754 386744
rect 122838 387640 122894 387696
rect 113822 295296 113878 295352
rect 112442 272584 112498 272640
rect 102138 263472 102194 263528
rect 105542 263472 105598 263528
rect 108946 263200 109002 263256
rect 105910 263064 105966 263120
rect 104806 262792 104862 262848
rect 107566 262928 107622 262984
rect 105910 261160 105966 261216
rect 103794 261024 103850 261080
rect 104806 261024 104862 261080
rect 108946 262248 109002 262304
rect 107566 260888 107622 260944
rect 125598 387504 125654 387560
rect 126426 387504 126482 387560
rect 124126 386824 124182 386880
rect 129738 387368 129794 387424
rect 134522 386688 134578 386744
rect 132590 386416 132646 386472
rect 133602 386416 133658 386472
rect 125598 301416 125654 301472
rect 135902 386552 135958 386608
rect 137282 386416 137338 386472
rect 135902 263064 135958 263120
rect 150438 387368 150494 387424
rect 158718 387368 158774 387424
rect 150438 386824 150494 386880
rect 151542 386824 151598 386880
rect 166262 388592 166318 388648
rect 179418 386688 179474 386744
rect 180246 386688 180302 386744
rect 173162 384920 173218 384976
rect 169022 383560 169078 383616
rect 166262 371864 166318 371920
rect 169022 319368 169078 319424
rect 183834 386552 183890 386608
rect 184846 386552 184902 386608
rect 186962 386416 187018 386472
rect 184846 386144 184902 386200
rect 179418 384784 179474 384840
rect 186962 383424 187018 383480
rect 173162 267008 173218 267064
rect 138662 263200 138718 263256
rect 137282 262928 137338 262984
rect 134522 262792 134578 262848
rect 117962 257896 118018 257952
rect 116398 252456 116454 252512
rect 113822 245656 113878 245712
rect 114650 245656 114706 245712
rect 114650 240080 114706 240136
rect 48226 215056 48282 215112
rect 50986 198464 51042 198520
rect 57886 198192 57942 198248
rect 56230 197784 56286 197840
rect 54574 197648 54630 197704
rect 52918 197376 52974 197432
rect 64510 198328 64566 198384
rect 59266 140256 59322 140312
rect 62578 138896 62634 138952
rect 60922 138760 60978 138816
rect 70398 198464 70454 198520
rect 69478 197920 69534 197976
rect 72790 198056 72846 198112
rect 71778 197784 71834 197840
rect 71134 197512 71190 197568
rect 75918 199960 75974 200016
rect 77758 198600 77814 198656
rect 79322 198192 79378 198248
rect 73158 197648 73214 197704
rect 74446 197648 74502 197704
rect 82726 199688 82782 199744
rect 84106 199280 84162 199336
rect 81070 198872 81126 198928
rect 85578 198328 85634 198384
rect 86038 198192 86094 198248
rect 87694 198464 87750 198520
rect 92386 199416 92442 199472
rect 94502 199960 94558 200016
rect 95974 199960 96030 200016
rect 95238 199280 95294 199336
rect 94318 199008 94374 199064
rect 91006 198736 91062 198792
rect 89350 198328 89406 198384
rect 88338 197920 88394 197976
rect 96618 197648 96674 197704
rect 97998 198056 98054 198112
rect 100620 199824 100676 199880
rect 100666 199724 100668 199744
rect 100668 199724 100720 199744
rect 100720 199724 100722 199744
rect 100666 199688 100722 199724
rect 102598 199688 102654 199744
rect 103426 198872 103482 198928
rect 99194 197920 99250 197976
rect 86958 197512 87014 197568
rect 97630 197512 97686 197568
rect 105910 199552 105966 199608
rect 104898 199416 104954 199472
rect 107658 199960 107714 200016
rect 107566 199416 107622 199472
rect 108946 199280 109002 199336
rect 106278 198736 106334 198792
rect 104254 197784 104310 197840
rect 78586 197376 78642 197432
rect 79414 197376 79470 197432
rect 104162 197376 104218 197432
rect 67546 197240 67602 197296
rect 95146 195200 95202 195256
rect 65890 137944 65946 138000
rect 66166 137536 66222 137592
rect 89166 130328 89222 130384
rect 85670 128968 85726 129024
rect 47582 110608 47638 110664
rect 46662 97144 46718 97200
rect 52918 87760 52974 87816
rect 50986 85720 51042 85776
rect 60646 87624 60702 87680
rect 57610 87352 57666 87408
rect 54666 87080 54722 87136
rect 56506 86128 56562 86184
rect 59266 87216 59322 87272
rect 62026 87488 62082 87544
rect 63866 85584 63922 85640
rect 65614 87896 65670 87952
rect 84842 87624 84898 87680
rect 68650 85856 68706 85912
rect 80748 84904 80804 84960
rect 77620 84768 77676 84824
rect 71364 84632 71420 84688
rect 79184 84496 79240 84552
rect 48226 81640 48282 81696
rect 47858 80280 47914 80336
rect 47490 63960 47546 64016
rect 47582 61240 47638 61296
rect 47766 58520 47822 58576
rect 47674 57160 47730 57216
rect 47674 28192 47730 28248
rect 48134 65320 48190 65376
rect 48042 62600 48098 62656
rect 47950 59880 48006 59936
rect 47858 46280 47914 46336
rect 47766 26832 47822 26888
rect 47950 25472 48006 25528
rect 85026 87352 85082 87408
rect 85026 80688 85082 80744
rect 84842 79328 84898 79384
rect 49422 78920 49478 78976
rect 49330 77560 49386 77616
rect 49238 69400 49294 69456
rect 49146 68040 49202 68096
rect 49054 55800 49110 55856
rect 48226 49000 48282 49056
rect 48134 43560 48190 43616
rect 48962 28464 49018 28520
rect 48042 22616 48098 22672
rect 47582 21256 47638 21312
rect 47490 15816 47546 15872
rect 47858 6296 47914 6352
rect 49146 39208 49202 39264
rect 49330 48864 49386 48920
rect 50434 75928 50490 75984
rect 49606 74840 49662 74896
rect 49514 72120 49570 72176
rect 49422 44784 49478 44840
rect 49238 37848 49294 37904
rect 49514 36488 49570 36544
rect 50158 70352 50214 70408
rect 50066 52536 50122 52592
rect 50066 42200 50122 42256
rect 49606 33768 49662 33824
rect 49054 24112 49110 24168
rect 50250 66272 50306 66328
rect 50158 18536 50214 18592
rect 50342 49136 50398 49192
rect 50250 17176 50306 17232
rect 50526 73208 50582 73264
rect 50618 53896 50674 53952
rect 50526 35128 50582 35184
rect 50434 30912 50490 30968
rect 84658 53216 84714 53272
rect 67914 50224 67970 50280
rect 50986 47776 51042 47832
rect 52366 47640 52422 47696
rect 53746 47504 53802 47560
rect 51354 38120 51410 38176
rect 50618 29552 50674 29608
rect 52550 29824 52606 29880
rect 54942 21528 54998 21584
rect 53746 2760 53802 2816
rect 56506 46144 56562 46200
rect 56046 31184 56102 31240
rect 55034 9016 55090 9072
rect 57242 14728 57298 14784
rect 58438 25608 58494 25664
rect 57794 8880 57850 8936
rect 60646 47912 60702 47968
rect 60830 44920 60886 44976
rect 59634 32680 59690 32736
rect 59174 10240 59230 10296
rect 62762 47912 62818 47968
rect 62026 22752 62082 22808
rect 61934 12960 61990 13016
rect 64786 46960 64842 47016
rect 65614 46960 65670 47016
rect 63314 43424 63370 43480
rect 65522 36624 65578 36680
rect 63222 28328 63278 28384
rect 62762 11600 62818 11656
rect 64326 3440 64382 3496
rect 66074 42064 66130 42120
rect 65614 19896 65670 19952
rect 67454 14456 67510 14512
rect 66718 10376 66774 10432
rect 68834 40568 68890 40624
rect 69110 33904 69166 33960
rect 71502 49272 71558 49328
rect 70214 32408 70270 32464
rect 70306 31048 70362 31104
rect 77206 48048 77262 48104
rect 79322 48048 79378 48104
rect 78586 47912 78642 47968
rect 74446 46960 74502 47016
rect 75182 46960 75238 47016
rect 74998 37984 75054 38040
rect 72974 13096 73030 13152
rect 72422 11736 72478 11792
rect 73802 7792 73858 7848
rect 72606 6432 72662 6488
rect 75182 20032 75238 20088
rect 78586 21392 78642 21448
rect 76562 14592 76618 14648
rect 76194 6568 76250 6624
rect 77390 5072 77446 5128
rect 79506 47912 79562 47968
rect 79506 24248 79562 24304
rect 84106 47912 84162 47968
rect 81254 40704 81310 40760
rect 83002 39344 83058 39400
rect 83278 35264 83334 35320
rect 82082 32544 82138 32600
rect 80886 29688 80942 29744
rect 80702 17312 80758 17368
rect 79322 15952 79378 16008
rect 79690 6704 79746 6760
rect 86866 93064 86922 93120
rect 86222 87760 86278 87816
rect 86222 51856 86278 51912
rect 87694 90480 87750 90536
rect 87602 87080 87658 87136
rect 87050 52536 87106 52592
rect 86958 51720 87014 51776
rect 87050 32816 87106 32872
rect 87786 87488 87842 87544
rect 87786 54576 87842 54632
rect 87694 52536 87750 52592
rect 88246 51740 88302 51776
rect 88246 51720 88248 51740
rect 88248 51720 88300 51740
rect 88300 51720 88302 51740
rect 87694 47912 87750 47968
rect 87694 18672 87750 18728
rect 87970 9152 88026 9208
rect 87602 4936 87658 4992
rect 92754 124752 92810 124808
rect 91558 123528 91614 123584
rect 90362 108296 90418 108352
rect 91742 87896 91798 87952
rect 91926 87216 91982 87272
rect 91926 53080 91982 53136
rect 91742 7520 91798 7576
rect 93950 117952 94006 118008
rect 105726 141344 105782 141400
rect 101402 133184 101458 133240
rect 98642 120808 98698 120864
rect 96250 119312 96306 119368
rect 97446 106800 97502 106856
rect 99838 102720 99894 102776
rect 101034 94424 101090 94480
rect 103334 131688 103390 131744
rect 102230 101496 102286 101552
rect 101402 3440 101458 3496
rect 104530 105440 104586 105496
rect 105542 80280 105598 80336
rect 105542 51720 105598 51776
rect 106922 98776 106978 98832
rect 108118 95784 108174 95840
rect 112810 192480 112866 192536
rect 110510 108432 110566 108488
rect 109314 3440 109370 3496
rect 111614 97280 111670 97336
rect 115846 137828 115902 137864
rect 115846 137808 115848 137828
rect 115848 137808 115900 137828
rect 115900 137808 115902 137828
rect 115202 137400 115258 137456
rect 114006 123392 114062 123448
rect 116582 240080 116638 240136
rect 116582 224168 116638 224224
rect 178682 256808 178738 256864
rect 123482 254632 123538 254688
rect 120722 224168 120778 224224
rect 121458 211112 121514 211168
rect 118790 137536 118846 137592
rect 118698 137128 118754 137184
rect 117962 3304 118018 3360
rect 117594 2896 117650 2952
rect 122286 104216 122342 104272
rect 119894 102856 119950 102912
rect 121090 90344 121146 90400
rect 163502 250280 163558 250336
rect 126242 243752 126298 243808
rect 123574 211112 123630 211168
rect 123574 200640 123630 200696
rect 124678 100136 124734 100192
rect 142802 240488 142858 240544
rect 140042 237224 140098 237280
rect 138662 231784 138718 231840
rect 126978 134544 127034 134600
rect 126242 9152 126298 9208
rect 130566 127744 130622 127800
rect 134154 119448 134210 119504
rect 137650 118088 137706 118144
rect 138662 28464 138718 28520
rect 141238 130464 141294 130520
rect 140042 10376 140098 10432
rect 151082 239400 151138 239456
rect 146942 233960 146998 234016
rect 144182 228520 144238 228576
rect 144734 138216 144790 138272
rect 144182 113736 144238 113792
rect 142802 5072 142858 5128
rect 148322 116592 148378 116648
rect 146942 31184 146998 31240
rect 152462 229608 152518 229664
rect 151818 129104 151874 129160
rect 151082 7792 151138 7848
rect 155222 227432 155278 227488
rect 152462 111016 152518 111072
rect 158718 218728 158774 218784
rect 162490 136040 162546 136096
rect 155406 111016 155462 111072
rect 155222 109656 155278 109712
rect 158902 109656 158958 109712
rect 174542 232872 174598 232928
rect 166078 136176 166134 136232
rect 163502 3440 163558 3496
rect 176658 138352 176714 138408
rect 174542 29824 174598 29880
rect 173162 3440 173218 3496
rect 169574 3304 169630 3360
rect 214654 382880 214710 382936
rect 212538 265512 212594 265568
rect 208950 264424 209006 264480
rect 205362 263336 205418 263392
rect 201774 262112 201830 262168
rect 198186 261160 198242 261216
rect 194598 260208 194654 260264
rect 198002 253544 198058 253600
rect 188342 242664 188398 242720
rect 187330 139032 187386 139088
rect 183742 138624 183798 138680
rect 178682 26968 178738 27024
rect 180246 3576 180302 3632
rect 191102 230696 191158 230752
rect 190826 129240 190882 129296
rect 188342 53216 188398 53272
rect 195242 220768 195298 220824
rect 194414 134680 194470 134736
rect 191102 124888 191158 124944
rect 197910 131824 197966 131880
rect 195242 98640 195298 98696
rect 202142 249192 202198 249248
rect 199382 235048 199438 235104
rect 198002 102856 198058 102912
rect 209042 248104 209098 248160
rect 206282 224168 206338 224224
rect 203522 221992 203578 222048
rect 202142 141344 202198 141400
rect 201498 139984 201554 140040
rect 199382 32680 199438 32736
rect 206282 144064 206338 144120
rect 206282 139304 206338 139360
rect 205638 138216 205694 138272
rect 203522 100000 203578 100056
rect 208582 131960 208638 132016
rect 205086 3712 205142 3768
rect 206282 3712 206338 3768
rect 211802 244840 211858 244896
rect 210422 241440 210478 241496
rect 209042 101496 209098 101552
rect 214562 238312 214618 238368
rect 213182 219816 213238 219872
rect 212170 126384 212226 126440
rect 211802 123528 211858 123584
rect 210422 29688 210478 29744
rect 213182 90480 213238 90536
rect 219714 267688 219770 267744
rect 216126 266600 216182 266656
rect 216034 245928 216090 245984
rect 215942 223080 215998 223136
rect 214654 205536 214710 205592
rect 215666 138488 215722 138544
rect 215298 138352 215354 138408
rect 214562 31048 214618 31104
rect 219438 200640 219494 200696
rect 222934 342352 222990 342408
rect 222842 258984 222898 259040
rect 219438 199144 219494 199200
rect 216034 195200 216090 195256
rect 218058 138624 218114 138680
rect 219254 138624 219310 138680
rect 215942 122168 215998 122224
rect 222750 124888 222806 124944
rect 223210 340856 223266 340912
rect 226338 342352 226394 342408
rect 226614 342216 226670 342272
rect 225050 341808 225106 341864
rect 224958 341536 225014 341592
rect 225142 341672 225198 341728
rect 225786 341400 225842 341456
rect 225602 340040 225658 340096
rect 225418 339768 225474 339824
rect 223302 268776 223358 268832
rect 223302 226208 223358 226264
rect 223210 198600 223266 198656
rect 222934 198192 222990 198248
rect 225418 199552 225474 199608
rect 225970 341128 226026 341184
rect 226154 340720 226210 340776
rect 225970 199416 226026 199472
rect 228914 380704 228970 380760
rect 228730 380296 228786 380352
rect 228638 377304 228694 377360
rect 227626 342216 227682 342272
rect 227534 338408 227590 338464
rect 226890 269864 226946 269920
rect 227718 342080 227774 342136
rect 228362 340992 228418 341048
rect 227810 340856 227866 340912
rect 228178 340856 228234 340912
rect 227626 257760 227682 257816
rect 227534 256672 227590 256728
rect 226982 246880 227038 246936
rect 226154 199280 226210 199336
rect 226338 199144 226394 199200
rect 226338 198056 226394 198112
rect 225786 197784 225842 197840
rect 225602 197240 225658 197296
rect 223302 181328 223358 181384
rect 226338 123528 226394 123584
rect 222842 91704 222898 91760
rect 228270 339632 228326 339688
rect 228270 199824 228326 199880
rect 228178 199688 228234 199744
rect 228546 340312 228602 340368
rect 228362 197920 228418 197976
rect 228638 327528 228694 327584
rect 228822 380160 228878 380216
rect 228822 322088 228878 322144
rect 228730 317736 228786 317792
rect 230386 380568 230442 380624
rect 230202 378664 230258 378720
rect 229006 374584 229062 374640
rect 228730 316648 228786 316704
rect 228914 316648 228970 316704
rect 230294 377440 230350 377496
rect 230202 328616 230258 328672
rect 230294 323176 230350 323232
rect 230386 318688 230442 318744
rect 229006 309032 229062 309088
rect 231766 387776 231822 387832
rect 231582 382880 231638 382936
rect 231490 376760 231546 376816
rect 231030 338816 231086 338872
rect 230938 338544 230994 338600
rect 230478 270952 230534 271008
rect 228914 251368 228970 251424
rect 228730 202408 228786 202464
rect 228546 197512 228602 197568
rect 231122 236136 231178 236192
rect 230938 199008 230994 199064
rect 228914 192480 228970 192536
rect 226982 120808 227038 120864
rect 231214 198464 231270 198520
rect 231490 329568 231546 329624
rect 231674 380432 231730 380488
rect 231674 319912 231730 319968
rect 231582 313384 231638 313440
rect 231398 198328 231454 198384
rect 233146 383288 233202 383344
rect 233054 383016 233110 383072
rect 232962 380840 233018 380896
rect 232870 377712 232926 377768
rect 232870 324264 232926 324320
rect 232962 314472 233018 314528
rect 233054 311208 233110 311264
rect 232594 222672 232650 222728
rect 232502 221040 232558 221096
rect 231766 193704 231822 193760
rect 232686 219408 232742 219464
rect 232778 216144 232834 216200
rect 232594 141888 232650 141944
rect 232962 214512 233018 214568
rect 233698 377576 233754 377632
rect 233882 364928 233938 364984
rect 233790 351328 233846 351384
rect 233698 325352 233754 325408
rect 233974 352552 234030 352608
rect 233882 307944 233938 308000
rect 233790 297064 233846 297120
rect 233974 295976 234030 296032
rect 234526 388456 234582 388512
rect 234434 380024 234490 380080
rect 234250 362480 234306 362536
rect 234158 356904 234214 356960
rect 234158 294888 234214 294944
rect 234342 360984 234398 361040
rect 234250 290536 234306 290592
rect 234434 306856 234490 306912
rect 234342 287272 234398 287328
rect 234066 274488 234122 274544
rect 233146 194792 233202 194848
rect 232962 140120 233018 140176
rect 232778 139712 232834 139768
rect 233146 139032 233202 139088
rect 232502 138216 232558 138272
rect 235538 388320 235594 388376
rect 235078 377848 235134 377904
rect 235446 374720 235502 374776
rect 235354 359352 235410 359408
rect 235262 354048 235318 354104
rect 235170 349968 235226 350024
rect 235078 326440 235134 326496
rect 235170 304680 235226 304736
rect 235354 305768 235410 305824
rect 235262 303456 235318 303512
rect 235446 301416 235502 301472
rect 239218 387368 239274 387424
rect 236458 386824 236514 386880
rect 237654 386824 237710 386880
rect 239034 386824 239090 386880
rect 235814 356632 235870 356688
rect 235630 343712 235686 343768
rect 235538 300328 235594 300384
rect 235538 207032 235594 207088
rect 234894 206352 234950 206408
rect 234526 195880 234582 195936
rect 235262 201456 235318 201512
rect 235630 204856 235686 204912
rect 235538 192616 235594 192672
rect 235906 348472 235962 348528
rect 235814 187176 235870 187232
rect 235722 184864 235778 184920
rect 238574 375944 238630 376000
rect 236826 369144 236882 369200
rect 236734 362208 236790 362264
rect 236550 345616 236606 345672
rect 236458 329704 236514 329760
rect 236550 310120 236606 310176
rect 237930 369008 237986 369064
rect 237286 355272 237342 355328
rect 237194 353912 237250 353968
rect 237010 351056 237066 351112
rect 236826 321000 236882 321056
rect 236734 315560 236790 315616
rect 236918 312296 236974 312352
rect 236642 299240 236698 299296
rect 237010 289720 237066 289776
rect 237102 191528 237158 191584
rect 237194 190304 237250 190360
rect 237378 341436 237380 341456
rect 237380 341436 237432 341456
rect 237432 341436 237434 341456
rect 237378 341400 237434 341436
rect 237746 341400 237802 341456
rect 237470 340992 237526 341048
rect 237470 340312 237526 340368
rect 237378 340040 237434 340096
rect 237562 339632 237618 339688
rect 237654 333240 237710 333296
rect 237838 340040 237894 340096
rect 238482 351192 238538 351248
rect 238022 345888 238078 345944
rect 238206 341536 238262 341592
rect 238206 340312 238262 340368
rect 238114 340176 238170 340232
rect 237930 331880 237986 331936
rect 237930 331064 237986 331120
rect 237838 291624 237894 291680
rect 237746 285096 237802 285152
rect 238022 329704 238078 329760
rect 237930 279656 237986 279712
rect 237654 275304 237710 275360
rect 237378 274488 237434 274544
rect 238114 289448 238170 289504
rect 238390 337456 238446 337512
rect 238298 292712 238354 292768
rect 238206 288360 238262 288416
rect 238666 339360 238722 339416
rect 238574 332968 238630 333024
rect 238482 330792 238538 330848
rect 238390 286184 238446 286240
rect 239126 341672 239182 341728
rect 239034 333240 239090 333296
rect 239586 346024 239642 346080
rect 239494 344256 239550 344312
rect 239402 342896 239458 342952
rect 239310 340584 239366 340640
rect 239218 331064 239274 331120
rect 239402 282784 239458 282840
rect 240046 342216 240102 342272
rect 240046 340856 240102 340912
rect 239954 340720 240010 340776
rect 239678 340448 239734 340504
rect 239586 284008 239642 284064
rect 239494 281832 239550 281888
rect 239310 280744 239366 280800
rect 240046 339924 240102 339960
rect 240046 339904 240048 339924
rect 240048 339904 240100 339924
rect 240100 339904 240102 339924
rect 239862 339768 239918 339824
rect 240046 339768 240102 339824
rect 244830 386824 244886 386880
rect 249890 387640 249946 387696
rect 241794 363704 241850 363760
rect 246302 357992 246358 358048
rect 242714 344936 242770 344992
rect 242806 343712 242862 343768
rect 245842 343168 245898 343224
rect 245658 343032 245714 343088
rect 244830 342760 244886 342816
rect 243542 342624 243598 342680
rect 244278 342488 244334 342544
rect 243818 342216 243874 342272
rect 247038 343576 247094 343632
rect 247866 343032 247922 343088
rect 246854 342488 246910 342544
rect 246302 342216 246358 342272
rect 248878 342624 248934 342680
rect 248510 340448 248566 340504
rect 249706 342352 249762 342408
rect 251914 387504 251970 387560
rect 251086 343440 251142 343496
rect 250902 343304 250958 343360
rect 254950 369280 255006 369336
rect 253938 367648 253994 367704
rect 252926 344800 252982 344856
rect 252190 339904 252246 339960
rect 253202 344528 253258 344584
rect 255318 344120 255374 344176
rect 259182 387368 259238 387424
rect 256054 386824 256110 386880
rect 255962 344664 256018 344720
rect 255594 341672 255650 341728
rect 258722 386688 258778 386744
rect 257986 381656 258042 381712
rect 256974 344528 257030 344584
rect 256698 344392 256754 344448
rect 256054 343032 256110 343088
rect 260010 377168 260066 377224
rect 258998 371864 259054 371920
rect 258722 343168 258778 343224
rect 260746 376760 260802 376816
rect 261022 373360 261078 373416
rect 262034 342216 262090 342272
rect 264242 370640 264298 370696
rect 262862 359488 262918 359544
rect 264058 344392 264114 344448
rect 263598 344004 263654 344040
rect 263598 343984 263600 344004
rect 263600 343984 263652 344004
rect 263652 343984 263654 344004
rect 262862 342216 262918 342272
rect 263046 342216 263102 342272
rect 262770 340584 262826 340640
rect 265070 366288 265126 366344
rect 264242 342216 264298 342272
rect 267094 365064 267150 365120
rect 267002 360848 267058 360904
rect 266358 344256 266414 344312
rect 268106 344256 268162 344312
rect 270130 387368 270186 387424
rect 269946 342896 270002 342952
rect 269118 342216 269174 342272
rect 270406 387232 270462 387288
rect 273166 387232 273222 387288
rect 272522 386960 272578 387016
rect 271234 378800 271290 378856
rect 271142 376216 271198 376272
rect 271234 342216 271290 342272
rect 272154 342216 272210 342272
rect 274638 387096 274694 387152
rect 275190 386960 275246 387016
rect 273902 362344 273958 362400
rect 273534 346024 273590 346080
rect 274178 356768 274234 356824
rect 273902 342216 273958 342272
rect 276202 343168 276258 343224
rect 277122 341400 277178 341456
rect 278226 343032 278282 343088
rect 279238 342896 279294 342952
rect 241242 339360 241298 339416
rect 280158 338408 280214 338464
rect 239862 278500 239918 278556
rect 239862 277412 239918 277468
rect 239678 276324 239734 276380
rect 238666 274216 238722 274272
rect 238022 273128 238078 273184
rect 237378 272040 237434 272096
rect 238206 260072 238262 260128
rect 238114 255584 238170 255640
rect 238022 225120 238078 225176
rect 237378 214240 237434 214296
rect 237378 201320 237434 201376
rect 237378 199144 237434 199200
rect 237286 146920 237342 146976
rect 280342 295160 280398 295216
rect 280526 338544 280582 338600
rect 280434 293800 280490 293856
rect 282182 384376 282238 384432
rect 280710 341536 280766 341592
rect 280894 341128 280950 341184
rect 280710 297744 280766 297800
rect 280618 296384 280674 296440
rect 280894 299376 280950 299432
rect 280986 298016 281042 298072
rect 280802 295976 280858 296032
rect 280526 292440 280582 292496
rect 282274 383152 282330 383208
rect 282826 379480 282882 379536
rect 282826 376760 282882 376816
rect 282918 376080 282974 376136
rect 282366 338816 282422 338872
rect 282274 323584 282330 323640
rect 282182 319504 282238 319560
rect 282458 331744 282514 331800
rect 282366 317056 282422 317112
rect 282550 330384 282606 330440
rect 282458 315424 282514 315480
rect 282550 313792 282606 313848
rect 282182 299412 282184 299432
rect 282184 299412 282236 299432
rect 282236 299412 282238 299432
rect 282182 299376 282238 299412
rect 281722 293528 281778 293584
rect 281630 291080 281686 291136
rect 282182 289756 282184 289776
rect 282184 289756 282236 289776
rect 282236 289756 282238 289776
rect 282182 289720 282238 289756
rect 281538 289448 281594 289504
rect 282090 288224 282146 288280
rect 282734 287952 282790 288008
rect 282642 286592 282698 286648
rect 281538 285504 281594 285560
rect 282642 285540 282644 285560
rect 282644 285540 282696 285560
rect 282696 285540 282698 285560
rect 282642 285504 282698 285540
rect 282090 284144 282146 284200
rect 281998 281460 282000 281480
rect 282000 281460 282052 281480
rect 282052 281460 282054 281480
rect 281998 281424 282054 281460
rect 281998 279656 282054 279712
rect 282826 277752 282882 277808
rect 282734 277344 282790 277400
rect 282826 276256 282882 276312
rect 282826 275168 282882 275224
rect 282734 273672 282790 273728
rect 282826 273300 282828 273320
rect 282828 273300 282880 273320
rect 282880 273300 282882 273320
rect 282826 273264 282882 273300
rect 282826 272176 282882 272232
rect 282734 271088 282790 271144
rect 282826 270680 282882 270736
rect 281906 270000 281962 270056
rect 281906 267552 281962 267608
rect 281814 265920 281870 265976
rect 280250 263472 280306 263528
rect 282826 261976 282882 262032
rect 282550 260788 282552 260808
rect 282552 260788 282604 260808
rect 282604 260788 282606 260808
rect 282550 260752 282606 260788
rect 282550 257352 282606 257408
rect 282826 256400 282882 256456
rect 280158 255992 280214 256048
rect 282826 253408 282882 253464
rect 282826 242956 282882 242992
rect 282826 242936 282828 242956
rect 282828 242936 282880 242956
rect 282880 242936 282882 242956
rect 281538 239264 281594 239320
rect 280158 237360 280214 237416
rect 238666 216688 238722 216744
rect 238390 204856 238446 204912
rect 238206 200232 238262 200288
rect 238114 193840 238170 193896
rect 235906 143656 235962 143712
rect 235906 140664 235962 140720
rect 235262 139848 235318 139904
rect 235722 139304 235778 139360
rect 235630 138760 235686 138816
rect 237746 140664 237802 140720
rect 236826 139168 236882 139224
rect 235906 138896 235962 138952
rect 235906 138660 235908 138680
rect 235908 138660 235960 138680
rect 235960 138660 235962 138680
rect 235906 138624 235962 138660
rect 235814 138488 235870 138544
rect 235078 138216 235134 138272
rect 233882 138080 233938 138136
rect 238666 203496 238722 203552
rect 280066 201456 280122 201512
rect 238390 196968 238446 197024
rect 238574 183776 238630 183832
rect 238206 145696 238262 145752
rect 238390 141752 238446 141808
rect 239770 178404 239826 178460
rect 238574 141616 238630 141672
rect 238482 140684 238538 140720
rect 238482 140664 238484 140684
rect 238484 140664 238536 140684
rect 238536 140664 238538 140684
rect 239586 141344 239642 141400
rect 239678 140664 239734 140720
rect 238758 138216 238814 138272
rect 239862 177316 239918 177372
rect 233146 136992 233202 137048
rect 237378 136856 237434 136912
rect 233422 133320 233478 133376
rect 231122 28328 231178 28384
rect 229834 3712 229890 3768
rect 239678 135904 239734 135960
rect 238022 112376 238078 112432
rect 266910 140528 266966 140584
rect 275282 140528 275338 140584
rect 240782 139576 240838 139632
rect 239862 33088 239918 33144
rect 247590 137128 247646 137184
rect 247038 136720 247094 136776
rect 244094 136312 244150 136368
rect 242622 6160 242678 6216
rect 241426 4800 241482 4856
rect 237010 3848 237066 3904
rect 240506 3168 240562 3224
rect 241426 2760 241482 2816
rect 246302 134816 246358 134872
rect 246302 3168 246358 3224
rect 252190 137264 252246 137320
rect 254674 137264 254730 137320
rect 254582 38120 254638 38176
rect 253386 6296 253442 6352
rect 256974 25608 257030 25664
rect 258722 69400 258778 69456
rect 258170 22752 258226 22808
rect 255778 21528 255834 21584
rect 260102 54440 260158 54496
rect 259366 36624 259422 36680
rect 258722 6160 258778 6216
rect 262126 137964 262182 138000
rect 260562 33904 260618 33960
rect 262126 137944 262128 137964
rect 262128 137944 262180 137964
rect 262180 137944 262182 137964
rect 262310 137944 262366 138000
rect 261666 6432 261722 6488
rect 260102 4800 260158 4856
rect 258262 3168 258318 3224
rect 267002 139576 267058 139632
rect 266542 93064 266598 93120
rect 265346 35264 265402 35320
rect 264150 6704 264206 6760
rect 262954 6568 263010 6624
rect 268934 117952 268990 118008
rect 267738 108296 267794 108352
rect 270130 106800 270186 106856
rect 271142 105440 271198 105496
rect 274914 97280 274970 97336
rect 273718 95784 273774 95840
rect 271326 94424 271382 94480
rect 273902 85856 273958 85912
rect 271142 85720 271198 85776
rect 267186 46280 267242 46336
rect 267186 3984 267242 4040
rect 268842 3984 268898 4040
rect 267002 3168 267058 3224
rect 265346 3032 265402 3088
rect 264978 2896 265034 2952
rect 271142 3168 271198 3224
rect 272430 3168 272486 3224
rect 273902 3168 273958 3224
rect 277306 137536 277362 137592
rect 276110 137400 276166 137456
rect 278502 104216 278558 104272
rect 280342 236000 280398 236056
rect 280250 234640 280306 234696
rect 280158 137264 280214 137320
rect 280526 224984 280582 225040
rect 280434 222808 280490 222864
rect 280250 136312 280306 136368
rect 280802 216688 280858 216744
rect 280618 213152 280674 213208
rect 280526 139984 280582 140040
rect 280434 134680 280490 134736
rect 280618 129104 280674 129160
rect 280066 102720 280122 102776
rect 278042 32408 278098 32464
rect 277858 3984 277914 4040
rect 280986 205672 281042 205728
rect 281170 204176 281226 204232
rect 280986 3848 281042 3904
rect 280802 3712 280858 3768
rect 281354 196016 281410 196072
rect 281814 237632 281870 237688
rect 281722 235184 281778 235240
rect 281630 233552 281686 233608
rect 281538 140528 281594 140584
rect 281998 233280 282054 233336
rect 281906 231104 281962 231160
rect 281906 216688 281962 216744
rect 281906 212608 281962 212664
rect 281814 139576 281870 139632
rect 281722 137128 281778 137184
rect 281630 134816 281686 134872
rect 282182 229200 282238 229256
rect 282274 227840 282330 227896
rect 282090 225256 282146 225312
rect 281998 205672 282054 205728
rect 281998 203224 282054 203280
rect 281906 116592 281962 116648
rect 282182 220904 282238 220960
rect 282458 219816 282514 219872
rect 282366 218048 282422 218104
rect 282826 219444 282828 219464
rect 282828 219444 282880 219464
rect 282880 219444 282882 219464
rect 282826 219408 282882 219444
rect 282826 211656 282882 211712
rect 282826 204856 282882 204912
rect 282458 204176 282514 204232
rect 282366 196016 282422 196072
rect 282274 193296 282330 193352
rect 282366 190576 282422 190632
rect 282458 178084 282514 178120
rect 282458 178064 282460 178084
rect 282460 178064 282512 178084
rect 282512 178064 282514 178084
rect 282826 176840 282882 176896
rect 284298 360984 284354 361040
rect 283194 270408 283250 270464
rect 283562 283600 283618 283656
rect 283470 282648 283526 282704
rect 283654 281016 283710 281072
rect 283378 280064 283434 280120
rect 283286 268912 283342 268968
rect 283102 267280 283158 267336
rect 283010 255040 283066 255096
rect 285862 238856 285918 238912
rect 283102 230560 283158 230616
rect 283010 190984 283066 191040
rect 282918 173576 282974 173632
rect 282826 172216 282882 172272
rect 282734 171808 282790 171864
rect 282826 170720 282882 170776
rect 282826 169668 282828 169688
rect 282828 169668 282880 169688
rect 282880 169668 282882 169688
rect 282826 169632 282882 169668
rect 282826 169224 282882 169280
rect 282826 168136 282882 168192
rect 282734 167728 282790 167784
rect 282274 133184 282330 133240
rect 281998 108432 282054 108488
rect 282182 43560 282238 43616
rect 281354 3984 281410 4040
rect 281170 3576 281226 3632
rect 284482 229472 284538 229528
rect 283286 222264 283342 222320
rect 283194 213968 283250 214024
rect 283102 123528 283158 123584
rect 283378 221312 283434 221368
rect 283470 216688 283526 216744
rect 283562 215600 283618 215656
rect 283470 136176 283526 136232
rect 284390 215328 284446 215384
rect 283654 207440 283710 207496
rect 283562 136040 283618 136096
rect 284298 193568 284354 193624
rect 283654 134544 283710 134600
rect 283286 129240 283342 129296
rect 283194 111016 283250 111072
rect 284666 227024 284722 227080
rect 284574 202952 284630 203008
rect 284482 124888 284538 124944
rect 284390 109656 284446 109712
rect 284758 226344 284814 226400
rect 284850 223624 284906 223680
rect 284758 131960 284814 132016
rect 285034 208936 285090 208992
rect 284850 131824 284906 131880
rect 284666 126384 284722 126440
rect 285770 197376 285826 197432
rect 285678 196016 285734 196072
rect 285034 119448 285090 119504
rect 284574 98776 284630 98832
rect 284298 50224 284354 50280
rect 285954 231920 286010 231976
rect 285862 137944 285918 138000
rect 286046 204312 286102 204368
rect 285954 133320 286010 133376
rect 286322 201728 286378 201784
rect 286138 200368 286194 200424
rect 286046 123392 286102 123448
rect 286230 199280 286286 199336
rect 286414 198736 286470 198792
rect 286322 131688 286378 131744
rect 286506 197648 286562 197704
rect 286414 130328 286470 130384
rect 287518 207168 287574 207224
rect 287426 206352 287482 206408
rect 286506 128968 286562 129024
rect 286230 124752 286286 124808
rect 286138 119312 286194 119368
rect 287886 340312 287942 340368
rect 288438 217776 288494 217832
rect 287794 188400 287850 188456
rect 287610 187584 287666 187640
rect 287702 186768 287758 186824
rect 287886 185952 287942 186008
rect 287794 122032 287850 122088
rect 287702 120672 287758 120728
rect 287610 104080 287666 104136
rect 287886 101360 287942 101416
rect 287518 100136 287574 100192
rect 287426 90344 287482 90400
rect 285770 32544 285826 32600
rect 285678 21392 285734 21448
rect 283010 14728 283066 14784
rect 286598 6160 286654 6216
rect 283102 4800 283158 4856
rect 277858 3440 277914 3496
rect 278042 3440 278098 3496
rect 279514 3440 279570 3496
rect 282182 3440 282238 3496
rect 276018 3168 276074 3224
rect 275282 3032 275338 3088
rect 288806 274896 288862 274952
rect 288806 140256 288862 140312
rect 289818 190032 289874 190088
rect 289082 181056 289138 181112
rect 289082 139440 289138 139496
rect 290094 250280 290150 250336
rect 290002 141752 290058 141808
rect 289910 141616 289966 141672
rect 290186 249464 290242 249520
rect 290278 247832 290334 247888
rect 290370 240624 290426 240680
rect 290278 141344 290334 141400
rect 290370 139848 290426 139904
rect 290186 139168 290242 139224
rect 295062 362480 295118 362536
rect 291474 340176 291530 340232
rect 291658 247016 291714 247072
rect 291658 140120 291714 140176
rect 290094 138352 290150 138408
rect 289818 49136 289874 49192
rect 289082 49000 289138 49056
rect 290186 9016 290242 9072
rect 288438 3304 288494 3360
rect 289082 3304 289138 3360
rect 292670 251232 292726 251288
rect 305826 382744 305882 382800
rect 309414 356904 309470 356960
rect 313002 352552 313058 352608
rect 320178 355408 320234 355464
rect 316590 351328 316646 351384
rect 302238 345888 302294 345944
rect 327354 357992 327410 358048
rect 323766 344936 323822 344992
rect 334530 386688 334586 386744
rect 330942 342760 330998 342816
rect 341706 386824 341762 386880
rect 348882 387640 348938 387696
rect 356058 387504 356114 387560
rect 366822 369280 366878 369336
rect 363234 367648 363290 367704
rect 359646 344800 359702 344856
rect 370410 344664 370466 344720
rect 377586 381656 377642 381712
rect 384762 377168 384818 377224
rect 388350 373360 388406 373416
rect 381174 371864 381230 371920
rect 392582 387096 392638 387152
rect 391938 359488 391994 359544
rect 373998 344528 374054 344584
rect 352470 343304 352526 343360
rect 395526 370640 395582 370696
rect 402702 366288 402758 366344
rect 409878 365064 409934 365120
rect 406290 360848 406346 360904
rect 399114 344392 399170 344448
rect 417422 387504 417478 387560
rect 417054 378800 417110 378856
rect 413466 344256 413522 344312
rect 392582 343168 392638 343224
rect 420642 387368 420698 387424
rect 424230 376216 424286 376272
rect 431406 387232 431462 387288
rect 427818 362344 427874 362400
rect 452934 387640 452990 387696
rect 449346 387504 449402 387560
rect 442170 387096 442226 387152
rect 438582 386960 438638 387016
rect 454682 386824 454738 386880
rect 456522 386824 456578 386880
rect 452934 384240 452990 384296
rect 454682 363704 454738 363760
rect 434994 356768 435050 356824
rect 458178 355952 458234 356008
rect 456798 347656 456854 347712
rect 417422 343032 417478 343088
rect 345294 342624 345350 342680
rect 338118 342488 338174 342544
rect 298650 340040 298706 340096
rect 453302 339360 453358 339416
rect 456798 339360 456854 339416
rect 447782 332424 447838 332480
rect 453302 332424 453358 332480
rect 456062 326984 456118 327040
rect 457442 326984 457498 327040
rect 454682 318688 454738 318744
rect 456062 318688 456118 318744
rect 442262 270408 442318 270464
rect 447782 270408 447838 270464
rect 451922 253136 451978 253192
rect 454682 253136 454738 253192
rect 440882 238720 440938 238776
rect 442262 238720 442318 238776
rect 439502 231784 439558 231840
rect 440882 231784 440938 231840
rect 450542 224848 450598 224904
rect 451922 224848 451978 224904
rect 449162 204176 449218 204232
rect 450542 204176 450598 204232
rect 445390 198736 445446 198792
rect 449162 198736 449218 198792
rect 442906 194792 442962 194848
rect 445390 194792 445446 194848
rect 436006 191664 436062 191720
rect 439502 191664 439558 191720
rect 434626 187720 434682 187776
rect 429198 185544 429254 185600
rect 428462 184864 428518 184920
rect 426438 183096 426494 183152
rect 442906 190440 442962 190496
rect 436098 190304 436154 190360
rect 436098 187720 436154 187776
rect 436006 185544 436062 185600
rect 434626 184864 434682 184920
rect 429198 183096 429254 183152
rect 427082 179424 427138 179480
rect 428462 179424 428518 179480
rect 425702 176024 425758 176080
rect 421562 175888 421618 175944
rect 421562 166368 421618 166424
rect 427082 176024 427138 176080
rect 426346 175888 426402 175944
rect 425702 165552 425758 165608
rect 292670 141888 292726 141944
rect 462962 368328 463018 368384
rect 462962 358944 463018 359000
rect 459558 358672 459614 358728
rect 462318 357312 462374 357368
rect 459558 355952 459614 356008
rect 458914 350376 458970 350432
rect 462318 350376 462374 350432
rect 467102 377984 467158 378040
rect 465078 371456 465134 371512
rect 467102 371456 467158 371512
rect 464342 371184 464398 371240
rect 464986 368328 465042 368384
rect 464342 357312 464398 357368
rect 463698 348472 463754 348528
rect 458914 347656 458970 347712
rect 469218 382744 469274 382800
rect 469218 377984 469274 378040
rect 467838 375400 467894 375456
rect 467838 371320 467894 371376
rect 473174 388728 473230 388784
rect 473358 388728 473414 388784
rect 473266 388456 473322 388512
rect 473174 388184 473230 388240
rect 471242 384648 471298 384704
rect 473542 388456 473598 388512
rect 473266 384648 473322 384704
rect 471242 375400 471298 375456
rect 479614 411848 479670 411904
rect 479614 403008 479670 403064
rect 476118 389136 476174 389192
rect 479522 389136 479578 389192
rect 476118 388456 476174 388512
rect 474646 387776 474702 387832
rect 479890 501608 479946 501664
rect 480074 517520 480130 517576
rect 480166 516840 480222 516896
rect 479982 479848 480038 479904
rect 480350 474408 480406 474464
rect 484122 657192 484178 657248
rect 484030 600208 484086 600264
rect 484214 657056 484270 657112
rect 484122 599936 484178 599992
rect 484306 655560 484362 655616
rect 484214 562944 484270 563000
rect 482282 554512 482338 554568
rect 481730 550432 481786 550488
rect 480442 474000 480498 474056
rect 480258 465704 480314 465760
rect 480534 405592 480590 405648
rect 479798 405184 479854 405240
rect 480626 404232 480682 404288
rect 480810 403688 480866 403744
rect 480718 402872 480774 402928
rect 481086 532072 481142 532128
rect 481638 523096 481694 523152
rect 481822 542272 481878 542328
rect 482006 536424 482062 536480
rect 481914 533840 481970 533896
rect 481822 514664 481878 514720
rect 481730 513304 481786 513360
rect 481638 511808 481694 511864
rect 482098 530440 482154 530496
rect 482190 523640 482246 523696
rect 482006 515208 482062 515264
rect 481914 511536 481970 511592
rect 482190 515752 482246 515808
rect 482190 514800 482246 514856
rect 481638 507048 481694 507104
rect 482098 479304 482154 479360
rect 482098 478216 482154 478272
rect 482098 474700 482154 474736
rect 482098 474680 482100 474700
rect 482100 474680 482152 474700
rect 482152 474680 482154 474700
rect 482098 472232 482154 472288
rect 482006 471688 482062 471744
rect 482098 471144 482154 471200
rect 482006 470328 482062 470384
rect 482098 469512 482154 469568
rect 482098 468968 482154 469024
rect 482006 468560 482062 468616
rect 482006 467764 482062 467800
rect 482006 467744 482008 467764
rect 482008 467744 482060 467764
rect 482060 467744 482062 467764
rect 482098 466792 482154 466848
rect 482098 464924 482100 464944
rect 482100 464924 482152 464944
rect 482152 464924 482154 464944
rect 482098 464888 482154 464924
rect 482006 464616 482062 464672
rect 482098 464072 482154 464128
rect 482098 463392 482154 463448
rect 482098 462984 482154 463040
rect 482098 462032 482154 462088
rect 482006 461896 482062 461952
rect 481914 461352 481970 461408
rect 482098 460672 482154 460728
rect 482098 459312 482154 459368
rect 482006 458632 482062 458688
rect 482098 457952 482154 458008
rect 482006 457544 482062 457600
rect 482098 456592 482154 456648
rect 482098 455268 482100 455288
rect 482100 455268 482152 455288
rect 482152 455268 482154 455288
rect 482098 455232 482154 455268
rect 482006 454824 482062 454880
rect 482098 453736 482154 453792
rect 482098 452548 482100 452568
rect 482100 452548 482152 452568
rect 482152 452548 482154 452568
rect 482098 452512 482154 452548
rect 482098 451560 482154 451616
rect 483754 554104 483810 554160
rect 483202 550160 483258 550216
rect 482558 523504 482614 523560
rect 482374 522144 482430 522200
rect 482466 520920 482522 520976
rect 482374 514120 482430 514176
rect 482374 511944 482430 512000
rect 482282 510856 482338 510912
rect 482282 510448 482338 510504
rect 482190 449928 482246 449984
rect 482190 449828 482192 449848
rect 482192 449828 482244 449848
rect 482244 449828 482246 449848
rect 482190 449792 482246 449828
rect 482098 449384 482154 449440
rect 482190 448840 482246 448896
rect 482190 448296 482246 448352
rect 482098 447888 482154 447944
rect 482006 446664 482062 446720
rect 482190 446956 482246 446992
rect 482190 446936 482192 446956
rect 482192 446936 482244 446956
rect 482244 446936 482246 446956
rect 482098 446120 482154 446176
rect 482190 445440 482246 445496
rect 482098 445168 482154 445224
rect 482190 444216 482246 444272
rect 482098 443944 482154 444000
rect 482190 442720 482246 442776
rect 482098 441224 482154 441280
rect 482190 440680 482246 440736
rect 482190 440000 482246 440056
rect 482190 438796 482246 438832
rect 482190 438776 482192 438796
rect 482192 438776 482244 438796
rect 482244 438776 482246 438796
rect 482098 438504 482154 438560
rect 482190 424496 482246 424552
rect 482190 417288 482246 417344
rect 482190 414568 482246 414624
rect 482190 413616 482246 413672
rect 481086 412936 481142 412992
rect 482190 411032 482246 411088
rect 482190 410760 482246 410816
rect 482190 408348 482192 408368
rect 482192 408348 482244 408368
rect 482244 408348 482246 408368
rect 482190 408312 482246 408348
rect 480994 408176 481050 408232
rect 482190 406544 482246 406600
rect 480902 402600 480958 402656
rect 482190 399336 482246 399392
rect 482006 398384 482062 398440
rect 482190 397704 482246 397760
rect 482190 396616 482246 396672
rect 482190 395664 482246 395720
rect 482190 393896 482246 393952
rect 482098 392264 482154 392320
rect 482190 388320 482246 388376
rect 479798 388184 479854 388240
rect 482282 387640 482338 387696
rect 477498 386008 477554 386064
rect 479706 386008 479762 386064
rect 477498 382744 477554 382800
rect 474462 355272 474518 355328
rect 482926 520784 482982 520840
rect 483018 519016 483074 519072
rect 483018 517520 483074 517576
rect 482926 514800 482982 514856
rect 482558 513032 482614 513088
rect 482466 510312 482522 510368
rect 482466 495488 482522 495544
rect 483018 510448 483074 510504
rect 482650 508544 482706 508600
rect 482926 506232 482982 506288
rect 482834 506096 482890 506152
rect 482926 500520 482982 500576
rect 482834 499976 482890 500032
rect 482834 494672 482890 494728
rect 482742 491952 482798 492008
rect 482926 491816 482982 491872
rect 482834 424768 482890 424824
rect 482834 423408 482890 423464
rect 482834 423308 482836 423328
rect 482836 423308 482888 423328
rect 482888 423308 482890 423328
rect 482834 423272 482890 423308
rect 482834 417968 482890 418024
rect 482834 416608 482890 416664
rect 482834 415112 482890 415168
rect 482834 413752 482890 413808
rect 482834 412392 482890 412448
rect 482834 410352 482890 410408
rect 482834 409536 482890 409592
rect 482834 407496 482890 407552
rect 482834 406816 482890 406872
rect 482834 404776 482890 404832
rect 482834 402056 482890 402112
rect 482834 401376 482890 401432
rect 482834 400968 482890 401024
rect 482834 399880 482890 399936
rect 482834 398692 482836 398712
rect 482836 398692 482888 398712
rect 482888 398692 482890 398712
rect 482834 398656 482890 398692
rect 482834 397160 482890 397216
rect 482834 395800 482890 395856
rect 482834 394304 482890 394360
rect 482834 393252 482836 393272
rect 482836 393252 482888 393272
rect 482888 393252 482890 393272
rect 482834 393216 482890 393252
rect 483294 541864 483350 541920
rect 483202 426672 483258 426728
rect 483478 538872 483534 538928
rect 483386 537784 483442 537840
rect 483570 535336 483626 535392
rect 483662 530304 483718 530360
rect 483846 545808 483902 545864
rect 483754 437008 483810 437064
rect 483662 436192 483718 436248
rect 483570 432112 483626 432168
rect 483478 430752 483534 430808
rect 483386 428304 483442 428360
rect 483294 426128 483350 426184
rect 485962 640736 486018 640792
rect 485778 638968 485834 639024
rect 485134 558456 485190 558512
rect 484398 551520 484454 551576
rect 484306 532072 484362 532128
rect 484490 548664 484546 548720
rect 484398 431024 484454 431080
rect 484582 543224 484638 543280
rect 484490 429392 484546 429448
rect 484674 540640 484730 540696
rect 484766 537920 484822 537976
rect 484950 532208 485006 532264
rect 484858 526768 484914 526824
rect 484766 436464 484822 436520
rect 484674 429936 484730 429992
rect 484582 428848 484638 428904
rect 485042 525272 485098 525328
rect 484950 434832 485006 434888
rect 485778 545128 485834 545184
rect 485226 523912 485282 523968
rect 485226 503376 485282 503432
rect 485134 494672 485190 494728
rect 485962 479984 486018 480040
rect 485042 432656 485098 432712
rect 484858 428032 484914 428088
rect 483846 421504 483902 421560
rect 486330 544584 486386 544640
rect 486238 541728 486294 541784
rect 486422 533704 486478 533760
rect 486330 435376 486386 435432
rect 486514 529624 486570 529680
rect 486422 433472 486478 433528
rect 486606 526904 486662 526960
rect 501786 657736 501842 657792
rect 486974 599800 487030 599856
rect 497646 655968 497702 656024
rect 494886 655832 494942 655888
rect 492126 655560 492182 655616
rect 496266 655696 496322 655752
rect 503166 657192 503222 657248
rect 508502 657328 508558 657384
rect 504546 657056 504602 657112
rect 514206 657600 514262 657656
rect 534906 657600 534962 657656
rect 515586 657464 515642 657520
rect 532146 657464 532202 657520
rect 529386 657328 529442 657384
rect 530766 657192 530822 657248
rect 536286 657056 536342 657112
rect 537666 656920 537722 656976
rect 493506 654608 493562 654664
rect 488446 654472 488502 654528
rect 500406 654472 500462 654528
rect 487526 640600 487582 640656
rect 487158 637608 487214 637664
rect 487158 613672 487214 613728
rect 487158 559000 487214 559056
rect 487710 551248 487766 551304
rect 487526 475088 487582 475144
rect 486606 433744 486662 433800
rect 486514 431568 486570 431624
rect 486238 422048 486294 422104
rect 490746 654200 490802 654256
rect 540242 652840 540298 652896
rect 488998 641824 489054 641880
rect 488538 641688 488594 641744
rect 488722 639920 488778 639976
rect 488538 637608 488594 637664
rect 488446 600072 488502 600128
rect 488906 639104 488962 639160
rect 488998 476720 489054 476776
rect 488906 472912 488962 472968
rect 488722 469648 488778 469704
rect 487710 408720 487766 408776
rect 489182 525136 489238 525192
rect 539782 630536 539838 630592
rect 539598 627816 539654 627872
rect 539506 612720 539562 612776
rect 539414 610680 539470 610736
rect 539322 604424 539378 604480
rect 539414 601840 539470 601896
rect 539506 601704 539562 601760
rect 497370 600208 497426 600264
rect 490378 547168 490434 547224
rect 490286 543088 490342 543144
rect 489182 425584 489238 425640
rect 490470 536288 490526 536344
rect 490470 437688 490526 437744
rect 490378 434424 490434 434480
rect 490286 425176 490342 425232
rect 482926 392808 482982 392864
rect 482926 391584 482982 391640
rect 482834 391176 482890 391232
rect 482926 390360 482982 390416
rect 482834 386280 482890 386336
rect 482742 383288 482798 383344
rect 482466 342896 482522 342952
rect 495714 599528 495770 599584
rect 492126 598168 492182 598224
rect 493506 598168 493562 598224
rect 494886 598168 494942 598224
rect 494610 558728 494666 558784
rect 492126 549888 492182 549944
rect 491574 526496 491630 526552
rect 491942 546352 491998 546408
rect 492034 520104 492090 520160
rect 491942 509496 491998 509552
rect 492034 491544 492090 491600
rect 492126 422456 492182 422512
rect 491574 417560 491630 417616
rect 494610 490456 494666 490512
rect 495622 526360 495678 526416
rect 496082 535064 496138 535120
rect 495990 521328 496046 521384
rect 495806 520104 495862 520160
rect 495714 491952 495770 492008
rect 495622 418648 495678 418704
rect 496082 499160 496138 499216
rect 495990 478488 496046 478544
rect 495806 415384 495862 415440
rect 496818 522280 496874 522336
rect 496818 508408 496874 508464
rect 497646 598168 497702 598224
rect 497370 491816 497426 491872
rect 497646 521600 497702 521656
rect 498382 531936 498438 531992
rect 498566 527856 498622 527912
rect 498750 522008 498806 522064
rect 498750 477400 498806 477456
rect 498566 419736 498622 419792
rect 498382 405048 498438 405104
rect 497462 363568 497518 363624
rect 496266 354048 496322 354104
rect 492586 278024 492642 278080
rect 482374 164736 482430 164792
rect 311438 86128 311494 86184
rect 293682 3440 293738 3496
rect 304354 51856 304410 51912
rect 297270 42200 297326 42256
rect 300766 3304 300822 3360
rect 307942 4936 307998 4992
rect 329194 85584 329250 85640
rect 315026 80688 315082 80744
rect 322110 79328 322166 79384
rect 318522 53080 318578 53136
rect 325606 54576 325662 54632
rect 343362 84632 343418 84688
rect 334622 58520 334678 58576
rect 332690 7520 332746 7576
rect 334622 7520 334678 7576
rect 499578 599664 499634 599720
rect 499026 359352 499082 359408
rect 497462 298696 497518 298752
rect 499762 536152 499818 536208
rect 499946 530848 500002 530904
rect 499762 419192 499818 419248
rect 500222 457408 500278 457464
rect 499946 420280 500002 420336
rect 500222 390088 500278 390144
rect 501234 525000 501290 525056
rect 501326 522688 501382 522744
rect 501418 521192 501474 521248
rect 501510 519696 501566 519752
rect 501510 482296 501566 482352
rect 501418 480664 501474 480720
rect 501326 476312 501382 476368
rect 501234 427352 501290 427408
rect 500406 380024 500462 380080
rect 502706 522552 502762 522608
rect 502706 472504 502762 472560
rect 501786 364928 501842 364984
rect 503074 511944 503130 512000
rect 503074 389000 503130 389056
rect 504086 599936 504142 599992
rect 503810 562944 503866 563000
rect 503166 374584 503222 374640
rect 504178 564304 504234 564360
rect 504178 562944 504234 563000
rect 504086 511944 504142 512000
rect 504086 511264 504142 511320
rect 504362 521464 504418 521520
rect 504362 481752 504418 481808
rect 503810 388864 503866 388920
rect 505466 555872 505522 555928
rect 505558 521056 505614 521112
rect 505466 502968 505522 503024
rect 505558 481208 505614 481264
rect 505926 383016 505982 383072
rect 506938 540504 506994 540560
rect 506938 494808 506994 494864
rect 504546 345616 504602 345672
rect 507858 600072 507914 600128
rect 508042 599800 508098 599856
rect 507950 532072 508006 532128
rect 507858 405184 507914 405240
rect 508042 457408 508098 457464
rect 508686 382880 508742 382936
rect 510066 380840 510122 380896
rect 511906 598984 511962 599040
rect 511906 485832 511962 485888
rect 512826 380704 512882 380760
rect 515586 380568 515642 380624
rect 516966 380432 517022 380488
rect 514206 380296 514262 380352
rect 519726 380160 519782 380216
rect 523682 598304 523738 598360
rect 522486 377712 522542 377768
rect 521106 377440 521162 377496
rect 518346 369144 518402 369200
rect 525246 377848 525302 377904
rect 523866 377576 523922 377632
rect 529202 598032 529258 598088
rect 528006 378664 528062 378720
rect 526626 377304 526682 377360
rect 523682 369008 523738 369064
rect 511446 362208 511502 362264
rect 531962 599800 532018 599856
rect 532146 598304 532202 598360
rect 531962 386144 532018 386200
rect 533526 375944 533582 376000
rect 530766 351192 530822 351248
rect 529202 349832 529258 349888
rect 536010 600208 536066 600264
rect 535734 599120 535790 599176
rect 536102 383424 536158 383480
rect 534906 348336 534962 348392
rect 536838 598984 536894 599040
rect 538586 600072 538642 600128
rect 537666 598032 537722 598088
rect 536286 347112 536342 347168
rect 507950 346976 508006 347032
rect 539690 625096 539746 625152
rect 539598 331744 539654 331800
rect 539966 622376 540022 622432
rect 539874 621016 539930 621072
rect 539782 338816 539838 338872
rect 539690 330384 539746 330440
rect 507858 278024 507914 278080
rect 499578 163920 499634 163976
rect 559654 700304 559710 700360
rect 545118 657328 545174 657384
rect 543738 657192 543794 657248
rect 543462 652840 543518 652896
rect 542358 651208 542414 651264
rect 541162 641688 541218 641744
rect 541070 640328 541126 640384
rect 540978 638968 541034 639024
rect 541254 637608 541310 637664
rect 541162 383152 541218 383208
rect 541346 634888 541402 634944
rect 542818 649848 542874 649904
rect 542450 648488 542506 648544
rect 542358 598304 542414 598360
rect 542634 647128 542690 647184
rect 542542 645768 542598 645824
rect 542450 598168 542506 598224
rect 542726 643048 542782 643104
rect 542910 644408 542966 644464
rect 542818 612720 542874 612776
rect 543370 615848 543426 615904
rect 543002 614488 543058 614544
rect 542910 610680 542966 610736
rect 542542 596808 542598 596864
rect 543186 613128 543242 613184
rect 543094 611768 543150 611824
rect 543094 601024 543150 601080
rect 543186 600208 543242 600264
rect 543002 594768 543058 594824
rect 543370 593408 543426 593464
rect 541346 384376 541402 384432
rect 543922 656920 543978 656976
rect 543922 600208 543978 600264
rect 545210 657056 545266 657112
rect 545210 599800 545266 599856
rect 580262 697176 580318 697232
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 546590 657600 546646 657656
rect 545118 388592 545174 388648
rect 546682 657464 546738 657520
rect 546682 384920 546738 384976
rect 546590 384784 546646 384840
rect 580170 617516 580172 617536
rect 580172 617516 580224 617536
rect 580224 617516 580226 617536
rect 580170 617480 580226 617516
rect 543738 383560 543794 383616
rect 541254 380976 541310 381032
rect 580354 644000 580410 644056
rect 580262 373224 580318 373280
rect 580170 351872 580226 351928
rect 580446 590960 580502 591016
rect 580538 537784 580594 537840
rect 580446 353912 580502 353968
rect 580630 431568 580686 431624
rect 580630 356632 580686 356688
rect 580538 351056 580594 351112
rect 580262 325216 580318 325272
rect 541070 322224 541126 322280
rect 540978 321408 541034 321464
rect 580262 272176 580318 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 205672 580226 205728
rect 580170 165824 580226 165880
rect 540242 163104 540298 163160
rect 580354 232328 580410 232384
rect 580446 192480 580502 192536
rect 580538 152632 580594 152688
rect 580262 135904 580318 135960
rect 492586 86128 492642 86184
rect 364614 84904 364670 84960
rect 357530 84768 357586 84824
rect 355322 55800 355378 55856
rect 355322 4800 355378 4856
rect 361118 84496 361174 84552
rect 432602 83000 432658 83056
rect 428554 81640 428610 81696
rect 421562 78920 421618 78976
rect 417422 77560 417478 77616
rect 414662 76200 414718 76256
rect 410522 74840 410578 74896
rect 400126 40704 400182 40760
rect 393042 24248 393098 24304
rect 382370 20032 382426 20088
rect 378874 13096 378930 13152
rect 375286 11736 375342 11792
rect 389454 15952 389510 16008
rect 385958 14592 386014 14648
rect 396538 17312 396594 17368
rect 403622 39344 403678 39400
rect 407210 18672 407266 18728
rect 411902 57160 411958 57216
rect 410798 4800 410854 4856
rect 411902 4800 411958 4856
rect 414294 4800 414350 4856
rect 410522 3576 410578 3632
rect 418802 59880 418858 59936
rect 417882 7520 417938 7576
rect 417422 3440 417478 3496
rect 414662 3032 414718 3088
rect 418802 4120 418858 4176
rect 421378 4120 421434 4176
rect 425702 68040 425758 68096
rect 422942 61240 422998 61296
rect 427082 62600 427138 62656
rect 425702 7520 425758 7576
rect 422942 4120 422998 4176
rect 424966 4120 425022 4176
rect 427082 4120 427138 4176
rect 428462 4120 428518 4176
rect 421562 3848 421618 3904
rect 431222 65320 431278 65376
rect 429842 63960 429898 64016
rect 431222 4936 431278 4992
rect 429842 4800 429898 4856
rect 432050 4800 432106 4856
rect 428554 3712 428610 3768
rect 450542 73480 450598 73536
rect 446402 72120 446458 72176
rect 443642 70760 443698 70816
rect 436742 66680 436798 66736
rect 435362 47776 435418 47832
rect 435546 4936 435602 4992
rect 435362 3984 435418 4040
rect 432602 3168 432658 3224
rect 439502 47640 439558 47696
rect 436742 4120 436798 4176
rect 439134 4120 439190 4176
rect 438858 3984 438914 4040
rect 442262 47504 442318 47560
rect 442630 7520 442686 7576
rect 439502 3304 439558 3360
rect 580262 72936 580318 72992
rect 471058 51720 471114 51776
rect 450542 4800 450598 4856
rect 453302 4800 453358 4856
rect 443642 4120 443698 4176
rect 446218 4120 446274 4176
rect 446402 4120 446458 4176
rect 449806 4120 449862 4176
rect 467470 3848 467526 3904
rect 456890 3576 456946 3632
rect 463974 3440 464030 3496
rect 460386 3032 460442 3088
rect 545486 48864 545542 48920
rect 481730 46144 481786 46200
rect 474554 3712 474610 3768
rect 478142 3168 478198 3224
rect 499394 43424 499450 43480
rect 495898 12960 495954 13016
rect 492310 11600 492366 11656
rect 488814 10240 488870 10296
rect 485226 8880 485282 8936
rect 506478 42064 506534 42120
rect 502982 19896 503038 19952
rect 512642 40568 512698 40624
rect 508502 14456 508558 14512
rect 508502 3984 508558 4040
rect 510066 3984 510122 4040
rect 520738 39208 520794 39264
rect 517150 17176 517206 17232
rect 512642 3440 512698 3496
rect 513562 3440 513618 3496
rect 524234 37848 524290 37904
rect 531318 36488 531374 36544
rect 527822 18536 527878 18592
rect 534906 35128 534962 35184
rect 538402 33768 538458 33824
rect 541990 30912 542046 30968
rect 549074 44784 549130 44840
rect 552662 29552 552718 29608
rect 559746 28192 559802 28248
rect 556158 24112 556214 24168
rect 562322 26832 562378 26888
rect 566830 25472 566886 25528
rect 562322 3440 562378 3496
rect 563242 3440 563298 3496
rect 573914 22616 573970 22672
rect 570326 21256 570382 21312
rect 576122 15816 576178 15872
rect 580170 6568 580226 6624
rect 576122 3984 576178 4040
rect 577410 3984 577466 4040
rect 582194 3304 582250 3360
<< metal3 >>
rect 176929 700498 176995 700501
rect 218973 700498 219039 700501
rect 176929 700496 219039 700498
rect 176929 700440 176934 700496
rect 176990 700440 218978 700496
rect 219034 700440 219039 700496
rect 176929 700438 219039 700440
rect 176929 700435 176995 700438
rect 218973 700435 219039 700438
rect 413645 700498 413711 700501
rect 483054 700498 483060 700500
rect 413645 700496 483060 700498
rect 413645 700440 413650 700496
rect 413706 700440 483060 700496
rect 413645 700438 483060 700440
rect 413645 700435 413711 700438
rect 483054 700436 483060 700438
rect 483124 700436 483130 700500
rect 24301 700362 24367 700365
rect 32397 700362 32463 700365
rect 24301 700360 32463 700362
rect 24301 700304 24306 700360
rect 24362 700304 32402 700360
rect 32458 700304 32463 700360
rect 24301 700302 32463 700304
rect 24301 700299 24367 700302
rect 32397 700299 32463 700302
rect 55990 700300 55996 700364
rect 56060 700362 56066 700364
rect 89161 700362 89227 700365
rect 56060 700360 89227 700362
rect 56060 700304 89166 700360
rect 89222 700304 89227 700360
rect 56060 700302 89227 700304
rect 56060 700300 56066 700302
rect 89161 700299 89227 700302
rect 160093 700362 160159 700365
rect 202781 700362 202847 700365
rect 160093 700360 202847 700362
rect 160093 700304 160098 700360
rect 160154 700304 202786 700360
rect 202842 700304 202847 700360
rect 160093 700302 202847 700304
rect 160093 700299 160159 700302
rect 202781 700299 202847 700302
rect 397453 700362 397519 700365
rect 479558 700362 479564 700364
rect 397453 700360 479564 700362
rect 397453 700304 397458 700360
rect 397514 700304 479564 700360
rect 397453 700302 479564 700304
rect 397453 700299 397519 700302
rect 479558 700300 479564 700302
rect 479628 700300 479634 700364
rect 508497 700362 508563 700365
rect 559649 700362 559715 700365
rect 508497 700360 559715 700362
rect 508497 700304 508502 700360
rect 508558 700304 559654 700360
rect 559710 700304 559715 700360
rect 508497 700302 559715 700304
rect 508497 700299 508563 700302
rect 559649 700299 559715 700302
rect 59118 699756 59124 699820
rect 59188 699818 59194 699820
rect 59261 699818 59327 699821
rect 141417 699818 141483 699821
rect 59188 699816 141483 699818
rect 59188 699760 59266 699816
rect 59322 699760 141422 699816
rect 141478 699760 141483 699816
rect 59188 699758 141483 699760
rect 59188 699756 59194 699758
rect 59261 699755 59327 699758
rect 141417 699755 141483 699758
rect 156597 698322 156663 698325
rect 160093 698322 160159 698325
rect 156597 698320 160159 698322
rect 156597 698264 156602 698320
rect 156658 698264 160098 698320
rect 160154 698264 160159 698320
rect 156597 698262 160159 698264
rect 156597 698259 156663 698262
rect 160093 698259 160159 698262
rect 173157 698322 173223 698325
rect 176929 698322 176995 698325
rect 173157 698320 176995 698322
rect 173157 698264 173162 698320
rect 173218 698264 176934 698320
rect 176990 698264 176995 698320
rect 173157 698262 176995 698264
rect 173157 698259 173223 698262
rect 176929 698259 176995 698262
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect 173157 687306 173223 687309
rect 168422 687304 173223 687306
rect 168422 687248 173162 687304
rect 173218 687248 173223 687304
rect 168422 687246 173223 687248
rect 167637 687170 167703 687173
rect 168422 687170 168482 687246
rect 173157 687243 173223 687246
rect 167637 687168 168482 687170
rect 167637 687112 167642 687168
rect 167698 687112 168482 687168
rect 167637 687110 168482 687112
rect 167637 687107 167703 687110
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 555366 683844 555372 683908
rect 555436 683906 555442 683908
rect 583520 683906 584960 683996
rect 555436 683846 584960 683906
rect 555436 683844 555442 683846
rect 583520 683756 584960 683846
rect 153193 681866 153259 681869
rect 156597 681866 156663 681869
rect 153193 681864 156663 681866
rect 153193 681808 153198 681864
rect 153254 681808 156602 681864
rect 156658 681808 156663 681864
rect 153193 681806 156663 681808
rect 153193 681803 153259 681806
rect 156597 681803 156663 681806
rect 283833 681730 283899 681733
rect 288341 681730 288407 681733
rect 283833 681728 288407 681730
rect 283833 681672 283838 681728
rect 283894 681672 288346 681728
rect 288402 681672 288407 681728
rect 283833 681670 288407 681672
rect 283833 681667 283899 681670
rect 288341 681667 288407 681670
rect 167637 679010 167703 679013
rect 164558 679008 167703 679010
rect 164558 678952 167642 679008
rect 167698 678952 167703 679008
rect 164558 678950 167703 678952
rect 158897 678194 158963 678197
rect 164558 678194 164618 678950
rect 167637 678947 167703 678950
rect 288341 678738 288407 678741
rect 290457 678738 290523 678741
rect 288341 678736 290523 678738
rect 288341 678680 288346 678736
rect 288402 678680 290462 678736
rect 290518 678680 290523 678736
rect 288341 678678 290523 678680
rect 288341 678675 288407 678678
rect 290457 678675 290523 678678
rect 158897 678192 164618 678194
rect 158897 678136 158902 678192
rect 158958 678136 164618 678192
rect 158897 678134 164618 678136
rect 158897 678131 158963 678134
rect 157977 675882 158043 675885
rect 158897 675882 158963 675885
rect 157977 675880 158963 675882
rect 157977 675824 157982 675880
rect 158038 675824 158902 675880
rect 158958 675824 158963 675880
rect 157977 675822 158963 675824
rect 157977 675819 158043 675822
rect 158897 675819 158963 675822
rect -960 671258 480 671348
rect 31702 671258 31708 671260
rect -960 671198 31708 671258
rect -960 671108 480 671198
rect 31702 671196 31708 671198
rect 31772 671196 31778 671260
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 155309 666498 155375 666501
rect 157977 666498 158043 666501
rect 155309 666496 158043 666498
rect 155309 666440 155314 666496
rect 155370 666440 157982 666496
rect 158038 666440 158043 666496
rect 155309 666438 158043 666440
rect 155309 666435 155375 666438
rect 157977 666435 158043 666438
rect 150525 660922 150591 660925
rect 152457 660922 152523 660925
rect 150525 660920 152523 660922
rect 150525 660864 150530 660920
rect 150586 660864 152462 660920
rect 152518 660864 152523 660920
rect 150525 660862 152523 660864
rect 150525 660859 150591 660862
rect 152457 660859 152523 660862
rect -960 658202 480 658292
rect 14406 658202 14412 658204
rect -960 658142 14412 658202
rect -960 658052 480 658142
rect 14406 658140 14412 658142
rect 14476 658140 14482 658204
rect 290457 657794 290523 657797
rect 309777 657794 309843 657797
rect 290457 657792 309843 657794
rect 290457 657736 290462 657792
rect 290518 657736 309782 657792
rect 309838 657736 309843 657792
rect 290457 657734 309843 657736
rect 290457 657731 290523 657734
rect 309777 657731 309843 657734
rect 486969 657794 487035 657797
rect 501781 657794 501847 657797
rect 486969 657792 501847 657794
rect 486969 657736 486974 657792
rect 487030 657736 501786 657792
rect 501842 657736 501847 657792
rect 486969 657734 501847 657736
rect 486969 657731 487035 657734
rect 501781 657731 501847 657734
rect 55070 657596 55076 657660
rect 55140 657658 55146 657660
rect 300117 657658 300183 657661
rect 514201 657658 514267 657661
rect 55140 657656 514267 657658
rect 55140 657600 300122 657656
rect 300178 657600 514206 657656
rect 514262 657600 514267 657656
rect 55140 657598 514267 657600
rect 55140 657596 55146 657598
rect 300117 657595 300183 657598
rect 514201 657595 514267 657598
rect 534901 657658 534967 657661
rect 546585 657658 546651 657661
rect 534901 657656 546651 657658
rect 534901 657600 534906 657656
rect 534962 657600 546590 657656
rect 546646 657600 546651 657656
rect 534901 657598 546651 657600
rect 534901 657595 534967 657598
rect 546585 657595 546651 657598
rect 170990 657460 170996 657524
rect 171060 657522 171066 657524
rect 235165 657522 235231 657525
rect 515581 657522 515647 657525
rect 171060 657520 515647 657522
rect 171060 657464 235170 657520
rect 235226 657464 515586 657520
rect 515642 657464 515647 657520
rect 171060 657462 515647 657464
rect 171060 657460 171066 657462
rect 235165 657459 235231 657462
rect 515581 657459 515647 657462
rect 532141 657522 532207 657525
rect 546677 657522 546743 657525
rect 532141 657520 546743 657522
rect 532141 657464 532146 657520
rect 532202 657464 546682 657520
rect 546738 657464 546743 657520
rect 532141 657462 546743 657464
rect 532141 657459 532207 657462
rect 546677 657459 546743 657462
rect 484025 657386 484091 657389
rect 508497 657386 508563 657389
rect 484025 657384 508563 657386
rect 484025 657328 484030 657384
rect 484086 657328 508502 657384
rect 508558 657328 508563 657384
rect 484025 657326 508563 657328
rect 484025 657323 484091 657326
rect 508497 657323 508563 657326
rect 529381 657386 529447 657389
rect 545113 657386 545179 657389
rect 529381 657384 545179 657386
rect 529381 657328 529386 657384
rect 529442 657328 545118 657384
rect 545174 657328 545179 657384
rect 529381 657326 545179 657328
rect 529381 657323 529447 657326
rect 545113 657323 545179 657326
rect 484117 657250 484183 657253
rect 503161 657250 503227 657253
rect 484117 657248 503227 657250
rect 484117 657192 484122 657248
rect 484178 657192 503166 657248
rect 503222 657192 503227 657248
rect 484117 657190 503227 657192
rect 484117 657187 484183 657190
rect 503161 657187 503227 657190
rect 530761 657250 530827 657253
rect 543733 657250 543799 657253
rect 530761 657248 543799 657250
rect 530761 657192 530766 657248
rect 530822 657192 543738 657248
rect 543794 657192 543799 657248
rect 583520 657236 584960 657476
rect 530761 657190 543799 657192
rect 530761 657187 530827 657190
rect 543733 657187 543799 657190
rect 484209 657114 484275 657117
rect 504541 657114 504607 657117
rect 484209 657112 504607 657114
rect 484209 657056 484214 657112
rect 484270 657056 504546 657112
rect 504602 657056 504607 657112
rect 484209 657054 504607 657056
rect 484209 657051 484275 657054
rect 504541 657051 504607 657054
rect 536281 657114 536347 657117
rect 545205 657114 545271 657117
rect 536281 657112 545271 657114
rect 536281 657056 536286 657112
rect 536342 657056 545210 657112
rect 545266 657056 545271 657112
rect 536281 657054 545271 657056
rect 536281 657051 536347 657054
rect 545205 657051 545271 657054
rect 537661 656978 537727 656981
rect 543917 656978 543983 656981
rect 537661 656976 543983 656978
rect 537661 656920 537666 656976
rect 537722 656920 543922 656976
rect 543978 656920 543983 656976
rect 537661 656918 543983 656920
rect 537661 656915 537727 656918
rect 543917 656915 543983 656918
rect 473261 656026 473327 656029
rect 497641 656026 497707 656029
rect 473261 656024 497707 656026
rect 473261 655968 473266 656024
rect 473322 655968 497646 656024
rect 497702 655968 497707 656024
rect 473261 655966 497707 655968
rect 473261 655963 473327 655966
rect 497641 655963 497707 655966
rect 476021 655890 476087 655893
rect 494881 655890 494947 655893
rect 476021 655888 494947 655890
rect 476021 655832 476026 655888
rect 476082 655832 494886 655888
rect 494942 655832 494947 655888
rect 476021 655830 494947 655832
rect 476021 655827 476087 655830
rect 494881 655827 494947 655830
rect 477401 655754 477467 655757
rect 496261 655754 496327 655757
rect 477401 655752 496327 655754
rect 477401 655696 477406 655752
rect 477462 655696 496266 655752
rect 496322 655696 496327 655752
rect 477401 655694 496327 655696
rect 477401 655691 477467 655694
rect 496261 655691 496327 655694
rect 484301 655618 484367 655621
rect 492121 655618 492187 655621
rect 484301 655616 492187 655618
rect 484301 655560 484306 655616
rect 484362 655560 492126 655616
rect 492182 655560 492187 655616
rect 484301 655558 492187 655560
rect 484301 655555 484367 655558
rect 492121 655555 492187 655558
rect 475929 654666 475995 654669
rect 493501 654666 493567 654669
rect 475929 654664 493567 654666
rect 475929 654608 475934 654664
rect 475990 654608 493506 654664
rect 493562 654608 493567 654664
rect 475929 654606 493567 654608
rect 475929 654603 475995 654606
rect 493501 654603 493567 654606
rect 488441 654530 488507 654533
rect 500401 654530 500467 654533
rect 488441 654528 500467 654530
rect 488441 654472 488446 654528
rect 488502 654472 500406 654528
rect 500462 654472 500467 654528
rect 488441 654470 500467 654472
rect 488441 654467 488507 654470
rect 500401 654467 500467 654470
rect 489862 654196 489868 654260
rect 489932 654258 489938 654260
rect 490741 654258 490807 654261
rect 489932 654256 490807 654258
rect 489932 654200 490746 654256
rect 490802 654200 490807 654256
rect 489932 654198 490807 654200
rect 489932 654196 489938 654198
rect 490741 654195 490807 654198
rect 153561 652898 153627 652901
rect 155309 652898 155375 652901
rect 153561 652896 155375 652898
rect 153561 652840 153566 652896
rect 153622 652840 155314 652896
rect 155370 652840 155375 652896
rect 153561 652838 155375 652840
rect 153561 652835 153627 652838
rect 155309 652835 155375 652838
rect 540237 652898 540303 652901
rect 543457 652898 543523 652901
rect 540237 652896 543523 652898
rect 540237 652840 540242 652896
rect 540298 652840 543462 652896
rect 543518 652840 543523 652896
rect 540237 652838 543523 652840
rect 540237 652835 540303 652838
rect 543457 652835 543523 652838
rect 542353 651266 542419 651269
rect 539948 651264 542419 651266
rect 539948 651208 542358 651264
rect 542414 651208 542419 651264
rect 539948 651206 542419 651208
rect 542353 651203 542419 651206
rect 309777 650314 309843 650317
rect 312905 650314 312971 650317
rect 309777 650312 312971 650314
rect 309777 650256 309782 650312
rect 309838 650256 312910 650312
rect 312966 650256 312971 650312
rect 309777 650254 312971 650256
rect 309777 650251 309843 650254
rect 312905 650251 312971 650254
rect 38561 650178 38627 650181
rect 340045 650178 340111 650181
rect 38561 650176 340111 650178
rect 38561 650120 38566 650176
rect 38622 650120 340050 650176
rect 340106 650120 340111 650176
rect 38561 650118 340111 650120
rect 38561 650115 38627 650118
rect 340045 650115 340111 650118
rect 28901 650042 28967 650045
rect 368381 650042 368447 650045
rect 28901 650040 368447 650042
rect 28901 649984 28906 650040
rect 28962 649984 368386 650040
rect 368442 649984 368447 650040
rect 28901 649982 368447 649984
rect 28901 649979 28967 649982
rect 368381 649979 368447 649982
rect 149697 649906 149763 649909
rect 153561 649906 153627 649909
rect 542813 649906 542879 649909
rect 149697 649904 153627 649906
rect 149697 649848 149702 649904
rect 149758 649848 153566 649904
rect 153622 649848 153627 649904
rect 149697 649846 153627 649848
rect 539948 649904 542879 649906
rect 539948 649848 542818 649904
rect 542874 649848 542879 649904
rect 539948 649846 542879 649848
rect 149697 649843 149763 649846
rect 153561 649843 153627 649846
rect 542813 649843 542879 649846
rect 37181 648682 37247 648685
rect 360653 648682 360719 648685
rect 37181 648680 360719 648682
rect 37181 648624 37186 648680
rect 37242 648624 360658 648680
rect 360714 648624 360719 648680
rect 37181 648622 360719 648624
rect 37181 648619 37247 648622
rect 360653 648619 360719 648622
rect 542445 648546 542511 648549
rect 539948 648544 542511 648546
rect 539948 648488 542450 648544
rect 542506 648488 542511 648544
rect 539948 648486 542511 648488
rect 542445 648483 542511 648486
rect 34421 648410 34487 648413
rect 204897 648410 204963 648413
rect 34421 648408 204963 648410
rect 34421 648352 34426 648408
rect 34482 648352 204902 648408
rect 204958 648352 204963 648408
rect 34421 648350 204963 648352
rect 34421 648347 34487 648350
rect 204897 648347 204963 648350
rect 193029 648274 193095 648277
rect 208393 648274 208459 648277
rect 193029 648272 208459 648274
rect 193029 648216 193034 648272
rect 193090 648216 208398 648272
rect 208454 648216 208459 648272
rect 193029 648214 208459 648216
rect 193029 648211 193095 648214
rect 208393 648211 208459 648214
rect 103881 648138 103947 648141
rect 280797 648138 280863 648141
rect 103881 648136 280863 648138
rect 103881 648080 103886 648136
rect 103942 648080 280802 648136
rect 280858 648080 280863 648136
rect 103881 648078 280863 648080
rect 103881 648075 103947 648078
rect 280797 648075 280863 648078
rect 96153 648002 96219 648005
rect 286317 648002 286383 648005
rect 96153 648000 286383 648002
rect 96153 647944 96158 648000
rect 96214 647944 286322 648000
rect 286378 647944 286383 648000
rect 96153 647942 286383 647944
rect 96153 647939 96219 647942
rect 286317 647939 286383 647942
rect 91001 647866 91067 647869
rect 289261 647866 289327 647869
rect 91001 647864 289327 647866
rect 91001 647808 91006 647864
rect 91062 647808 289266 647864
rect 289322 647808 289327 647864
rect 91001 647806 289327 647808
rect 91001 647803 91067 647806
rect 289261 647803 289327 647806
rect 65241 647730 65307 647733
rect 275277 647730 275343 647733
rect 65241 647728 275343 647730
rect 65241 647672 65246 647728
rect 65302 647672 275282 647728
rect 275338 647672 275343 647728
rect 65241 647670 275343 647672
rect 65241 647667 65307 647670
rect 275277 647667 275343 647670
rect 202045 647594 202111 647597
rect 233141 647594 233207 647597
rect 202045 647592 233207 647594
rect 202045 647536 202050 647592
rect 202106 647536 233146 647592
rect 233202 647536 233207 647592
rect 202045 647534 233207 647536
rect 202045 647531 202111 647534
rect 233141 647531 233207 647534
rect 233417 647594 233483 647597
rect 461669 647594 461735 647597
rect 233417 647592 461735 647594
rect 233417 647536 233422 647592
rect 233478 647536 461674 647592
rect 461730 647536 461735 647592
rect 233417 647534 461735 647536
rect 233417 647531 233483 647534
rect 461669 647531 461735 647534
rect 35801 647458 35867 647461
rect 202781 647458 202847 647461
rect 35801 647456 202847 647458
rect 35801 647400 35806 647456
rect 35862 647400 202786 647456
rect 202842 647400 202847 647456
rect 35801 647398 202847 647400
rect 35801 647395 35867 647398
rect 202781 647395 202847 647398
rect 208485 647458 208551 647461
rect 467281 647458 467347 647461
rect 208485 647456 467347 647458
rect 208485 647400 208490 647456
rect 208546 647400 467286 647456
rect 467342 647400 467347 647456
rect 208485 647398 467347 647400
rect 208485 647395 208551 647398
rect 467281 647395 467347 647398
rect 204621 647322 204687 647325
rect 467097 647322 467163 647325
rect 204621 647320 467163 647322
rect 204621 647264 204626 647320
rect 204682 647264 467102 647320
rect 467158 647264 467163 647320
rect 204621 647262 467163 647264
rect 204621 647259 204687 647262
rect 467097 647259 467163 647262
rect 542629 647186 542695 647189
rect 539948 647184 542695 647186
rect 539948 647128 542634 647184
rect 542690 647128 542695 647184
rect 539948 647126 542695 647128
rect 542629 647123 542695 647126
rect 212349 646914 212415 646917
rect 212349 646912 219450 646914
rect 212349 646856 212354 646912
rect 212410 646856 219450 646912
rect 212349 646854 219450 646856
rect 212349 646851 212415 646854
rect 50797 646778 50863 646781
rect 212441 646778 212507 646781
rect 50797 646776 212507 646778
rect 50797 646720 50802 646776
rect 50858 646720 212446 646776
rect 212502 646720 212507 646776
rect 50797 646718 212507 646720
rect 219390 646778 219450 646854
rect 464337 646778 464403 646781
rect 219390 646776 464403 646778
rect 219390 646720 464342 646776
rect 464398 646720 464403 646776
rect 219390 646718 464403 646720
rect 50797 646715 50863 646718
rect 212441 646715 212507 646718
rect 464337 646715 464403 646718
rect 53741 646642 53807 646645
rect 333605 646642 333671 646645
rect 53741 646640 333671 646642
rect 53741 646584 53746 646640
rect 53802 646584 333610 646640
rect 333666 646584 333671 646640
rect 53741 646582 333671 646584
rect 53741 646579 53807 646582
rect 333605 646579 333671 646582
rect 52177 646506 52243 646509
rect 332317 646506 332383 646509
rect 52177 646504 332383 646506
rect 52177 646448 52182 646504
rect 52238 646448 332322 646504
rect 332378 646448 332383 646504
rect 52177 646446 332383 646448
rect 52177 646443 52243 646446
rect 332317 646443 332383 646446
rect 53649 646370 53715 646373
rect 336181 646370 336247 646373
rect 53649 646368 336247 646370
rect 53649 646312 53654 646368
rect 53710 646312 336186 646368
rect 336242 646312 336247 646368
rect 53649 646310 336247 646312
rect 53649 646307 53715 646310
rect 336181 646307 336247 646310
rect 52085 646234 52151 646237
rect 334893 646234 334959 646237
rect 52085 646232 334959 646234
rect 52085 646176 52090 646232
rect 52146 646176 334898 646232
rect 334954 646176 334959 646232
rect 52085 646174 334959 646176
rect 52085 646171 52151 646174
rect 334893 646171 334959 646174
rect 53465 646098 53531 646101
rect 345197 646098 345263 646101
rect 53465 646096 345263 646098
rect 53465 646040 53470 646096
rect 53526 646040 345202 646096
rect 345258 646040 345263 646096
rect 53465 646038 345263 646040
rect 53465 646035 53531 646038
rect 345197 646035 345263 646038
rect 36997 645962 37063 645965
rect 351637 645962 351703 645965
rect 36997 645960 351703 645962
rect 36997 645904 37002 645960
rect 37058 645904 351642 645960
rect 351698 645904 351703 645960
rect 36997 645902 351703 645904
rect 36997 645899 37063 645902
rect 351637 645899 351703 645902
rect 542537 645826 542603 645829
rect 539948 645824 542603 645826
rect 539948 645768 542542 645824
rect 542598 645768 542603 645824
rect 539948 645766 542603 645768
rect 542537 645763 542603 645766
rect 35709 645554 35775 645557
rect 106181 645554 106247 645557
rect 35709 645552 106247 645554
rect 35709 645496 35714 645552
rect 35770 645496 106186 645552
rect 106242 645496 106247 645552
rect 35709 645494 106247 645496
rect 35709 645491 35775 645494
rect 106181 645491 106247 645494
rect 216213 645554 216279 645557
rect 227713 645554 227779 645557
rect 216213 645552 227779 645554
rect 216213 645496 216218 645552
rect 216274 645496 227718 645552
rect 227774 645496 227779 645552
rect 216213 645494 227779 645496
rect 216213 645491 216279 645494
rect 227713 645491 227779 645494
rect 102593 645418 102659 645421
rect 278313 645418 278379 645421
rect 102593 645416 278379 645418
rect 102593 645360 102598 645416
rect 102654 645360 278318 645416
rect 278374 645360 278379 645416
rect 102593 645358 278379 645360
rect 102593 645355 102659 645358
rect 278313 645355 278379 645358
rect 98729 645282 98795 645285
rect 275461 645282 275527 645285
rect 98729 645280 275527 645282
rect -960 644996 480 645236
rect 98729 645224 98734 645280
rect 98790 645224 275466 645280
rect 275522 645224 275527 645280
rect 98729 645222 275527 645224
rect 98729 645219 98795 645222
rect 275461 645219 275527 645222
rect 36905 645146 36971 645149
rect 102133 645146 102199 645149
rect 36905 645144 102199 645146
rect 36905 645088 36910 645144
rect 36966 645088 102138 645144
rect 102194 645088 102199 645144
rect 36905 645086 102199 645088
rect 36905 645083 36971 645086
rect 102133 645083 102199 645086
rect 105169 645146 105235 645149
rect 282177 645146 282243 645149
rect 105169 645144 282243 645146
rect 105169 645088 105174 645144
rect 105230 645088 282182 645144
rect 282238 645088 282243 645144
rect 105169 645086 282243 645088
rect 105169 645083 105235 645086
rect 282177 645083 282243 645086
rect 312905 645146 312971 645149
rect 331857 645146 331923 645149
rect 312905 645144 331923 645146
rect 312905 645088 312910 645144
rect 312966 645088 331862 645144
rect 331918 645088 331923 645144
rect 312905 645086 331923 645088
rect 312905 645083 312971 645086
rect 331857 645083 331923 645086
rect 44766 644948 44772 645012
rect 44836 645010 44842 645012
rect 231761 645010 231827 645013
rect 44836 645008 231827 645010
rect 44836 644952 231766 645008
rect 231822 644952 231827 645008
rect 44836 644950 231827 644952
rect 44836 644948 44842 644950
rect 231761 644947 231827 644950
rect 232037 645010 232103 645013
rect 461853 645010 461919 645013
rect 232037 645008 461919 645010
rect 232037 644952 232042 645008
rect 232098 644952 461858 645008
rect 461914 644952 461919 645008
rect 232037 644950 461919 644952
rect 232037 644947 232103 644950
rect 461853 644947 461919 644950
rect 54293 644874 54359 644877
rect 215293 644874 215359 644877
rect 54293 644872 215359 644874
rect 54293 644816 54298 644872
rect 54354 644816 215298 644872
rect 215354 644816 215359 644872
rect 54293 644814 215359 644816
rect 54293 644811 54359 644814
rect 215293 644811 215359 644814
rect 227805 644874 227871 644877
rect 461577 644874 461643 644877
rect 227805 644872 461643 644874
rect 227805 644816 227810 644872
rect 227866 644816 461582 644872
rect 461638 644816 461643 644872
rect 227805 644814 461643 644816
rect 227805 644811 227871 644814
rect 461577 644811 461643 644814
rect 52310 644676 52316 644740
rect 52380 644738 52386 644740
rect 296478 644738 296484 644740
rect 52380 644678 296484 644738
rect 52380 644676 52386 644678
rect 296478 644676 296484 644678
rect 296548 644676 296554 644740
rect 46790 644540 46796 644604
rect 46860 644602 46866 644604
rect 298001 644602 298067 644605
rect 46860 644600 298067 644602
rect 46860 644544 298006 644600
rect 298062 644544 298067 644600
rect 46860 644542 298067 644544
rect 46860 644540 46866 644542
rect 298001 644539 298067 644542
rect 542905 644466 542971 644469
rect 539948 644464 542971 644466
rect 539948 644408 542910 644464
rect 542966 644408 542971 644464
rect 539948 644406 542971 644408
rect 542905 644403 542971 644406
rect 44030 644268 44036 644332
rect 44100 644330 44106 644332
rect 375414 644330 375420 644332
rect 44100 644270 375420 644330
rect 44100 644268 44106 644270
rect 375414 644268 375420 644270
rect 375484 644268 375490 644332
rect 46841 644194 46907 644197
rect 86861 644194 86927 644197
rect 46841 644192 86927 644194
rect 46841 644136 46846 644192
rect 46902 644136 86866 644192
rect 86922 644136 86927 644192
rect 46841 644134 86927 644136
rect 46841 644131 46907 644134
rect 86861 644131 86927 644134
rect 45277 644058 45343 644061
rect 80053 644058 80119 644061
rect 45277 644056 80119 644058
rect 45277 644000 45282 644056
rect 45338 644000 80058 644056
rect 80114 644000 80119 644056
rect 45277 643998 80119 644000
rect 45277 643995 45343 643998
rect 80053 643995 80119 643998
rect 85849 644058 85915 644061
rect 276657 644058 276723 644061
rect 85849 644056 276723 644058
rect 85849 644000 85854 644056
rect 85910 644000 276662 644056
rect 276718 644000 276723 644056
rect 85849 643998 276723 644000
rect 85849 643995 85915 643998
rect 276657 643995 276723 643998
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 88425 643922 88491 643925
rect 287789 643922 287855 643925
rect 88425 643920 287855 643922
rect 88425 643864 88430 643920
rect 88486 643864 287794 643920
rect 287850 643864 287855 643920
rect 583520 643908 584960 643998
rect 88425 643862 287855 643864
rect 88425 643859 88491 643862
rect 287789 643859 287855 643862
rect 80697 643786 80763 643789
rect 291837 643786 291903 643789
rect 80697 643784 291903 643786
rect 80697 643728 80702 643784
rect 80758 643728 291842 643784
rect 291898 643728 291903 643784
rect 80697 643726 291903 643728
rect 80697 643723 80763 643726
rect 291837 643723 291903 643726
rect 31661 643650 31727 643653
rect 176653 643650 176719 643653
rect 31661 643648 176719 643650
rect 31661 643592 31666 643648
rect 31722 643592 176658 643648
rect 176714 643592 176719 643648
rect 31661 643590 176719 643592
rect 31661 643587 31727 643590
rect 176653 643587 176719 643590
rect 177665 643650 177731 643653
rect 204161 643650 204227 643653
rect 177665 643648 204227 643650
rect 177665 643592 177670 643648
rect 177726 643592 204166 643648
rect 204222 643592 204227 643648
rect 177665 643590 204227 643592
rect 177665 643587 177731 643590
rect 204161 643587 204227 643590
rect 207473 643650 207539 643653
rect 233877 643650 233943 643653
rect 207473 643648 233943 643650
rect 207473 643592 207478 643648
rect 207534 643592 233882 643648
rect 233938 643592 233943 643648
rect 207473 643590 233943 643592
rect 207473 643587 207539 643590
rect 233877 643587 233943 643590
rect 234521 643650 234587 643653
rect 472617 643650 472683 643653
rect 234521 643648 472683 643650
rect 234521 643592 234526 643648
rect 234582 643592 472622 643648
rect 472678 643592 472683 643648
rect 234521 643590 472683 643592
rect 234521 643587 234587 643590
rect 472617 643587 472683 643590
rect 46749 643514 46815 643517
rect 297449 643514 297515 643517
rect 46749 643512 297515 643514
rect 46749 643456 46754 643512
rect 46810 643456 297454 643512
rect 297510 643456 297515 643512
rect 46749 643454 297515 643456
rect 46749 643451 46815 643454
rect 297449 643451 297515 643454
rect 52361 643378 52427 643381
rect 303981 643378 304047 643381
rect 52361 643376 304047 643378
rect 52361 643320 52366 643376
rect 52422 643320 303986 643376
rect 304042 643320 304047 643376
rect 52361 643318 304047 643320
rect 52361 643315 52427 643318
rect 303981 643315 304047 643318
rect 45461 643242 45527 643245
rect 88977 643242 89043 643245
rect 179321 643244 179387 643245
rect 179270 643242 179276 643244
rect 45461 643240 89043 643242
rect 45461 643184 45466 643240
rect 45522 643184 88982 643240
rect 89038 643184 89043 643240
rect 45461 643182 89043 643184
rect 179230 643182 179276 643242
rect 179340 643240 179387 643244
rect 179382 643184 179387 643240
rect 45461 643179 45527 643182
rect 88977 643179 89043 643182
rect 179270 643180 179276 643182
rect 179340 643180 179387 643184
rect 179321 643179 179387 643180
rect 203793 643242 203859 643245
rect 207013 643242 207079 643245
rect 203793 643240 207079 643242
rect 203793 643184 203798 643240
rect 203854 643184 207018 643240
rect 207074 643184 207079 643240
rect 203793 643182 207079 643184
rect 203793 643179 203859 643182
rect 207013 643179 207079 643182
rect 542721 643106 542787 643109
rect 539948 643104 542787 643106
rect 539948 643048 542726 643104
rect 542782 643048 542787 643104
rect 539948 643046 542787 643048
rect 542721 643043 542787 643046
rect 53557 642834 53623 642837
rect 223481 642834 223547 642837
rect 53557 642832 223547 642834
rect 53557 642776 53562 642832
rect 53618 642776 223486 642832
rect 223542 642776 223547 642832
rect 53557 642774 223547 642776
rect 53557 642771 53623 642774
rect 223481 642771 223547 642774
rect 42609 642698 42675 642701
rect 376753 642698 376819 642701
rect 42609 642696 376819 642698
rect 42609 642640 42614 642696
rect 42670 642640 376758 642696
rect 376814 642640 376819 642696
rect 42609 642638 376819 642640
rect 42609 642635 42675 642638
rect 376753 642635 376819 642638
rect 54702 642500 54708 642564
rect 54772 642562 54778 642564
rect 92473 642562 92539 642565
rect 54772 642560 92539 642562
rect 54772 642504 92478 642560
rect 92534 642504 92539 642560
rect 54772 642502 92539 642504
rect 54772 642500 54778 642502
rect 92473 642499 92539 642502
rect 93577 642562 93643 642565
rect 278221 642562 278287 642565
rect 93577 642560 278287 642562
rect 93577 642504 93582 642560
rect 93638 642504 278226 642560
rect 278282 642504 278287 642560
rect 93577 642502 278287 642504
rect 93577 642499 93643 642502
rect 278221 642499 278287 642502
rect 84561 642426 84627 642429
rect 279509 642426 279575 642429
rect 84561 642424 279575 642426
rect 84561 642368 84566 642424
rect 84622 642368 279514 642424
rect 279570 642368 279575 642424
rect 84561 642366 279575 642368
rect 84561 642363 84627 642366
rect 279509 642363 279575 642366
rect 48630 642228 48636 642292
rect 48700 642290 48706 642292
rect 296846 642290 296852 642292
rect 48700 642230 296852 642290
rect 48700 642228 48706 642230
rect 296846 642228 296852 642230
rect 296916 642228 296922 642292
rect 46657 642154 46723 642157
rect 297633 642154 297699 642157
rect 46657 642152 297699 642154
rect 46657 642096 46662 642152
rect 46718 642096 297638 642152
rect 297694 642096 297699 642152
rect 46657 642094 297699 642096
rect 46657 642091 46723 642094
rect 297633 642091 297699 642094
rect 50981 642018 51047 642021
rect 309133 642018 309199 642021
rect 50981 642016 309199 642018
rect 50981 641960 50986 642016
rect 51042 641960 309138 642016
rect 309194 641960 309199 642016
rect 50981 641958 309199 641960
rect 50981 641955 51047 641958
rect 309133 641955 309199 641958
rect 222929 641882 222995 641885
rect 488993 641882 489059 641885
rect 222929 641880 489059 641882
rect 222929 641824 222934 641880
rect 222990 641824 488998 641880
rect 489054 641824 489059 641880
rect 222929 641822 489059 641824
rect 222929 641819 222995 641822
rect 488993 641819 489059 641822
rect 35617 641746 35683 641749
rect 85481 641746 85547 641749
rect 35617 641744 85547 641746
rect 35617 641688 35622 641744
rect 35678 641688 85486 641744
rect 85542 641688 85547 641744
rect 35617 641686 85547 641688
rect 35617 641683 35683 641686
rect 85481 641683 85547 641686
rect 177246 641684 177252 641748
rect 177316 641746 177322 641748
rect 177941 641746 178007 641749
rect 177316 641744 178007 641746
rect 177316 641688 177946 641744
rect 178002 641688 178007 641744
rect 177316 641686 178007 641688
rect 177316 641684 177322 641686
rect 177941 641683 178007 641686
rect 179086 641684 179092 641748
rect 179156 641746 179162 641748
rect 179321 641746 179387 641749
rect 179156 641744 179387 641746
rect 179156 641688 179326 641744
rect 179382 641688 179387 641744
rect 179156 641686 179387 641688
rect 179156 641684 179162 641686
rect 179321 641683 179387 641686
rect 488533 641746 488599 641749
rect 489494 641746 489500 641748
rect 488533 641744 489500 641746
rect 488533 641688 488538 641744
rect 488594 641688 489500 641744
rect 488533 641686 489500 641688
rect 488533 641683 488599 641686
rect 489494 641684 489500 641686
rect 489564 641684 489570 641748
rect 541157 641746 541223 641749
rect 539948 641744 541223 641746
rect 539948 641688 541162 641744
rect 541218 641688 541223 641744
rect 539948 641686 541223 641688
rect 541157 641683 541223 641686
rect 42701 641474 42767 641477
rect 218053 641474 218119 641477
rect 42701 641472 218119 641474
rect 42701 641416 42706 641472
rect 42762 641416 218058 641472
rect 218114 641416 218119 641472
rect 42701 641414 218119 641416
rect 42701 641411 42767 641414
rect 218053 641411 218119 641414
rect 36813 641338 36879 641341
rect 376937 641338 377003 641341
rect 36813 641336 377003 641338
rect 36813 641280 36818 641336
rect 36874 641280 376942 641336
rect 376998 641280 377003 641336
rect 36813 641278 377003 641280
rect 36813 641275 36879 641278
rect 376937 641275 377003 641278
rect 51993 641202 52059 641205
rect 91093 641202 91159 641205
rect 51993 641200 91159 641202
rect 51993 641144 51998 641200
rect 52054 641144 91098 641200
rect 91154 641144 91159 641200
rect 51993 641142 91159 641144
rect 51993 641139 52059 641142
rect 91093 641139 91159 641142
rect 92289 641202 92355 641205
rect 276749 641202 276815 641205
rect 92289 641200 276815 641202
rect 92289 641144 92294 641200
rect 92350 641144 276754 641200
rect 276810 641144 276815 641200
rect 92289 641142 276815 641144
rect 92289 641139 92355 641142
rect 276749 641139 276815 641142
rect 487654 641140 487660 641204
rect 487724 641202 487730 641204
rect 487724 641142 490084 641202
rect 487724 641140 487730 641142
rect 50838 641004 50844 641068
rect 50908 641066 50914 641068
rect 297357 641066 297423 641069
rect 50908 641064 297423 641066
rect 50908 641008 297362 641064
rect 297418 641008 297423 641064
rect 50908 641006 297423 641008
rect 50908 641004 50914 641006
rect 297357 641003 297423 641006
rect 52269 640930 52335 640933
rect 305269 640930 305335 640933
rect 52269 640928 305335 640930
rect 52269 640872 52274 640928
rect 52330 640872 305274 640928
rect 305330 640872 305335 640928
rect 52269 640870 305335 640872
rect 52269 640867 52335 640870
rect 305269 640867 305335 640870
rect 45369 640794 45435 640797
rect 56501 640794 56567 640797
rect 45369 640792 56567 640794
rect 45369 640736 45374 640792
rect 45430 640736 56506 640792
rect 56562 640736 56567 640792
rect 45369 640734 56567 640736
rect 45369 640731 45435 640734
rect 56501 640731 56567 640734
rect 217961 640794 218027 640797
rect 230381 640794 230447 640797
rect 217961 640792 230447 640794
rect 217961 640736 217966 640792
rect 218022 640736 230386 640792
rect 230442 640736 230447 640792
rect 217961 640734 230447 640736
rect 217961 640731 218027 640734
rect 230381 640731 230447 640734
rect 230657 640794 230723 640797
rect 485957 640794 486023 640797
rect 230657 640792 486023 640794
rect 230657 640736 230662 640792
rect 230718 640736 485962 640792
rect 486018 640736 486023 640792
rect 230657 640734 486023 640736
rect 230657 640731 230723 640734
rect 485957 640731 486023 640734
rect 219065 640658 219131 640661
rect 487521 640658 487587 640661
rect 219065 640656 487587 640658
rect 219065 640600 219070 640656
rect 219126 640600 487526 640656
rect 487582 640600 487587 640656
rect 219065 640598 487587 640600
rect 219065 640595 219131 640598
rect 487521 640595 487587 640598
rect 37089 640522 37155 640525
rect 310421 640522 310487 640525
rect 37089 640520 310487 640522
rect 37089 640464 37094 640520
rect 37150 640464 310426 640520
rect 310482 640464 310487 640520
rect 37089 640462 310487 640464
rect 37089 640459 37155 640462
rect 310421 640459 310487 640462
rect 55806 640324 55812 640388
rect 55876 640386 55882 640388
rect 214557 640386 214623 640389
rect 55876 640384 214623 640386
rect 55876 640328 214562 640384
rect 214618 640328 214623 640384
rect 55876 640326 214623 640328
rect 55876 640324 55882 640326
rect 214557 640323 214623 640326
rect 215201 640386 215267 640389
rect 216765 640386 216831 640389
rect 541065 640386 541131 640389
rect 215201 640384 216831 640386
rect 215201 640328 215206 640384
rect 215262 640328 216770 640384
rect 216826 640328 216831 640384
rect 215201 640326 216831 640328
rect 539948 640384 541131 640386
rect 539948 640328 541070 640384
rect 541126 640328 541131 640384
rect 539948 640326 541131 640328
rect 215201 640323 215267 640326
rect 216765 640323 216831 640326
rect 541065 640323 541131 640326
rect 41270 640052 41276 640116
rect 41340 640114 41346 640116
rect 125593 640114 125659 640117
rect 41340 640112 125659 640114
rect 41340 640056 125598 640112
rect 125654 640056 125659 640112
rect 41340 640054 125659 640056
rect 41340 640052 41346 640054
rect 125593 640051 125659 640054
rect 199745 640114 199811 640117
rect 251081 640114 251147 640117
rect 199745 640112 251147 640114
rect 199745 640056 199750 640112
rect 199806 640056 251086 640112
rect 251142 640056 251147 640112
rect 199745 640054 251147 640056
rect 199745 640051 199811 640054
rect 251081 640051 251147 640054
rect 41321 639978 41387 639981
rect 82813 639978 82879 639981
rect 41321 639976 82879 639978
rect 41321 639920 41326 639976
rect 41382 639920 82818 639976
rect 82874 639920 82879 639976
rect 41321 639918 82879 639920
rect 41321 639915 41387 639918
rect 82813 639915 82879 639918
rect 94865 639978 94931 639981
rect 206369 639978 206435 639981
rect 488717 639978 488783 639981
rect 94865 639976 103530 639978
rect 94865 639920 94870 639976
rect 94926 639920 103530 639976
rect 94865 639918 103530 639920
rect 94865 639915 94931 639918
rect 58934 639780 58940 639844
rect 59004 639842 59010 639844
rect 95141 639842 95207 639845
rect 59004 639840 95207 639842
rect 59004 639784 95146 639840
rect 95202 639784 95207 639840
rect 59004 639782 95207 639784
rect 103470 639842 103530 639918
rect 206369 639976 488783 639978
rect 206369 639920 206374 639976
rect 206430 639920 488722 639976
rect 488778 639920 488783 639976
rect 206369 639918 488783 639920
rect 206369 639915 206435 639918
rect 488717 639915 488783 639918
rect 152549 639842 152615 639845
rect 103470 639840 152615 639842
rect 103470 639784 152554 639840
rect 152610 639784 152615 639840
rect 103470 639782 152615 639784
rect 59004 639780 59010 639782
rect 95141 639779 95207 639782
rect 152549 639779 152615 639782
rect 250989 639842 251055 639845
rect 358721 639842 358787 639845
rect 250989 639840 358787 639842
rect 250989 639784 250994 639840
rect 251050 639784 358726 639840
rect 358782 639784 358787 639840
rect 250989 639782 358787 639784
rect 250989 639779 251055 639782
rect 358721 639779 358787 639782
rect 67817 639706 67883 639709
rect 287697 639706 287763 639709
rect 67817 639704 287763 639706
rect 67817 639648 67822 639704
rect 67878 639648 287702 639704
rect 287758 639648 287763 639704
rect 67817 639646 287763 639648
rect 67817 639643 67883 639646
rect 287697 639643 287763 639646
rect 121913 639570 121979 639573
rect 140773 639570 140839 639573
rect 121913 639568 140839 639570
rect 121913 639512 121918 639568
rect 121974 639512 140778 639568
rect 140834 639512 140839 639568
rect 121913 639510 140839 639512
rect 121913 639507 121979 639510
rect 140773 639507 140839 639510
rect 198641 639570 198707 639573
rect 234613 639570 234679 639573
rect 198641 639568 234679 639570
rect 198641 639512 198646 639568
rect 198702 639512 234618 639568
rect 234674 639512 234679 639568
rect 198641 639510 234679 639512
rect 198641 639507 198707 639510
rect 234613 639507 234679 639510
rect 235901 639570 235967 639573
rect 462957 639570 463023 639573
rect 235901 639568 463023 639570
rect 235901 639512 235906 639568
rect 235962 639512 462962 639568
rect 463018 639512 463023 639568
rect 235901 639510 463023 639512
rect 235901 639507 235967 639510
rect 462957 639507 463023 639510
rect 46473 639434 46539 639437
rect 297725 639434 297791 639437
rect 46473 639432 297791 639434
rect 46473 639376 46478 639432
rect 46534 639376 297730 639432
rect 297786 639376 297791 639432
rect 46473 639374 297791 639376
rect 46473 639371 46539 639374
rect 297725 639371 297791 639374
rect 55029 639298 55095 639301
rect 81433 639298 81499 639301
rect 55029 639296 81499 639298
rect 55029 639240 55034 639296
rect 55090 639240 81438 639296
rect 81494 639240 81499 639296
rect 55029 639238 81499 639240
rect 55029 639235 55095 639238
rect 81433 639235 81499 639238
rect 83273 639298 83339 639301
rect 155309 639298 155375 639301
rect 83273 639296 155375 639298
rect 83273 639240 83278 639296
rect 83334 639240 155314 639296
rect 155370 639240 155375 639296
rect 83273 639238 155375 639240
rect 83273 639235 83339 639238
rect 155309 639235 155375 639238
rect 213821 639298 213887 639301
rect 220353 639298 220419 639301
rect 479241 639298 479307 639301
rect 213821 639296 219450 639298
rect 213821 639240 213826 639296
rect 213882 639240 219450 639296
rect 213821 639238 219450 639240
rect 213821 639235 213887 639238
rect 81985 639162 82051 639165
rect 155493 639162 155559 639165
rect 81985 639160 155559 639162
rect 81985 639104 81990 639160
rect 82046 639104 155498 639160
rect 155554 639104 155559 639160
rect 81985 639102 155559 639104
rect 81985 639099 82051 639102
rect 155493 639099 155559 639102
rect 184289 639162 184355 639165
rect 213821 639162 213887 639165
rect 184289 639160 213887 639162
rect 184289 639104 184294 639160
rect 184350 639104 213826 639160
rect 213882 639104 213887 639160
rect 184289 639102 213887 639104
rect 219390 639162 219450 639238
rect 220353 639296 479307 639298
rect 220353 639240 220358 639296
rect 220414 639240 479246 639296
rect 479302 639240 479307 639296
rect 220353 639238 479307 639240
rect 220353 639235 220419 639238
rect 479241 639235 479307 639238
rect 488901 639162 488967 639165
rect 219390 639160 488967 639162
rect 219390 639104 488906 639160
rect 488962 639104 488967 639160
rect 219390 639102 488967 639104
rect 184289 639099 184355 639102
rect 213821 639099 213887 639102
rect 488901 639099 488967 639102
rect 50889 639026 50955 639029
rect 122741 639026 122807 639029
rect 50889 639024 122807 639026
rect 50889 638968 50894 639024
rect 50950 638968 122746 639024
rect 122802 638968 122807 639024
rect 50889 638966 122807 638968
rect 50889 638963 50955 638966
rect 122741 638963 122807 638966
rect 125777 639026 125843 639029
rect 138105 639026 138171 639029
rect 125777 639024 138171 639026
rect 125777 638968 125782 639024
rect 125838 638968 138110 639024
rect 138166 638968 138171 639024
rect 125777 638966 138171 638968
rect 125777 638963 125843 638966
rect 138105 638963 138171 638966
rect 197261 639026 197327 639029
rect 220721 639026 220787 639029
rect 197261 639024 220787 639026
rect 197261 638968 197266 639024
rect 197322 638968 220726 639024
rect 220782 638968 220787 639024
rect 197261 638966 220787 638968
rect 197261 638963 197327 638966
rect 220721 638963 220787 638966
rect 485773 639026 485839 639029
rect 486182 639026 486188 639028
rect 485773 639024 486188 639026
rect 485773 638968 485778 639024
rect 485834 638968 486188 639024
rect 485773 638966 486188 638968
rect 485773 638963 485839 638966
rect 486182 638964 486188 638966
rect 486252 638964 486258 639028
rect 540973 639026 541039 639029
rect 539948 639024 541039 639026
rect 539948 638968 540978 639024
rect 541034 638968 541039 639024
rect 539948 638966 541039 638968
rect 540973 638963 541039 638966
rect 39798 638692 39804 638756
rect 39868 638754 39874 638756
rect 109033 638754 109099 638757
rect 39868 638752 109099 638754
rect 39868 638696 109038 638752
rect 109094 638696 109099 638752
rect 39868 638694 109099 638696
rect 39868 638692 39874 638694
rect 109033 638691 109099 638694
rect 87137 638618 87203 638621
rect 155401 638618 155467 638621
rect 87137 638616 155467 638618
rect 87137 638560 87142 638616
rect 87198 638560 155406 638616
rect 155462 638560 155467 638616
rect 87137 638558 155467 638560
rect 87137 638555 87203 638558
rect 155401 638555 155467 638558
rect 210141 638618 210207 638621
rect 230381 638618 230447 638621
rect 210141 638616 230447 638618
rect 210141 638560 210146 638616
rect 210202 638560 230386 638616
rect 230442 638560 230447 638616
rect 210141 638558 230447 638560
rect 210141 638555 210207 638558
rect 230381 638555 230447 638558
rect 107745 638482 107811 638485
rect 129733 638482 129799 638485
rect 107745 638480 129799 638482
rect 107745 638424 107750 638480
rect 107806 638424 129738 638480
rect 129794 638424 129799 638480
rect 107745 638422 129799 638424
rect 107745 638419 107811 638422
rect 129733 638419 129799 638422
rect 130929 638482 130995 638485
rect 250989 638482 251055 638485
rect 130929 638480 251055 638482
rect 130929 638424 130934 638480
rect 130990 638424 250994 638480
rect 251050 638424 251055 638480
rect 130929 638422 251055 638424
rect 130929 638419 130995 638422
rect 250989 638419 251055 638422
rect 89713 638346 89779 638349
rect 279601 638346 279667 638349
rect 89713 638344 279667 638346
rect 89713 638288 89718 638344
rect 89774 638288 279606 638344
rect 279662 638288 279667 638344
rect 89713 638286 279667 638288
rect 89713 638283 89779 638286
rect 279601 638283 279667 638286
rect 76833 638210 76899 638213
rect 279417 638210 279483 638213
rect 76833 638208 279483 638210
rect 76833 638152 76838 638208
rect 76894 638152 279422 638208
rect 279478 638152 279483 638208
rect 76833 638150 279483 638152
rect 76833 638147 76899 638150
rect 279417 638147 279483 638150
rect 69105 638074 69171 638077
rect 278037 638074 278103 638077
rect 69105 638072 278103 638074
rect 69105 638016 69110 638072
rect 69166 638016 278042 638072
rect 278098 638016 278103 638072
rect 69105 638014 278103 638016
rect 69105 638011 69171 638014
rect 278037 638011 278103 638014
rect 66529 637938 66595 637941
rect 294597 637938 294663 637941
rect 66529 637936 294663 637938
rect 66529 637880 66534 637936
rect 66590 637880 294602 637936
rect 294658 637880 294663 637936
rect 66529 637878 294663 637880
rect 66529 637875 66595 637878
rect 294597 637875 294663 637878
rect 39849 637802 39915 637805
rect 108297 637802 108363 637805
rect 39849 637800 108363 637802
rect 39849 637744 39854 637800
rect 39910 637744 108302 637800
rect 108358 637744 108363 637800
rect 39849 637742 108363 637744
rect 39849 637739 39915 637742
rect 108297 637739 108363 637742
rect 123201 637802 123267 637805
rect 139393 637802 139459 637805
rect 123201 637800 139459 637802
rect 123201 637744 123206 637800
rect 123262 637744 139398 637800
rect 139454 637744 139459 637800
rect 123201 637742 139459 637744
rect 123201 637739 123267 637742
rect 139393 637739 139459 637742
rect 183185 637802 183251 637805
rect 211061 637802 211127 637805
rect 183185 637800 211127 637802
rect 183185 637744 183190 637800
rect 183246 637744 211066 637800
rect 211122 637744 211127 637800
rect 183185 637742 211127 637744
rect 183185 637739 183251 637742
rect 211061 637739 211127 637742
rect 224309 637802 224375 637805
rect 471513 637802 471579 637805
rect 224309 637800 471579 637802
rect 224309 637744 224314 637800
rect 224370 637744 471518 637800
rect 471574 637744 471579 637800
rect 224309 637742 471579 637744
rect 224309 637739 224375 637742
rect 471513 637739 471579 637742
rect 109493 637666 109559 637669
rect 123477 637666 123543 637669
rect 109493 637664 123543 637666
rect 109493 637608 109498 637664
rect 109554 637608 123482 637664
rect 123538 637608 123543 637664
rect 109493 637606 123543 637608
rect 109493 637603 109559 637606
rect 123477 637603 123543 637606
rect 195881 637666 195947 637669
rect 224217 637666 224283 637669
rect 195881 637664 224283 637666
rect 195881 637608 195886 637664
rect 195942 637608 224222 637664
rect 224278 637608 224283 637664
rect 195881 637606 224283 637608
rect 195881 637603 195947 637606
rect 224217 637603 224283 637606
rect 229553 637666 229619 637669
rect 479977 637666 480043 637669
rect 487153 637668 487219 637669
rect 229553 637664 480043 637666
rect 229553 637608 229558 637664
rect 229614 637608 479982 637664
rect 480038 637608 480043 637664
rect 229553 637606 480043 637608
rect 229553 637603 229619 637606
rect 479977 637603 480043 637606
rect 487102 637604 487108 637668
rect 487172 637666 487219 637668
rect 488533 637666 488599 637669
rect 489310 637666 489316 637668
rect 487172 637664 487264 637666
rect 487214 637608 487264 637664
rect 487172 637606 487264 637608
rect 488533 637664 489316 637666
rect 488533 637608 488538 637664
rect 488594 637608 489316 637664
rect 488533 637606 489316 637608
rect 487172 637604 487219 637606
rect 487153 637603 487219 637604
rect 488533 637603 488599 637606
rect 489310 637604 489316 637606
rect 489380 637604 489386 637668
rect 541249 637666 541315 637669
rect 539948 637664 541315 637666
rect 539948 637608 541254 637664
rect 541310 637608 541315 637664
rect 539948 637606 541315 637608
rect 541249 637603 541315 637606
rect 58750 637468 58756 637532
rect 58820 637530 58826 637532
rect 99373 637530 99439 637533
rect 58820 637528 99439 637530
rect 58820 637472 99378 637528
rect 99434 637472 99439 637528
rect 58820 637470 99439 637472
rect 58820 637468 58826 637470
rect 99373 637467 99439 637470
rect 71681 637394 71747 637397
rect 136081 637394 136147 637397
rect 71681 637392 136147 637394
rect 71681 637336 71686 637392
rect 71742 637336 136086 637392
rect 136142 637336 136147 637392
rect 71681 637334 136147 637336
rect 71681 637331 71747 637334
rect 136081 637331 136147 637334
rect 63953 637258 64019 637261
rect 152457 637258 152523 637261
rect 63953 637256 152523 637258
rect 63953 637200 63958 637256
rect 64014 637200 152462 637256
rect 152518 637200 152523 637256
rect 63953 637198 152523 637200
rect 63953 637195 64019 637198
rect 152457 637195 152523 637198
rect 245009 637258 245075 637261
rect 249609 637258 249675 637261
rect 245009 637256 249675 637258
rect 245009 637200 245014 637256
rect 245070 637200 249614 637256
rect 249670 637200 249675 637256
rect 245009 637198 249675 637200
rect 245009 637195 245075 637198
rect 249609 637195 249675 637198
rect 100017 637122 100083 637125
rect 124213 637122 124279 637125
rect 100017 637120 124279 637122
rect 100017 637064 100022 637120
rect 100078 637064 124218 637120
rect 124274 637064 124279 637120
rect 100017 637062 124279 637064
rect 100017 637059 100083 637062
rect 124213 637059 124279 637062
rect 177573 637122 177639 637125
rect 485814 637122 485820 637124
rect 177573 637120 485820 637122
rect 177573 637064 177578 637120
rect 177634 637064 485820 637120
rect 177573 637062 485820 637064
rect 177573 637059 177639 637062
rect 485814 637060 485820 637062
rect 485884 637060 485890 637124
rect 75545 636986 75611 636989
rect 78121 636986 78187 636989
rect 131113 636986 131179 636989
rect 75545 636984 76114 636986
rect 75545 636928 75550 636984
rect 75606 636928 76114 636984
rect 75545 636926 76114 636928
rect 75545 636923 75611 636926
rect 58566 636788 58572 636852
rect 58636 636850 58642 636852
rect 75821 636850 75887 636853
rect 58636 636848 75887 636850
rect 58636 636792 75826 636848
rect 75882 636792 75887 636848
rect 58636 636790 75887 636792
rect 76054 636850 76114 636926
rect 78121 636984 131179 636986
rect 78121 636928 78126 636984
rect 78182 636928 131118 636984
rect 131174 636928 131179 636984
rect 78121 636926 131179 636928
rect 78121 636923 78187 636926
rect 131113 636923 131179 636926
rect 178902 636924 178908 636988
rect 178972 636986 178978 636988
rect 282862 636986 282868 636988
rect 178972 636926 282868 636986
rect 178972 636924 178978 636926
rect 282862 636924 282868 636926
rect 282932 636924 282938 636988
rect 134609 636850 134675 636853
rect 76054 636848 134675 636850
rect 76054 636792 134614 636848
rect 134670 636792 134675 636848
rect 76054 636790 134675 636792
rect 58636 636788 58642 636790
rect 75821 636787 75887 636790
rect 134609 636787 134675 636790
rect 176561 636850 176627 636853
rect 295057 636850 295123 636853
rect 176561 636848 295123 636850
rect 176561 636792 176566 636848
rect 176622 636792 295062 636848
rect 295118 636792 295123 636848
rect 176561 636790 295123 636792
rect 176561 636787 176627 636790
rect 295057 636787 295123 636790
rect 358721 636850 358787 636853
rect 370957 636850 371023 636853
rect 358721 636848 371023 636850
rect 358721 636792 358726 636848
rect 358782 636792 370962 636848
rect 371018 636792 371023 636848
rect 358721 636790 371023 636792
rect 358721 636787 358787 636790
rect 370957 636787 371023 636790
rect 62665 636714 62731 636717
rect 254577 636714 254643 636717
rect 62665 636712 254643 636714
rect 62665 636656 62670 636712
rect 62726 636656 254582 636712
rect 254638 636656 254643 636712
rect 62665 636654 254643 636656
rect 62665 636651 62731 636654
rect 254577 636651 254643 636654
rect 52126 636516 52132 636580
rect 52196 636578 52202 636580
rect 73153 636578 73219 636581
rect 52196 636576 73219 636578
rect 52196 636520 73158 636576
rect 73214 636520 73219 636576
rect 52196 636518 73219 636520
rect 52196 636516 52202 636518
rect 73153 636515 73219 636518
rect 132217 636578 132283 636581
rect 163589 636578 163655 636581
rect 132217 636576 163655 636578
rect 132217 636520 132222 636576
rect 132278 636520 163594 636576
rect 163650 636520 163655 636576
rect 132217 636518 163655 636520
rect 132217 636515 132283 636518
rect 163589 636515 163655 636518
rect 221825 636578 221891 636581
rect 464613 636578 464679 636581
rect 221825 636576 464679 636578
rect 221825 636520 221830 636576
rect 221886 636520 464618 636576
rect 464674 636520 464679 636576
rect 221825 636518 464679 636520
rect 221825 636515 221891 636518
rect 464613 636515 464679 636518
rect 74257 636442 74323 636445
rect 159449 636442 159515 636445
rect 74257 636440 159515 636442
rect 74257 636384 74262 636440
rect 74318 636384 159454 636440
rect 159510 636384 159515 636440
rect 74257 636382 159515 636384
rect 74257 636379 74323 636382
rect 159449 636379 159515 636382
rect 177614 636380 177620 636444
rect 177684 636442 177690 636444
rect 479374 636442 479380 636444
rect 177684 636382 479380 636442
rect 177684 636380 177690 636382
rect 479374 636380 479380 636382
rect 479444 636380 479450 636444
rect 53281 636306 53347 636309
rect 78581 636306 78647 636309
rect 53281 636304 78647 636306
rect 53281 636248 53286 636304
rect 53342 636248 78586 636304
rect 78642 636248 78647 636304
rect 53281 636246 78647 636248
rect 53281 636243 53347 636246
rect 78581 636243 78647 636246
rect 124489 636306 124555 636309
rect 135253 636306 135319 636309
rect 124489 636304 135319 636306
rect 124489 636248 124494 636304
rect 124550 636248 135258 636304
rect 135314 636248 135319 636304
rect 124489 636246 135319 636248
rect 124489 636243 124555 636246
rect 135253 636243 135319 636246
rect 225689 636306 225755 636309
rect 248781 636306 248847 636309
rect 262857 636306 262923 636309
rect 541014 636306 541020 636308
rect 225689 636304 244290 636306
rect 225689 636248 225694 636304
rect 225750 636248 244290 636304
rect 225689 636246 244290 636248
rect 225689 636243 225755 636246
rect 244230 636170 244290 636246
rect 248781 636304 262923 636306
rect 248781 636248 248786 636304
rect 248842 636248 262862 636304
rect 262918 636248 262923 636304
rect 248781 636246 262923 636248
rect 539948 636246 541020 636306
rect 248781 636243 248847 636246
rect 262857 636243 262923 636246
rect 541014 636244 541020 636246
rect 541084 636244 541090 636308
rect 252461 636170 252527 636173
rect 244230 636168 252527 636170
rect 244230 636112 252466 636168
rect 252522 636112 252527 636168
rect 244230 636110 252527 636112
rect 252461 636107 252527 636110
rect 331857 636170 331923 636173
rect 335169 636170 335235 636173
rect 331857 636168 335235 636170
rect 331857 636112 331862 636168
rect 331918 636112 335174 636168
rect 335230 636112 335235 636168
rect 331857 636110 335235 636112
rect 331857 636107 331923 636110
rect 335169 636107 335235 636110
rect 54845 636034 54911 636037
rect 140037 636034 140103 636037
rect 54845 636032 140103 636034
rect 54845 635976 54850 636032
rect 54906 635976 140042 636032
rect 140098 635976 140103 636032
rect 54845 635974 140103 635976
rect 54845 635971 54911 635974
rect 140037 635971 140103 635974
rect 70393 635898 70459 635901
rect 256141 635898 256207 635901
rect 70393 635896 256207 635898
rect 70393 635840 70398 635896
rect 70454 635840 256146 635896
rect 256202 635840 256207 635896
rect 70393 635838 256207 635840
rect 70393 635835 70459 635838
rect 256141 635835 256207 635838
rect 43989 635762 44055 635765
rect 70577 635762 70643 635765
rect 43989 635760 70643 635762
rect 43989 635704 43994 635760
rect 44050 635704 70582 635760
rect 70638 635704 70643 635760
rect 43989 635702 70643 635704
rect 43989 635699 44055 635702
rect 70577 635699 70643 635702
rect 79409 635762 79475 635765
rect 121361 635762 121427 635765
rect 79409 635760 121427 635762
rect 79409 635704 79414 635760
rect 79470 635704 121366 635760
rect 121422 635704 121427 635760
rect 79409 635702 121427 635704
rect 79409 635699 79475 635702
rect 121361 635699 121427 635702
rect 201125 635762 201191 635765
rect 244273 635762 244339 635765
rect 201125 635760 244339 635762
rect 201125 635704 201130 635760
rect 201186 635704 244278 635760
rect 244334 635704 244339 635760
rect 201125 635702 244339 635704
rect 201125 635699 201191 635702
rect 244273 635699 244339 635702
rect 48446 635564 48452 635628
rect 48516 635626 48522 635628
rect 97901 635626 97967 635629
rect 48516 635624 97967 635626
rect 48516 635568 97906 635624
rect 97962 635568 97967 635624
rect 48516 635566 97967 635568
rect 48516 635564 48522 635566
rect 97901 635563 97967 635566
rect 98085 635626 98151 635629
rect 119981 635626 120047 635629
rect 98085 635624 120047 635626
rect 98085 635568 98090 635624
rect 98146 635568 119986 635624
rect 120042 635568 120047 635624
rect 98085 635566 120047 635568
rect 98085 635563 98151 635566
rect 119981 635563 120047 635566
rect 179045 635626 179111 635629
rect 291929 635626 291995 635629
rect 179045 635624 291995 635626
rect 179045 635568 179050 635624
rect 179106 635568 291934 635624
rect 291990 635568 291995 635624
rect 179045 635566 291995 635568
rect 179045 635563 179111 635566
rect 291929 635563 291995 635566
rect 54937 635490 55003 635493
rect 136909 635490 136975 635493
rect 54937 635488 136975 635490
rect 54937 635432 54942 635488
rect 54998 635432 136914 635488
rect 136970 635432 136975 635488
rect 54937 635430 136975 635432
rect 54937 635427 55003 635430
rect 136909 635427 136975 635430
rect 179229 635490 179295 635493
rect 294689 635490 294755 635493
rect 179229 635488 294755 635490
rect 179229 635432 179234 635488
rect 179290 635432 294694 635488
rect 294750 635432 294755 635488
rect 179229 635430 294755 635432
rect 179229 635427 179295 635430
rect 294689 635427 294755 635430
rect 46565 635354 46631 635357
rect 53833 635354 53899 635357
rect 46565 635352 53899 635354
rect 46565 635296 46570 635352
rect 46626 635296 53838 635352
rect 53894 635296 53899 635352
rect 46565 635294 53899 635296
rect 46565 635291 46631 635294
rect 53833 635291 53899 635294
rect 54661 635354 54727 635357
rect 138841 635354 138907 635357
rect 54661 635352 138907 635354
rect 54661 635296 54666 635352
rect 54722 635296 138846 635352
rect 138902 635296 138907 635352
rect 54661 635294 138907 635296
rect 54661 635291 54727 635294
rect 138841 635291 138907 635294
rect 179321 635354 179387 635357
rect 294873 635354 294939 635357
rect 179321 635352 294939 635354
rect 179321 635296 179326 635352
rect 179382 635296 294878 635352
rect 294934 635296 294939 635352
rect 179321 635294 294939 635296
rect 179321 635291 179387 635294
rect 294873 635291 294939 635294
rect 44950 635156 44956 635220
rect 45020 635218 45026 635220
rect 71865 635218 71931 635221
rect 45020 635216 71931 635218
rect 45020 635160 71870 635216
rect 71926 635160 71931 635216
rect 45020 635158 71931 635160
rect 45020 635156 45026 635158
rect 71865 635155 71931 635158
rect 72969 635218 73035 635221
rect 255957 635218 256023 635221
rect 72969 635216 256023 635218
rect 72969 635160 72974 635216
rect 73030 635160 255962 635216
rect 256018 635160 256023 635216
rect 72969 635158 256023 635160
rect 72969 635155 73035 635158
rect 255957 635155 256023 635158
rect 48221 635082 48287 635085
rect 79317 635082 79383 635085
rect 48221 635080 79383 635082
rect 48221 635024 48226 635080
rect 48282 635024 79322 635080
rect 79378 635024 79383 635080
rect 48221 635022 79383 635024
rect 48221 635019 48287 635022
rect 79317 635019 79383 635022
rect 121085 635082 121151 635085
rect 136633 635082 136699 635085
rect 121085 635080 136699 635082
rect 121085 635024 121090 635080
rect 121146 635024 136638 635080
rect 136694 635024 136699 635080
rect 121085 635022 136699 635024
rect 121085 635019 121151 635022
rect 136633 635019 136699 635022
rect 177798 635020 177804 635084
rect 177868 635082 177874 635084
rect 226333 635082 226399 635085
rect 177868 635080 226399 635082
rect 177868 635024 226338 635080
rect 226394 635024 226399 635080
rect 177868 635022 226399 635024
rect 177868 635020 177874 635022
rect 226333 635019 226399 635022
rect 252461 635082 252527 635085
rect 471421 635082 471487 635085
rect 252461 635080 471487 635082
rect 252461 635024 252466 635080
rect 252522 635024 471426 635080
rect 471482 635024 471487 635080
rect 252461 635022 471487 635024
rect 252461 635019 252527 635022
rect 471421 635019 471487 635022
rect 119337 634946 119403 634949
rect 135345 634946 135411 634949
rect 119337 634944 135411 634946
rect 119337 634888 119342 634944
rect 119398 634888 135350 634944
rect 135406 634888 135411 634944
rect 119337 634886 135411 634888
rect 119337 634883 119403 634886
rect 135345 634883 135411 634886
rect 226471 634946 226537 634949
rect 464521 634946 464587 634949
rect 541341 634946 541407 634949
rect 226471 634944 464587 634946
rect 226471 634888 226476 634944
rect 226532 634888 464526 634944
rect 464582 634888 464587 634944
rect 226471 634886 464587 634888
rect 539948 634944 541407 634946
rect 539948 634888 541346 634944
rect 541402 634888 541407 634944
rect 539948 634886 541407 634888
rect 226471 634883 226537 634886
rect 464521 634883 464587 634886
rect 541341 634883 541407 634886
rect 48078 634748 48084 634812
rect 48148 634810 48154 634812
rect 296478 634810 296484 634812
rect 48148 634750 296484 634810
rect 48148 634748 48154 634750
rect 296478 634748 296484 634750
rect 296548 634748 296554 634812
rect 296662 634748 296668 634812
rect 296732 634810 296738 634812
rect 297909 634810 297975 634813
rect 296732 634808 297975 634810
rect 296732 634752 297914 634808
rect 297970 634752 297975 634808
rect 296732 634750 297975 634752
rect 296732 634748 296738 634750
rect 297909 634747 297975 634750
rect 127065 634674 127131 634677
rect 140865 634674 140931 634677
rect 127065 634672 140931 634674
rect 127065 634616 127070 634672
rect 127126 634616 140870 634672
rect 140926 634616 140931 634672
rect 127065 634614 140931 634616
rect 127065 634611 127131 634614
rect 140865 634611 140931 634614
rect 177941 634674 178007 634677
rect 484342 634674 484348 634676
rect 177941 634672 484348 634674
rect 177941 634616 177946 634672
rect 178002 634616 484348 634672
rect 177941 634614 484348 634616
rect 177941 634611 178007 634614
rect 484342 634612 484348 634614
rect 484412 634612 484418 634676
rect 48129 634538 48195 634541
rect 129825 634538 129891 634541
rect 48129 634536 129891 634538
rect 48129 634480 48134 634536
rect 48190 634480 129830 634536
rect 129886 634480 129891 634536
rect 48129 634478 129891 634480
rect 48129 634475 48195 634478
rect 129825 634475 129891 634478
rect 130929 634538 130995 634541
rect 140957 634538 141023 634541
rect 130929 634536 141023 634538
rect 130929 634480 130934 634536
rect 130990 634480 140962 634536
rect 141018 634480 141023 634536
rect 130929 634478 141023 634480
rect 130929 634475 130995 634478
rect 140957 634475 141023 634478
rect 179137 634538 179203 634541
rect 294781 634538 294847 634541
rect 179137 634536 294847 634538
rect 179137 634480 179142 634536
rect 179198 634480 294786 634536
rect 294842 634480 294847 634536
rect 179137 634478 294847 634480
rect 179137 634475 179203 634478
rect 294781 634475 294847 634478
rect 335169 634538 335235 634541
rect 376017 634538 376083 634541
rect 335169 634536 376083 634538
rect 335169 634480 335174 634536
rect 335230 634480 376022 634536
rect 376078 634480 376083 634536
rect 335169 634478 376083 634480
rect 335169 634475 335235 634478
rect 376017 634475 376083 634478
rect 118049 634402 118115 634405
rect 121862 634402 121868 634404
rect 118049 634400 121868 634402
rect 118049 634344 118054 634400
rect 118110 634344 121868 634400
rect 118049 634342 121868 634344
rect 118049 634339 118115 634342
rect 121862 634340 121868 634342
rect 121932 634340 121938 634404
rect 116761 634266 116827 634269
rect 128353 634266 128419 634269
rect 139485 634266 139551 634269
rect 116761 634264 125610 634266
rect 116761 634208 116766 634264
rect 116822 634208 125610 634264
rect 116761 634206 125610 634208
rect 116761 634203 116827 634206
rect 125550 634130 125610 634206
rect 128353 634264 139551 634266
rect 128353 634208 128358 634264
rect 128414 634208 139490 634264
rect 139546 634208 139551 634264
rect 128353 634206 139551 634208
rect 128353 634203 128419 634206
rect 139485 634203 139551 634206
rect 241927 634266 241993 634269
rect 241927 634264 248430 634266
rect 241927 634208 241932 634264
rect 241988 634208 248430 634264
rect 241927 634206 248430 634208
rect 241927 634203 241993 634206
rect 125550 634070 128370 634130
rect 128310 633994 128370 634070
rect 136817 633994 136883 633997
rect 128310 633992 136883 633994
rect 128310 633936 136822 633992
rect 136878 633936 136883 633992
rect 128310 633934 136883 633936
rect 248370 633994 248430 634206
rect 279785 633994 279851 633997
rect 248370 633992 279851 633994
rect 248370 633936 279790 633992
rect 279846 633936 279851 633992
rect 248370 633934 279851 633936
rect 136817 633931 136883 633934
rect 279785 633931 279851 633934
rect 121862 633796 121868 633860
rect 121932 633858 121938 633860
rect 136725 633858 136791 633861
rect 121932 633856 136791 633858
rect 121932 633800 136730 633856
rect 136786 633800 136791 633856
rect 121932 633798 136791 633800
rect 121932 633796 121938 633798
rect 136725 633795 136791 633798
rect 178953 633586 179019 633589
rect 294965 633586 295031 633589
rect 543774 633586 543780 633588
rect 178953 633584 295031 633586
rect 178953 633528 178958 633584
rect 179014 633528 294970 633584
rect 295026 633528 295031 633584
rect 178953 633526 295031 633528
rect 539948 633526 543780 633586
rect 178953 633523 179019 633526
rect 294965 633523 295031 633526
rect 543774 633524 543780 633526
rect 543844 633524 543850 633588
rect 54753 633450 54819 633453
rect 138933 633450 138999 633453
rect 54753 633448 138999 633450
rect 54753 633392 54758 633448
rect 54814 633392 138938 633448
rect 138994 633392 138999 633448
rect 54753 633390 138999 633392
rect 54753 633387 54819 633390
rect 138933 633387 138999 633390
rect 144177 633450 144243 633453
rect 149789 633450 149855 633453
rect 144177 633448 149855 633450
rect 144177 633392 144182 633448
rect 144238 633392 149794 633448
rect 149850 633392 149855 633448
rect 144177 633390 149855 633392
rect 144177 633387 144243 633390
rect 149789 633387 149855 633390
rect 177430 633388 177436 633452
rect 177500 633450 177506 633452
rect 485998 633450 486004 633452
rect 177500 633390 486004 633450
rect 177500 633388 177506 633390
rect 485998 633388 486004 633390
rect 486068 633388 486074 633452
rect 55489 633314 55555 633317
rect 177757 633314 177823 633317
rect 297449 633314 297515 633317
rect 55489 633312 60076 633314
rect 55489 633256 55494 633312
rect 55550 633256 60076 633312
rect 55489 633254 60076 633256
rect 177757 633312 180044 633314
rect 177757 633256 177762 633312
rect 177818 633256 180044 633312
rect 177757 633254 180044 633256
rect 297449 633312 300196 633314
rect 297449 633256 297454 633312
rect 297510 633256 300196 633312
rect 297449 633254 300196 633256
rect 55489 633251 55555 633254
rect 177757 633251 177823 633254
rect 297449 633251 297515 633254
rect 55581 632770 55647 632773
rect 58617 632770 58683 632773
rect 55581 632768 58683 632770
rect 55581 632712 55586 632768
rect 55642 632712 58622 632768
rect 58678 632712 58683 632768
rect 55581 632710 58683 632712
rect 55581 632707 55647 632710
rect 58617 632707 58683 632710
rect -960 632090 480 632180
rect 179086 632164 179092 632228
rect 179156 632226 179162 632228
rect 297633 632226 297699 632229
rect 545062 632226 545068 632228
rect 179156 632166 180044 632226
rect 297633 632224 299674 632226
rect 297633 632168 297638 632224
rect 297694 632168 299674 632224
rect 297633 632166 299674 632168
rect 539948 632166 545068 632226
rect 179156 632164 179162 632166
rect 297633 632163 297699 632166
rect 299614 632158 299674 632166
rect 545062 632164 545068 632166
rect 545132 632164 545138 632228
rect 59494 632098 60076 632158
rect 299614 632098 300196 632158
rect 3417 632090 3483 632093
rect 55581 632092 55647 632093
rect 55581 632090 55628 632092
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect 55536 632088 55628 632090
rect 55536 632032 55586 632088
rect 55536 632030 55628 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 55581 632028 55628 632030
rect 55692 632028 55698 632092
rect 57830 632028 57836 632092
rect 57900 632090 57906 632092
rect 59494 632090 59554 632098
rect 57900 632030 59554 632090
rect 57900 632028 57906 632030
rect 55581 632027 55647 632028
rect 177849 631138 177915 631141
rect 297725 631138 297791 631141
rect 177849 631136 180044 631138
rect 177849 631080 177854 631136
rect 177910 631080 180044 631136
rect 177849 631078 180044 631080
rect 297725 631136 299674 631138
rect 297725 631080 297730 631136
rect 297786 631080 299674 631136
rect 297725 631078 299674 631080
rect 177849 631075 177915 631078
rect 297725 631075 297791 631078
rect 299614 631070 299674 631078
rect 59494 631010 60076 631070
rect 299614 631010 300196 631070
rect 57646 630940 57652 631004
rect 57716 631002 57722 631004
rect 59494 631002 59554 631010
rect 57716 630942 59554 631002
rect 57716 630940 57722 630942
rect 539734 630597 539794 630836
rect 551134 630804 551140 630868
rect 551204 630866 551210 630868
rect 583520 630866 584960 630956
rect 551204 630806 584960 630866
rect 551204 630804 551210 630806
rect 583520 630716 584960 630806
rect 539734 630592 539843 630597
rect 539734 630536 539782 630592
rect 539838 630536 539843 630592
rect 539734 630534 539843 630536
rect 539777 630531 539843 630534
rect 179270 629988 179276 630052
rect 179340 630050 179346 630052
rect 298001 630050 298067 630053
rect 179340 629990 180044 630050
rect 298001 630048 299674 630050
rect 298001 629992 298006 630048
rect 298062 629992 299674 630048
rect 298001 629990 299674 629992
rect 179340 629988 179346 629990
rect 298001 629987 298067 629990
rect 299614 629982 299674 629990
rect 59494 629922 60076 629982
rect 299614 629922 300196 629982
rect 56317 629914 56383 629917
rect 59494 629914 59554 629922
rect 56317 629912 59554 629914
rect 56317 629856 56322 629912
rect 56378 629856 59554 629912
rect 56317 629854 59554 629856
rect 56317 629851 56383 629854
rect 539542 629444 539548 629508
rect 539612 629444 539618 629508
rect 148409 629234 148475 629237
rect 149697 629234 149763 629237
rect 148409 629232 149763 629234
rect 148409 629176 148414 629232
rect 148470 629176 149702 629232
rect 149758 629176 149763 629232
rect 148409 629174 149763 629176
rect 148409 629171 148475 629174
rect 149697 629171 149763 629174
rect 178902 628900 178908 628964
rect 178972 628962 178978 628964
rect 296713 628962 296779 628965
rect 178972 628902 180044 628962
rect 296713 628960 299674 628962
rect 296713 628904 296718 628960
rect 296774 628904 299674 628960
rect 296713 628902 299674 628904
rect 178972 628900 178978 628902
rect 296713 628899 296779 628902
rect 299614 628894 299674 628902
rect 59494 628834 60076 628894
rect 299614 628834 300196 628894
rect 56409 628826 56475 628829
rect 59494 628826 59554 628834
rect 56409 628824 59554 628826
rect 56409 628768 56414 628824
rect 56470 628768 59554 628824
rect 56409 628766 59554 628768
rect 56409 628763 56475 628766
rect 539550 627877 539610 628116
rect 177941 627874 178007 627877
rect 297357 627874 297423 627877
rect 177941 627872 180044 627874
rect 177941 627816 177946 627872
rect 178002 627816 180044 627872
rect 177941 627814 180044 627816
rect 297357 627872 299674 627874
rect 297357 627816 297362 627872
rect 297418 627816 299674 627872
rect 297357 627814 299674 627816
rect 539550 627872 539659 627877
rect 539550 627816 539598 627872
rect 539654 627816 539659 627872
rect 539550 627814 539659 627816
rect 177941 627811 178007 627814
rect 297357 627811 297423 627814
rect 59670 627744 59676 627808
rect 59740 627806 59746 627808
rect 299614 627806 299674 627814
rect 539593 627811 539659 627814
rect 59740 627746 60076 627806
rect 299614 627746 300196 627806
rect 59740 627744 59746 627746
rect 177573 626786 177639 626789
rect 297173 626786 297239 626789
rect 177573 626784 180044 626786
rect 177573 626728 177578 626784
rect 177634 626728 180044 626784
rect 177573 626726 180044 626728
rect 297173 626784 299674 626786
rect 297173 626728 297178 626784
rect 297234 626728 299674 626784
rect 297173 626726 299674 626728
rect 177573 626723 177639 626726
rect 297173 626723 297239 626726
rect 59854 626656 59860 626720
rect 59924 626718 59930 626720
rect 299614 626718 299674 626726
rect 539726 626724 539732 626788
rect 539796 626724 539802 626788
rect 59924 626658 60076 626718
rect 299614 626658 300196 626718
rect 59924 626656 59930 626658
rect 163497 625970 163563 625973
rect 288382 625970 288388 625972
rect 142110 625968 163563 625970
rect 134934 625834 134994 625940
rect 142110 625912 163502 625968
rect 163558 625912 163563 625968
rect 142110 625910 163563 625912
rect 254932 625910 288388 625970
rect 142110 625834 142170 625910
rect 163497 625907 163563 625910
rect 288382 625908 288388 625910
rect 288452 625908 288458 625972
rect 377673 625970 377739 625973
rect 374900 625968 377739 625970
rect 374900 625912 377678 625968
rect 377734 625912 377739 625968
rect 374900 625910 377739 625912
rect 377673 625907 377739 625910
rect 134934 625774 142170 625834
rect 59169 625698 59235 625701
rect 177665 625698 177731 625701
rect 297541 625698 297607 625701
rect 59169 625696 60076 625698
rect 59169 625640 59174 625696
rect 59230 625640 60076 625696
rect 59169 625638 60076 625640
rect 177665 625696 180044 625698
rect 177665 625640 177670 625696
rect 177726 625640 180044 625696
rect 177665 625638 180044 625640
rect 297541 625696 300196 625698
rect 297541 625640 297546 625696
rect 297602 625640 300196 625696
rect 297541 625638 300196 625640
rect 59169 625635 59235 625638
rect 177665 625635 177731 625638
rect 297541 625635 297607 625638
rect 134934 625154 135178 625170
rect 539734 625157 539794 625396
rect 142797 625154 142863 625157
rect 286174 625154 286180 625156
rect 134934 625152 142863 625154
rect 134934 625110 142802 625152
rect 135118 625096 142802 625110
rect 142858 625096 142863 625152
rect 135118 625094 142863 625096
rect 254932 625094 286180 625154
rect 142797 625091 142863 625094
rect 286174 625092 286180 625094
rect 286244 625092 286250 625156
rect 377121 625154 377187 625157
rect 374900 625152 377187 625154
rect 374900 625096 377126 625152
rect 377182 625096 377187 625152
rect 374900 625094 377187 625096
rect 377121 625091 377187 625094
rect 539685 625152 539794 625157
rect 539685 625096 539690 625152
rect 539746 625096 539794 625152
rect 539685 625094 539794 625096
rect 539685 625091 539751 625094
rect 57605 624610 57671 624613
rect 57605 624608 60076 624610
rect 57605 624552 57610 624608
rect 57666 624552 60076 624608
rect 57605 624550 60076 624552
rect 57605 624547 57671 624550
rect 177798 624548 177804 624612
rect 177868 624610 177874 624612
rect 297541 624610 297607 624613
rect 177868 624550 180044 624610
rect 297541 624608 300196 624610
rect 297541 624552 297546 624608
rect 297602 624552 300196 624608
rect 297541 624550 300196 624552
rect 177868 624548 177874 624550
rect 297541 624547 297607 624550
rect 162209 624338 162275 624341
rect 283414 624338 283420 624340
rect 142110 624336 162275 624338
rect 134934 624202 134994 624308
rect 142110 624280 162214 624336
rect 162270 624280 162275 624336
rect 142110 624278 162275 624280
rect 254932 624278 283420 624338
rect 142110 624202 142170 624278
rect 162209 624275 162275 624278
rect 283414 624276 283420 624278
rect 283484 624276 283490 624340
rect 377673 624338 377739 624341
rect 374900 624336 377739 624338
rect 374900 624280 377678 624336
rect 377734 624280 377739 624336
rect 374900 624278 377739 624280
rect 377673 624275 377739 624278
rect 134934 624142 142170 624202
rect 539910 624004 539916 624068
rect 539980 624004 539986 624068
rect 59813 623522 59879 623525
rect 59813 623520 60076 623522
rect 59813 623464 59818 623520
rect 59874 623464 60076 623520
rect 59813 623462 60076 623464
rect 59813 623459 59879 623462
rect 134934 623386 134994 623492
rect 177430 623460 177436 623524
rect 177500 623522 177506 623524
rect 282126 623522 282132 623524
rect 177500 623462 180044 623522
rect 254932 623462 282132 623522
rect 177500 623460 177506 623462
rect 282126 623460 282132 623462
rect 282196 623460 282202 623524
rect 296846 623460 296852 623524
rect 296916 623522 296922 623524
rect 377765 623522 377831 623525
rect 296916 623462 300196 623522
rect 374900 623520 377831 623522
rect 374900 623464 377770 623520
rect 377826 623464 377831 623520
rect 374900 623462 377831 623464
rect 296916 623460 296922 623462
rect 377765 623459 377831 623462
rect 148317 623386 148383 623389
rect 134934 623384 148383 623386
rect 134934 623328 148322 623384
rect 148378 623328 148383 623384
rect 134934 623326 148383 623328
rect 148317 623323 148383 623326
rect 376017 622978 376083 622981
rect 384297 622978 384363 622981
rect 376017 622976 384363 622978
rect 376017 622920 376022 622976
rect 376078 622920 384302 622976
rect 384358 622920 384363 622976
rect 376017 622918 384363 622920
rect 376017 622915 376083 622918
rect 384297 622915 384363 622918
rect 152641 622706 152707 622709
rect 285622 622706 285628 622708
rect 142110 622704 152707 622706
rect 134934 622570 134994 622676
rect 142110 622648 152646 622704
rect 152702 622648 152707 622704
rect 142110 622646 152707 622648
rect 254932 622646 285628 622706
rect 142110 622570 142170 622646
rect 152641 622643 152707 622646
rect 285622 622644 285628 622646
rect 285692 622644 285698 622708
rect 377213 622706 377279 622709
rect 374900 622704 377279 622706
rect 374900 622648 377218 622704
rect 377274 622648 377279 622704
rect 374900 622646 377279 622648
rect 377213 622643 377279 622646
rect 134934 622510 142170 622570
rect 539918 622437 539978 622676
rect 59077 622434 59143 622437
rect 59077 622432 60076 622434
rect 59077 622376 59082 622432
rect 59138 622376 60076 622432
rect 59077 622374 60076 622376
rect 59077 622371 59143 622374
rect 177798 622372 177804 622436
rect 177868 622434 177874 622436
rect 297909 622434 297975 622437
rect 177868 622374 180044 622434
rect 297909 622432 300196 622434
rect 297909 622376 297914 622432
rect 297970 622376 300196 622432
rect 297909 622374 300196 622376
rect 539918 622432 540027 622437
rect 539918 622376 539966 622432
rect 540022 622376 540027 622432
rect 539918 622374 540027 622376
rect 177868 622372 177874 622374
rect 297909 622371 297975 622374
rect 539961 622371 540027 622374
rect 174537 621890 174603 621893
rect 288566 621890 288572 621892
rect 142110 621888 174603 621890
rect 134934 621754 134994 621860
rect 142110 621832 174542 621888
rect 174598 621832 174603 621888
rect 142110 621830 174603 621832
rect 254932 621830 288572 621890
rect 142110 621754 142170 621830
rect 174537 621827 174603 621830
rect 288566 621828 288572 621830
rect 288636 621828 288642 621892
rect 377029 621890 377095 621893
rect 374900 621888 377095 621890
rect 374900 621832 377034 621888
rect 377090 621832 377095 621888
rect 374900 621830 377095 621832
rect 377029 621827 377095 621830
rect 134934 621694 142170 621754
rect 296478 621692 296484 621756
rect 296548 621692 296554 621756
rect 296486 621618 296546 621692
rect 296486 621558 296730 621618
rect 57789 621346 57855 621349
rect 57789 621344 60076 621346
rect 57789 621288 57794 621344
rect 57850 621288 60076 621344
rect 57789 621286 60076 621288
rect 57789 621283 57855 621286
rect 177246 621284 177252 621348
rect 177316 621346 177322 621348
rect 296670 621346 296730 621558
rect 177316 621286 180044 621346
rect 296670 621286 300196 621346
rect 177316 621284 177322 621286
rect 146937 621210 147003 621213
rect 134934 621208 147003 621210
rect 134934 621152 146942 621208
rect 146998 621152 147003 621208
rect 134934 621150 147003 621152
rect 134934 621044 134994 621150
rect 146937 621147 147003 621150
rect 539918 621077 539978 621316
rect 285806 621074 285812 621076
rect 254932 621014 285812 621074
rect 285806 621012 285812 621014
rect 285876 621012 285882 621076
rect 377029 621074 377095 621077
rect 374900 621072 377095 621074
rect 374900 621016 377034 621072
rect 377090 621016 377095 621072
rect 374900 621014 377095 621016
rect 377029 621011 377095 621014
rect 539869 621072 539978 621077
rect 539869 621016 539874 621072
rect 539930 621016 539978 621072
rect 539869 621014 539978 621016
rect 539869 621011 539935 621014
rect 58433 620258 58499 620261
rect 58433 620256 60076 620258
rect 58433 620200 58438 620256
rect 58494 620200 60076 620256
rect 58433 620198 60076 620200
rect 58433 620195 58499 620198
rect 134934 619714 134994 620228
rect 163998 620196 164004 620260
rect 164068 620258 164074 620260
rect 297449 620258 297515 620261
rect 164068 620198 180044 620258
rect 297449 620256 300196 620258
rect 164068 620196 164074 620198
rect 254902 620122 254962 620228
rect 297449 620200 297454 620256
rect 297510 620200 300196 620256
rect 297449 620198 300196 620200
rect 297449 620195 297515 620198
rect 298134 620122 298140 620124
rect 254902 620062 298140 620122
rect 298134 620060 298140 620062
rect 298204 620060 298210 620124
rect 137277 619714 137343 619717
rect 134934 619712 137343 619714
rect 134934 619656 137282 619712
rect 137338 619656 137343 619712
rect 134934 619654 137343 619656
rect 374870 619714 374930 620228
rect 541198 619986 541204 619988
rect 539948 619926 541204 619986
rect 541198 619924 541204 619926
rect 541268 619924 541274 619988
rect 378041 619714 378107 619717
rect 374870 619712 378107 619714
rect 374870 619656 378046 619712
rect 378102 619656 378107 619712
rect 374870 619654 378107 619656
rect 137277 619651 137343 619654
rect 378041 619651 378107 619654
rect 164877 619442 164943 619445
rect 291142 619442 291148 619444
rect 142110 619440 164943 619442
rect 134934 619306 134994 619412
rect 142110 619384 164882 619440
rect 164938 619384 164943 619440
rect 142110 619382 164943 619384
rect 254932 619382 291148 619442
rect 142110 619306 142170 619382
rect 164877 619379 164943 619382
rect 291142 619380 291148 619382
rect 291212 619380 291218 619444
rect 375373 619442 375439 619445
rect 374900 619440 375439 619442
rect 374900 619384 375378 619440
rect 375434 619384 375439 619440
rect 374900 619382 375439 619384
rect 375373 619379 375439 619382
rect -960 619170 480 619260
rect 134934 619246 142170 619306
rect 29126 619170 29132 619172
rect -960 619110 29132 619170
rect -960 619020 480 619110
rect 29126 619108 29132 619110
rect 29196 619108 29202 619172
rect 58985 619170 59051 619173
rect 58985 619168 60076 619170
rect 58985 619112 58990 619168
rect 59046 619112 60076 619168
rect 58985 619110 60076 619112
rect 58985 619107 59051 619110
rect 177614 619108 177620 619172
rect 177684 619170 177690 619172
rect 297633 619170 297699 619173
rect 177684 619110 180044 619170
rect 297633 619168 300196 619170
rect 297633 619112 297638 619168
rect 297694 619112 300196 619168
rect 297633 619110 300196 619112
rect 177684 619108 177690 619110
rect 297633 619107 297699 619110
rect 169017 618626 169083 618629
rect 291326 618626 291332 618628
rect 142110 618624 169083 618626
rect 134934 618490 134994 618596
rect 142110 618568 169022 618624
rect 169078 618568 169083 618624
rect 142110 618566 169083 618568
rect 254932 618566 291332 618626
rect 142110 618490 142170 618566
rect 169017 618563 169083 618566
rect 291326 618564 291332 618566
rect 291396 618564 291402 618628
rect 375649 618626 375715 618629
rect 543958 618626 543964 618628
rect 374900 618624 375715 618626
rect 374900 618568 375654 618624
rect 375710 618568 375715 618624
rect 374900 618566 375715 618568
rect 539948 618566 543964 618626
rect 375649 618563 375715 618566
rect 543958 618564 543964 618566
rect 544028 618564 544034 618628
rect 134934 618430 142170 618490
rect 49601 618082 49667 618085
rect 49601 618080 60076 618082
rect 49601 618024 49606 618080
rect 49662 618024 60076 618080
rect 49601 618022 60076 618024
rect 49601 618019 49667 618022
rect 177430 618020 177436 618084
rect 177500 618082 177506 618084
rect 297357 618082 297423 618085
rect 177500 618022 180044 618082
rect 297357 618080 300196 618082
rect 297357 618024 297362 618080
rect 297418 618024 300196 618080
rect 297357 618022 300196 618024
rect 177500 618020 177506 618022
rect 297357 618019 297423 618022
rect 173249 617810 173315 617813
rect 293861 617810 293927 617813
rect 378317 617810 378383 617813
rect 142110 617808 173315 617810
rect 134934 617674 134994 617780
rect 142110 617752 173254 617808
rect 173310 617752 173315 617808
rect 142110 617750 173315 617752
rect 254932 617808 293927 617810
rect 254932 617752 293866 617808
rect 293922 617752 293927 617808
rect 254932 617750 293927 617752
rect 374900 617808 378383 617810
rect 374900 617752 378322 617808
rect 378378 617752 378383 617808
rect 374900 617750 378383 617752
rect 142110 617674 142170 617750
rect 173249 617747 173315 617750
rect 293861 617747 293927 617750
rect 378317 617747 378383 617750
rect 134934 617614 142170 617674
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 545246 617266 545252 617268
rect 539948 617206 545252 617266
rect 545246 617204 545252 617206
rect 545316 617204 545322 617268
rect 134934 617070 142170 617130
rect 57881 616994 57947 616997
rect 57881 616992 60076 616994
rect 57881 616936 57886 616992
rect 57942 616936 60076 616992
rect 134934 616964 134994 617070
rect 142110 616994 142170 617070
rect 273846 617068 273852 617132
rect 273916 617130 273922 617132
rect 273916 617070 296730 617130
rect 273916 617068 273922 617070
rect 166349 616994 166415 616997
rect 142110 616992 166415 616994
rect 57881 616934 60076 616936
rect 142110 616936 166354 616992
rect 166410 616936 166415 616992
rect 142110 616934 166415 616936
rect 57881 616931 57947 616934
rect 166349 616931 166415 616934
rect 177614 616932 177620 616996
rect 177684 616994 177690 616996
rect 292798 616994 292804 616996
rect 177684 616934 180044 616994
rect 254932 616934 292804 616994
rect 177684 616932 177690 616934
rect 292798 616932 292804 616934
rect 292868 616932 292874 616996
rect 296670 616994 296730 617070
rect 296670 616934 300196 616994
rect 374502 616725 374562 616964
rect 374502 616720 374611 616725
rect 374502 616664 374550 616720
rect 374606 616664 374611 616720
rect 374502 616662 374611 616664
rect 374545 616659 374611 616662
rect 167637 616178 167703 616181
rect 292614 616178 292620 616180
rect 142110 616176 167703 616178
rect 134934 616042 134994 616148
rect 142110 616120 167642 616176
rect 167698 616120 167703 616176
rect 142110 616118 167703 616120
rect 254932 616118 292620 616178
rect 142110 616042 142170 616118
rect 167637 616115 167703 616118
rect 292614 616116 292620 616118
rect 292684 616116 292690 616180
rect 378041 616178 378107 616181
rect 374900 616176 378107 616178
rect 374900 616120 378046 616176
rect 378102 616120 378107 616176
rect 374900 616118 378107 616120
rect 378041 616115 378107 616118
rect 134934 615982 142170 616042
rect 57513 615906 57579 615909
rect 57513 615904 60076 615906
rect 57513 615848 57518 615904
rect 57574 615848 60076 615904
rect 57513 615846 60076 615848
rect 57513 615843 57579 615846
rect 177062 615844 177068 615908
rect 177132 615906 177138 615908
rect 281441 615906 281507 615909
rect 543365 615906 543431 615909
rect 177132 615846 180044 615906
rect 281441 615904 300196 615906
rect 281441 615848 281446 615904
rect 281502 615848 300196 615904
rect 281441 615846 300196 615848
rect 539948 615904 543431 615906
rect 539948 615848 543370 615904
rect 543426 615848 543431 615904
rect 539948 615846 543431 615848
rect 177132 615844 177138 615846
rect 281441 615843 281507 615846
rect 543365 615843 543431 615846
rect 134934 615438 142170 615498
rect 134934 615332 134994 615438
rect 142110 615362 142170 615438
rect 173934 615362 173940 615364
rect 142110 615302 173940 615362
rect 173934 615300 173940 615302
rect 174004 615300 174010 615364
rect 294454 615362 294460 615364
rect 254932 615302 294460 615362
rect 294454 615300 294460 615302
rect 294524 615300 294530 615364
rect 374686 614821 374746 615332
rect 58893 614818 58959 614821
rect 58893 614816 60076 614818
rect 58893 614760 58898 614816
rect 58954 614760 60076 614816
rect 58893 614758 60076 614760
rect 58893 614755 58959 614758
rect 166758 614756 166764 614820
rect 166828 614818 166834 614820
rect 298001 614818 298067 614821
rect 166828 614758 180044 614818
rect 298001 614816 300196 614818
rect 298001 614760 298006 614816
rect 298062 614760 300196 614816
rect 298001 614758 300196 614760
rect 374686 614816 374795 614821
rect 374686 614760 374734 614816
rect 374790 614760 374795 614816
rect 374686 614758 374795 614760
rect 166828 614756 166834 614758
rect 298001 614755 298067 614758
rect 374729 614755 374795 614758
rect 134934 614622 142170 614682
rect 134934 614516 134994 614622
rect 142110 614546 142170 614622
rect 171777 614546 171843 614549
rect 294822 614546 294828 614548
rect 142110 614544 171843 614546
rect 142110 614488 171782 614544
rect 171838 614488 171843 614544
rect 142110 614486 171843 614488
rect 254932 614486 294828 614546
rect 171777 614483 171843 614486
rect 294822 614484 294828 614486
rect 294892 614484 294898 614548
rect 375925 614546 375991 614549
rect 542997 614546 543063 614549
rect 374900 614544 375991 614546
rect 374900 614488 375930 614544
rect 375986 614488 375991 614544
rect 374900 614486 375991 614488
rect 539948 614544 543063 614546
rect 539948 614488 543002 614544
rect 543058 614488 543063 614544
rect 539948 614486 543063 614488
rect 375925 614483 375991 614486
rect 542997 614483 543063 614486
rect 298502 613866 298508 613868
rect 296670 613806 298508 613866
rect 57697 613730 57763 613733
rect 57697 613728 60076 613730
rect 57697 613672 57702 613728
rect 57758 613672 60076 613728
rect 57697 613670 60076 613672
rect 57697 613667 57763 613670
rect 134934 613594 134994 613700
rect 177982 613668 177988 613732
rect 178052 613730 178058 613732
rect 296670 613730 296730 613806
rect 298502 613804 298508 613806
rect 298572 613804 298578 613868
rect 378685 613730 378751 613733
rect 178052 613670 180044 613730
rect 254932 613670 296730 613730
rect 298326 613670 300196 613730
rect 374900 613728 378751 613730
rect 374900 613672 378690 613728
rect 378746 613672 378751 613728
rect 374900 613670 378751 613672
rect 178052 613668 178058 613670
rect 178166 613594 178172 613596
rect 134934 613534 178172 613594
rect 178166 613532 178172 613534
rect 178236 613532 178242 613596
rect 271086 613532 271092 613596
rect 271156 613594 271162 613596
rect 298326 613594 298386 613670
rect 378685 613667 378751 613670
rect 487153 613730 487219 613733
rect 487153 613728 490084 613730
rect 487153 613672 487158 613728
rect 487214 613672 490084 613728
rect 487153 613670 490084 613672
rect 487153 613667 487219 613670
rect 271156 613534 298386 613594
rect 271156 613532 271162 613534
rect 543181 613186 543247 613189
rect 539948 613184 543247 613186
rect 539948 613128 543186 613184
rect 543242 613128 543247 613184
rect 539948 613126 543247 613128
rect 543181 613123 543247 613126
rect 134934 612990 142170 613050
rect 134934 612884 134994 612990
rect 142110 612914 142170 612990
rect 166257 612914 166323 612917
rect 293166 612914 293172 612916
rect 142110 612912 166323 612914
rect 142110 612856 166262 612912
rect 166318 612856 166323 612912
rect 142110 612854 166323 612856
rect 254932 612854 293172 612914
rect 166257 612851 166323 612854
rect 293166 612852 293172 612854
rect 293236 612852 293242 612916
rect 378409 612914 378475 612917
rect 374900 612912 378475 612914
rect 374900 612856 378414 612912
rect 378470 612856 378475 612912
rect 374900 612854 378475 612856
rect 378409 612851 378475 612854
rect 177297 612778 177363 612781
rect 177798 612778 177804 612780
rect 177297 612776 177804 612778
rect 177297 612720 177302 612776
rect 177358 612720 177804 612776
rect 177297 612718 177804 612720
rect 177297 612715 177363 612718
rect 177798 612716 177804 612718
rect 177868 612716 177874 612780
rect 292798 612716 292804 612780
rect 292868 612778 292874 612780
rect 293769 612778 293835 612781
rect 292868 612776 293835 612778
rect 292868 612720 293774 612776
rect 293830 612720 293835 612776
rect 292868 612718 293835 612720
rect 292868 612716 292874 612718
rect 293769 612715 293835 612718
rect 539501 612778 539567 612781
rect 542813 612778 542879 612781
rect 539501 612776 542879 612778
rect 539501 612720 539506 612776
rect 539562 612720 542818 612776
rect 542874 612720 542879 612776
rect 539501 612718 542879 612720
rect 539501 612715 539567 612718
rect 542813 612715 542879 612718
rect 57329 612642 57395 612645
rect 57329 612640 60076 612642
rect 57329 612584 57334 612640
rect 57390 612584 60076 612640
rect 57329 612582 60076 612584
rect 57329 612579 57395 612582
rect 177798 612580 177804 612644
rect 177868 612642 177874 612644
rect 298001 612642 298067 612645
rect 177868 612582 180044 612642
rect 298001 612640 300196 612642
rect 298001 612584 298006 612640
rect 298062 612584 300196 612640
rect 298001 612582 300196 612584
rect 177868 612580 177874 612582
rect 298001 612579 298067 612582
rect 134934 612174 142170 612234
rect 134934 612068 134994 612174
rect 142110 612098 142170 612174
rect 175774 612098 175780 612100
rect 142110 612038 175780 612098
rect 175774 612036 175780 612038
rect 175844 612036 175850 612100
rect 295558 612098 295564 612100
rect 254932 612038 295564 612098
rect 295558 612036 295564 612038
rect 295628 612036 295634 612100
rect 377121 612098 377187 612101
rect 374900 612096 377187 612098
rect 374900 612040 377126 612096
rect 377182 612040 377187 612096
rect 374900 612038 377187 612040
rect 377121 612035 377187 612038
rect 543089 611826 543155 611829
rect 539948 611824 543155 611826
rect 539948 611768 543094 611824
rect 543150 611768 543155 611824
rect 539948 611766 543155 611768
rect 543089 611763 543155 611766
rect 177614 611628 177620 611692
rect 177684 611690 177690 611692
rect 177941 611690 178007 611693
rect 177684 611688 178007 611690
rect 177684 611632 177946 611688
rect 178002 611632 178007 611688
rect 177684 611630 178007 611632
rect 177684 611628 177690 611630
rect 177941 611627 178007 611630
rect 59721 611554 59787 611557
rect 59721 611552 60076 611554
rect 59721 611496 59726 611552
rect 59782 611496 60076 611552
rect 59721 611494 60076 611496
rect 59721 611491 59787 611494
rect 177246 611492 177252 611556
rect 177316 611554 177322 611556
rect 177316 611494 180044 611554
rect 177316 611492 177322 611494
rect 286358 611492 286364 611556
rect 286428 611554 286434 611556
rect 286428 611494 300196 611554
rect 286428 611492 286434 611494
rect 177430 611356 177436 611420
rect 177500 611418 177506 611420
rect 177665 611418 177731 611421
rect 177500 611416 177731 611418
rect 177500 611360 177670 611416
rect 177726 611360 177731 611416
rect 177500 611358 177731 611360
rect 177500 611356 177506 611358
rect 177665 611355 177731 611358
rect 384297 611418 384363 611421
rect 391197 611418 391263 611421
rect 384297 611416 391263 611418
rect 384297 611360 384302 611416
rect 384358 611360 391202 611416
rect 391258 611360 391263 611416
rect 384297 611358 391263 611360
rect 384297 611355 384363 611358
rect 391197 611355 391263 611358
rect 170254 611282 170260 611284
rect 134934 611146 134994 611252
rect 142110 611222 170260 611282
rect 142110 611146 142170 611222
rect 170254 611220 170260 611222
rect 170324 611220 170330 611284
rect 295374 611282 295380 611284
rect 254932 611222 295380 611282
rect 295374 611220 295380 611222
rect 295444 611220 295450 611284
rect 376937 611282 377003 611285
rect 374900 611280 377003 611282
rect 374900 611224 376942 611280
rect 376998 611224 377003 611280
rect 374900 611222 377003 611224
rect 376937 611219 377003 611222
rect 134934 611086 142170 611146
rect 177062 610676 177068 610740
rect 177132 610738 177138 610740
rect 177205 610738 177271 610741
rect 177132 610736 177271 610738
rect 177132 610680 177210 610736
rect 177266 610680 177271 610736
rect 177132 610678 177271 610680
rect 177132 610676 177138 610678
rect 177205 610675 177271 610678
rect 539409 610738 539475 610741
rect 542905 610738 542971 610741
rect 539409 610736 542971 610738
rect 539409 610680 539414 610736
rect 539470 610680 542910 610736
rect 542966 610680 542971 610736
rect 539409 610678 542971 610680
rect 539409 610675 539475 610678
rect 542905 610675 542971 610678
rect 134934 610542 142170 610602
rect 58801 610466 58867 610469
rect 58801 610464 60076 610466
rect 58801 610408 58806 610464
rect 58862 610408 60076 610464
rect 134934 610436 134994 610542
rect 142110 610466 142170 610542
rect 174629 610466 174695 610469
rect 142110 610464 174695 610466
rect 58801 610406 60076 610408
rect 142110 610408 174634 610464
rect 174690 610408 174695 610464
rect 142110 610406 174695 610408
rect 58801 610403 58867 610406
rect 174629 610403 174695 610406
rect 177614 610404 177620 610468
rect 177684 610466 177690 610468
rect 298001 610466 298067 610469
rect 375465 610466 375531 610469
rect 543222 610466 543228 610468
rect 177684 610406 180044 610466
rect 298001 610464 300196 610466
rect 177684 610404 177690 610406
rect 254902 610330 254962 610436
rect 298001 610408 298006 610464
rect 298062 610408 300196 610464
rect 298001 610406 300196 610408
rect 374900 610464 375531 610466
rect 374900 610408 375470 610464
rect 375526 610408 375531 610464
rect 374900 610406 375531 610408
rect 539948 610406 543228 610466
rect 298001 610403 298067 610406
rect 375465 610403 375531 610406
rect 543222 610404 543228 610406
rect 543292 610404 543298 610468
rect 298318 610330 298324 610332
rect 254902 610270 298324 610330
rect 298318 610268 298324 610270
rect 298388 610268 298394 610332
rect 177849 609786 177915 609789
rect 177982 609786 177988 609788
rect 134934 609726 142170 609786
rect 134934 609620 134994 609726
rect 142110 609650 142170 609726
rect 177849 609784 177988 609786
rect 177849 609728 177854 609784
rect 177910 609728 177988 609784
rect 177849 609726 177988 609728
rect 177849 609723 177915 609726
rect 177982 609724 177988 609726
rect 178052 609724 178058 609788
rect 174813 609650 174879 609653
rect 299606 609650 299612 609652
rect 142110 609648 174879 609650
rect 142110 609592 174818 609648
rect 174874 609592 174879 609648
rect 142110 609590 174879 609592
rect 254932 609590 299612 609650
rect 174813 609587 174879 609590
rect 299606 609588 299612 609590
rect 299676 609588 299682 609652
rect 375557 609650 375623 609653
rect 374900 609648 375623 609650
rect 374900 609592 375562 609648
rect 375618 609592 375623 609648
rect 374900 609590 375623 609592
rect 375557 609587 375623 609590
rect 56133 609378 56199 609381
rect 56133 609376 60076 609378
rect 56133 609320 56138 609376
rect 56194 609320 60076 609376
rect 56133 609318 60076 609320
rect 56133 609315 56199 609318
rect 177798 609316 177804 609380
rect 177868 609378 177874 609380
rect 177868 609318 180044 609378
rect 177868 609316 177874 609318
rect 296846 609316 296852 609380
rect 296916 609378 296922 609380
rect 296916 609318 300196 609378
rect 296916 609316 296922 609318
rect 542854 609106 542860 609108
rect 539948 609046 542860 609106
rect 542854 609044 542860 609046
rect 542924 609044 542930 609108
rect 134934 608910 142170 608970
rect 134934 608804 134994 608910
rect 142110 608834 142170 608910
rect 169293 608834 169359 608837
rect 299238 608834 299244 608836
rect 142110 608832 169359 608834
rect 142110 608776 169298 608832
rect 169354 608776 169359 608832
rect 142110 608774 169359 608776
rect 254932 608774 299244 608834
rect 169293 608771 169359 608774
rect 299238 608772 299244 608774
rect 299308 608772 299314 608836
rect 375414 608834 375420 608836
rect 374900 608774 375420 608834
rect 375414 608772 375420 608774
rect 375484 608772 375490 608836
rect 298134 608500 298140 608564
rect 298204 608562 298210 608564
rect 299289 608562 299355 608565
rect 298204 608560 299355 608562
rect 298204 608504 299294 608560
rect 299350 608504 299355 608560
rect 298204 608502 299355 608504
rect 298204 608500 298210 608502
rect 299289 608499 299355 608502
rect 58709 608290 58775 608293
rect 58709 608288 60076 608290
rect 58709 608232 58714 608288
rect 58770 608232 60076 608288
rect 58709 608230 60076 608232
rect 58709 608227 58775 608230
rect 165470 608228 165476 608292
rect 165540 608290 165546 608292
rect 297817 608290 297883 608293
rect 165540 608230 180044 608290
rect 297817 608288 300196 608290
rect 297817 608232 297822 608288
rect 297878 608232 300196 608288
rect 297817 608230 300196 608232
rect 165540 608228 165546 608230
rect 297817 608227 297883 608230
rect 134934 608094 142170 608154
rect 134934 607988 134994 608094
rect 142110 608018 142170 608094
rect 178677 608018 178743 608021
rect 298686 608018 298692 608020
rect 142110 608016 178743 608018
rect 142110 607960 178682 608016
rect 178738 607960 178743 608016
rect 142110 607958 178743 607960
rect 254932 607958 298692 608018
rect 178677 607955 178743 607958
rect 298686 607956 298692 607958
rect 298756 607956 298762 608020
rect 376753 608018 376819 608021
rect 374900 608016 376819 608018
rect 374900 607960 376758 608016
rect 376814 607960 376819 608016
rect 374900 607958 376819 607960
rect 376753 607955 376819 607958
rect 539358 607684 539364 607748
rect 539428 607684 539434 607748
rect 57237 607202 57303 607205
rect 173157 607202 173223 607205
rect 57237 607200 60076 607202
rect 57237 607144 57242 607200
rect 57298 607144 60076 607200
rect 142110 607200 173223 607202
rect 57237 607142 60076 607144
rect 57237 607139 57303 607142
rect 134934 607066 134994 607172
rect 142110 607144 173162 607200
rect 173218 607144 173223 607200
rect 142110 607142 173223 607144
rect 142110 607066 142170 607142
rect 173157 607139 173223 607142
rect 176878 607140 176884 607204
rect 176948 607202 176954 607204
rect 294638 607202 294644 607204
rect 176948 607142 180044 607202
rect 254932 607142 294644 607202
rect 176948 607140 176954 607142
rect 294638 607140 294644 607142
rect 294708 607140 294714 607204
rect 376845 607202 376911 607205
rect 296670 607142 300196 607202
rect 374900 607200 376911 607202
rect 374900 607144 376850 607200
rect 376906 607144 376911 607200
rect 374900 607142 376911 607144
rect 134934 607006 142170 607066
rect 177246 607004 177252 607068
rect 177316 607066 177322 607068
rect 177389 607066 177455 607069
rect 177316 607064 177455 607066
rect 177316 607008 177394 607064
rect 177450 607008 177455 607064
rect 177316 607006 177455 607008
rect 177316 607004 177322 607006
rect 177389 607003 177455 607006
rect 177573 607066 177639 607069
rect 177982 607066 177988 607068
rect 177573 607064 177988 607066
rect 177573 607008 177578 607064
rect 177634 607008 177988 607064
rect 177573 607006 177988 607008
rect 177573 607003 177639 607006
rect 177982 607004 177988 607006
rect 178052 607004 178058 607068
rect 271270 607004 271276 607068
rect 271340 607066 271346 607068
rect 296670 607066 296730 607142
rect 376845 607139 376911 607142
rect 271340 607006 296730 607066
rect 271340 607004 271346 607006
rect 134934 606462 142170 606522
rect 134934 606356 134994 606462
rect 142110 606386 142170 606462
rect 171869 606386 171935 606389
rect 272006 606386 272012 606388
rect 142110 606384 171935 606386
rect 142110 606328 171874 606384
rect 171930 606328 171935 606384
rect 142110 606326 171935 606328
rect 254932 606326 272012 606386
rect 171869 606323 171935 606326
rect 272006 606324 272012 606326
rect 272076 606324 272082 606388
rect 378041 606386 378107 606389
rect 542670 606386 542676 606388
rect 374900 606384 378107 606386
rect 374900 606328 378046 606384
rect 378102 606328 378107 606384
rect 374900 606326 378107 606328
rect 539948 606326 542676 606386
rect 378041 606323 378107 606326
rect 542670 606324 542676 606326
rect 542740 606324 542746 606388
rect -960 606114 480 606204
rect 11646 606114 11652 606116
rect -960 606054 11652 606114
rect -960 605964 480 606054
rect 11646 606052 11652 606054
rect 11716 606052 11722 606116
rect 59813 606114 59879 606117
rect 297725 606114 297791 606117
rect 59813 606112 60076 606114
rect 59813 606056 59818 606112
rect 59874 606056 60076 606112
rect 59813 606054 60076 606056
rect 177622 606054 180044 606114
rect 297725 606112 300196 606114
rect 297725 606056 297730 606112
rect 297786 606056 300196 606112
rect 297725 606054 300196 606056
rect 59813 606051 59879 606054
rect 177430 605780 177436 605844
rect 177500 605842 177506 605844
rect 177622 605842 177682 606054
rect 297725 606051 297791 606054
rect 177500 605782 177682 605842
rect 177500 605780 177506 605782
rect 170489 605570 170555 605573
rect 299054 605570 299060 605572
rect 142110 605568 170555 605570
rect 134934 605434 134994 605540
rect 142110 605512 170494 605568
rect 170550 605512 170555 605568
rect 142110 605510 170555 605512
rect 254932 605510 299060 605570
rect 142110 605434 142170 605510
rect 170489 605507 170555 605510
rect 299054 605508 299060 605510
rect 299124 605508 299130 605572
rect 377949 605570 378015 605573
rect 374900 605568 378015 605570
rect 374900 605512 377954 605568
rect 378010 605512 378015 605568
rect 374900 605510 378015 605512
rect 377949 605507 378015 605510
rect 134934 605374 142170 605434
rect 136909 605162 136975 605165
rect 179321 605162 179387 605165
rect 136909 605160 179387 605162
rect 136909 605104 136914 605160
rect 136970 605104 179326 605160
rect 179382 605104 179387 605160
rect 136909 605102 179387 605104
rect 136909 605099 136975 605102
rect 179321 605099 179387 605102
rect 57053 605026 57119 605029
rect 57053 605024 60076 605026
rect 57053 604968 57058 605024
rect 57114 604968 60076 605024
rect 57053 604966 60076 604968
rect 57053 604963 57119 604966
rect 177062 604964 177068 605028
rect 177132 605026 177138 605028
rect 177132 604966 180044 605026
rect 177132 604964 177138 604966
rect 296662 604964 296668 605028
rect 296732 605026 296738 605028
rect 296732 604966 300196 605026
rect 296732 604964 296738 604966
rect 175958 604754 175964 604756
rect 134934 604618 134994 604724
rect 142110 604694 175964 604754
rect 142110 604618 142170 604694
rect 175958 604692 175964 604694
rect 176028 604692 176034 604756
rect 269798 604754 269804 604756
rect 254932 604694 269804 604754
rect 269798 604692 269804 604694
rect 269868 604692 269874 604756
rect 378041 604754 378107 604757
rect 374900 604752 378107 604754
rect 374900 604696 378046 604752
rect 378102 604696 378107 604752
rect 374900 604694 378107 604696
rect 378041 604691 378107 604694
rect 134934 604558 142170 604618
rect 134793 604482 134859 604485
rect 136909 604482 136975 604485
rect 134793 604480 136975 604482
rect 134793 604424 134798 604480
rect 134854 604424 136914 604480
rect 136970 604424 136975 604480
rect 134793 604422 136975 604424
rect 134793 604419 134859 604422
rect 136909 604419 136975 604422
rect 177614 604420 177620 604484
rect 177684 604482 177690 604484
rect 177757 604482 177823 604485
rect 177684 604480 177823 604482
rect 177684 604424 177762 604480
rect 177818 604424 177823 604480
rect 177684 604422 177823 604424
rect 177684 604420 177690 604422
rect 177757 604419 177823 604422
rect 298502 604420 298508 604484
rect 298572 604482 298578 604484
rect 299381 604482 299447 604485
rect 298572 604480 299447 604482
rect 298572 604424 299386 604480
rect 299442 604424 299447 604480
rect 298572 604422 299447 604424
rect 298572 604420 298578 604422
rect 299381 604419 299447 604422
rect 539317 604482 539383 604485
rect 539550 604482 539610 604996
rect 539317 604480 539610 604482
rect 539317 604424 539322 604480
rect 539378 604424 539610 604480
rect 539317 604422 539610 604424
rect 539317 604419 539383 604422
rect 583520 604060 584960 604300
rect 57421 603938 57487 603941
rect 167729 603938 167795 603941
rect 57421 603936 60076 603938
rect 57421 603880 57426 603936
rect 57482 603880 60076 603936
rect 142110 603936 167795 603938
rect 57421 603878 60076 603880
rect 57421 603875 57487 603878
rect 134934 603802 134994 603908
rect 142110 603880 167734 603936
rect 167790 603880 167795 603936
rect 142110 603878 167795 603880
rect 142110 603802 142170 603878
rect 167729 603875 167795 603878
rect 173750 603876 173756 603940
rect 173820 603938 173826 603940
rect 262806 603938 262812 603940
rect 173820 603878 180044 603938
rect 254932 603878 262812 603938
rect 173820 603876 173826 603878
rect 262806 603876 262812 603878
rect 262876 603876 262882 603940
rect 280654 603876 280660 603940
rect 280724 603938 280730 603940
rect 378041 603938 378107 603941
rect 280724 603878 300196 603938
rect 374900 603936 378107 603938
rect 374900 603880 378046 603936
rect 378102 603880 378107 603936
rect 374900 603878 378107 603880
rect 280724 603876 280730 603878
rect 378041 603875 378107 603878
rect 134934 603742 142170 603802
rect 540094 603666 540100 603668
rect 539948 603606 540100 603666
rect 540094 603604 540100 603606
rect 540164 603604 540170 603668
rect 146293 603258 146359 603261
rect 148409 603258 148475 603261
rect 134934 603198 142170 603258
rect 134934 603092 134994 603198
rect 142110 603122 142170 603198
rect 146293 603256 148475 603258
rect 146293 603200 146298 603256
rect 146354 603200 148414 603256
rect 148470 603200 148475 603256
rect 146293 603198 148475 603200
rect 146293 603195 146359 603198
rect 148409 603195 148475 603198
rect 169201 603122 169267 603125
rect 265934 603122 265940 603124
rect 142110 603120 169267 603122
rect 142110 603064 169206 603120
rect 169262 603064 169267 603120
rect 142110 603062 169267 603064
rect 254932 603062 265940 603122
rect 169201 603059 169267 603062
rect 265934 603060 265940 603062
rect 266004 603060 266010 603124
rect 378041 603122 378107 603125
rect 374900 603120 378107 603122
rect 374900 603064 378046 603120
rect 378102 603064 378107 603120
rect 374900 603062 378107 603064
rect 378041 603059 378107 603062
rect 138841 602986 138907 602989
rect 176561 602986 176627 602989
rect 138841 602984 176627 602986
rect 138841 602928 138846 602984
rect 138902 602928 176566 602984
rect 176622 602928 176627 602984
rect 138841 602926 176627 602928
rect 138841 602923 138907 602926
rect 176561 602923 176627 602926
rect 57145 602850 57211 602853
rect 57145 602848 60076 602850
rect 57145 602792 57150 602848
rect 57206 602792 60076 602848
rect 57145 602790 60076 602792
rect 57145 602787 57211 602790
rect 177614 602788 177620 602852
rect 177684 602850 177690 602852
rect 177684 602790 180044 602850
rect 177684 602788 177690 602790
rect 255814 602788 255820 602852
rect 255884 602850 255890 602852
rect 255884 602790 300196 602850
rect 255884 602788 255890 602790
rect 176193 602306 176259 602309
rect 280838 602306 280844 602308
rect 142110 602304 176259 602306
rect 134934 602170 134994 602276
rect 142110 602248 176198 602304
rect 176254 602248 176259 602304
rect 142110 602246 176259 602248
rect 254932 602246 280844 602306
rect 142110 602170 142170 602246
rect 176193 602243 176259 602246
rect 280838 602244 280844 602246
rect 280908 602244 280914 602308
rect 377622 602306 377628 602308
rect 374900 602246 377628 602306
rect 377622 602244 377628 602246
rect 377692 602244 377698 602308
rect 134934 602110 142170 602170
rect 176561 601898 176627 601901
rect 176561 601896 178050 601898
rect 176561 601840 176566 601896
rect 176622 601840 178050 601896
rect 176561 601838 178050 601840
rect 176561 601835 176627 601838
rect 54661 601762 54727 601765
rect 177573 601762 177639 601765
rect 177798 601762 177804 601764
rect 54661 601760 60076 601762
rect 54661 601704 54666 601760
rect 54722 601704 60076 601760
rect 54661 601702 60076 601704
rect 177573 601760 177804 601762
rect 177573 601704 177578 601760
rect 177634 601704 177804 601760
rect 177573 601702 177804 601704
rect 54661 601699 54727 601702
rect 177573 601699 177639 601702
rect 177798 601700 177804 601702
rect 177868 601700 177874 601764
rect 177990 601762 178050 601838
rect 538254 601836 538260 601900
rect 538324 601898 538330 601900
rect 539409 601898 539475 601901
rect 538324 601896 539475 601898
rect 538324 601840 539414 601896
rect 539470 601840 539475 601896
rect 538324 601838 539475 601840
rect 538324 601836 538330 601838
rect 539409 601835 539475 601838
rect 295057 601762 295123 601765
rect 177990 601702 180044 601762
rect 295057 601760 300196 601762
rect 295057 601704 295062 601760
rect 295118 601704 300196 601760
rect 295057 601702 300196 601704
rect 295057 601699 295123 601702
rect 538438 601700 538444 601764
rect 538508 601762 538514 601764
rect 539501 601762 539567 601765
rect 538508 601760 539567 601762
rect 538508 601704 539506 601760
rect 539562 601704 539567 601760
rect 538508 601702 539567 601704
rect 538508 601700 538514 601702
rect 539501 601699 539567 601702
rect 140037 601626 140103 601629
rect 178033 601626 178099 601629
rect 140037 601624 178099 601626
rect 140037 601568 140042 601624
rect 140098 601568 178038 601624
rect 178094 601568 178099 601624
rect 140037 601566 178099 601568
rect 140037 601563 140103 601566
rect 178033 601563 178099 601566
rect 164969 601490 165035 601493
rect 266854 601490 266860 601492
rect 142110 601488 165035 601490
rect 134934 601354 134994 601460
rect 142110 601432 164974 601488
rect 165030 601432 165035 601488
rect 142110 601430 165035 601432
rect 254932 601430 266860 601490
rect 142110 601354 142170 601430
rect 164969 601427 165035 601430
rect 266854 601428 266860 601430
rect 266924 601428 266930 601492
rect 376753 601490 376819 601493
rect 374900 601488 376819 601490
rect 374900 601432 376758 601488
rect 376814 601432 376819 601488
rect 374900 601430 376819 601432
rect 376753 601427 376819 601430
rect 134934 601294 142170 601354
rect 543089 601084 543155 601085
rect 543038 601082 543044 601084
rect 542998 601022 543044 601082
rect 543108 601080 543155 601084
rect 543150 601024 543155 601080
rect 543038 601020 543044 601022
rect 543108 601020 543155 601024
rect 543089 601019 543155 601020
rect 54845 600674 54911 600677
rect 171961 600674 172027 600677
rect 54845 600672 60076 600674
rect 54845 600616 54850 600672
rect 54906 600616 60076 600672
rect 142110 600672 172027 600674
rect 54845 600614 60076 600616
rect 54845 600611 54911 600614
rect 134934 600538 134994 600644
rect 142110 600616 171966 600672
rect 172022 600616 172027 600672
rect 142110 600614 172027 600616
rect 142110 600538 142170 600614
rect 171961 600611 172027 600614
rect 178033 600674 178099 600677
rect 179045 600674 179111 600677
rect 277894 600674 277900 600676
rect 178033 600672 180044 600674
rect 178033 600616 178038 600672
rect 178094 600616 179050 600672
rect 179106 600616 180044 600672
rect 178033 600614 180044 600616
rect 254932 600614 277900 600674
rect 178033 600611 178099 600614
rect 179045 600611 179111 600614
rect 277894 600612 277900 600614
rect 277964 600612 277970 600676
rect 291929 600674 291995 600677
rect 375465 600674 375531 600677
rect 291929 600672 300196 600674
rect 291929 600616 291934 600672
rect 291990 600616 300196 600672
rect 291929 600614 300196 600616
rect 374900 600672 375531 600674
rect 374900 600616 375470 600672
rect 375526 600616 375531 600672
rect 374900 600614 375531 600616
rect 291929 600611 291995 600614
rect 375465 600611 375531 600614
rect 134934 600478 142170 600538
rect 537334 600476 537340 600540
rect 537404 600538 537410 600540
rect 542670 600538 542676 600540
rect 537404 600478 542676 600538
rect 537404 600476 537410 600478
rect 542670 600476 542676 600478
rect 542740 600476 542746 600540
rect 138933 600266 138999 600269
rect 484025 600266 484091 600269
rect 497365 600266 497431 600269
rect 138933 600264 171150 600266
rect 138933 600208 138938 600264
rect 138994 600208 171150 600264
rect 138933 600206 171150 600208
rect 138933 600203 138999 600206
rect 170581 599858 170647 599861
rect 142110 599856 170647 599858
rect 134934 599722 134994 599828
rect 142110 599800 170586 599856
rect 170642 599800 170647 599856
rect 142110 599798 170647 599800
rect 142110 599722 142170 599798
rect 170581 599795 170647 599798
rect 134934 599662 142170 599722
rect 54753 599586 54819 599589
rect 171090 599586 171150 600206
rect 484025 600264 497431 600266
rect 484025 600208 484030 600264
rect 484086 600208 497370 600264
rect 497426 600208 497431 600264
rect 484025 600206 497431 600208
rect 484025 600203 484091 600206
rect 497365 600203 497431 600206
rect 536005 600266 536071 600269
rect 536005 600264 538874 600266
rect 536005 600208 536010 600264
rect 536066 600208 538874 600264
rect 536005 600206 538874 600208
rect 536005 600203 536071 600206
rect 488441 600130 488507 600133
rect 507853 600130 507919 600133
rect 488441 600128 507919 600130
rect 488441 600072 488446 600128
rect 488502 600072 507858 600128
rect 507914 600072 507919 600128
rect 488441 600070 507919 600072
rect 488441 600067 488507 600070
rect 507853 600067 507919 600070
rect 534574 600068 534580 600132
rect 534644 600130 534650 600132
rect 538581 600130 538647 600133
rect 534644 600128 538647 600130
rect 534644 600072 538586 600128
rect 538642 600072 538647 600128
rect 534644 600070 538647 600072
rect 538814 600130 538874 600206
rect 542670 600204 542676 600268
rect 542740 600266 542746 600268
rect 543181 600266 543247 600269
rect 543917 600266 543983 600269
rect 542740 600264 543247 600266
rect 542740 600208 543186 600264
rect 543242 600208 543247 600264
rect 542740 600206 543247 600208
rect 542740 600204 542746 600206
rect 543181 600203 543247 600206
rect 543414 600264 543983 600266
rect 543414 600208 543922 600264
rect 543978 600208 543983 600264
rect 543414 600206 543983 600208
rect 543414 600130 543474 600206
rect 543917 600203 543983 600206
rect 538814 600070 543474 600130
rect 534644 600068 534650 600070
rect 538581 600067 538647 600070
rect 484117 599994 484183 599997
rect 504081 599994 504147 599997
rect 484117 599992 504147 599994
rect 484117 599936 484122 599992
rect 484178 599936 504086 599992
rect 504142 599936 504147 599992
rect 484117 599934 504147 599936
rect 484117 599931 484183 599934
rect 504081 599931 504147 599934
rect 526294 599932 526300 599996
rect 526364 599994 526370 599996
rect 540094 599994 540100 599996
rect 526364 599934 540100 599994
rect 526364 599932 526370 599934
rect 540094 599932 540100 599934
rect 540164 599932 540170 599996
rect 256734 599858 256740 599860
rect 254932 599798 256740 599858
rect 256734 599796 256740 599798
rect 256804 599796 256810 599860
rect 378593 599858 378659 599861
rect 374900 599856 378659 599858
rect 374900 599800 378598 599856
rect 378654 599800 378659 599856
rect 374900 599798 378659 599800
rect 378593 599795 378659 599798
rect 486969 599858 487035 599861
rect 508037 599858 508103 599861
rect 486969 599856 508103 599858
rect 486969 599800 486974 599856
rect 487030 599800 508042 599856
rect 508098 599800 508103 599856
rect 486969 599798 508103 599800
rect 486969 599795 487035 599798
rect 508037 599795 508103 599798
rect 531957 599858 532023 599861
rect 545205 599858 545271 599861
rect 531957 599856 545271 599858
rect 531957 599800 531962 599856
rect 532018 599800 545210 599856
rect 545266 599800 545271 599856
rect 531957 599798 545271 599800
rect 531957 599795 532023 599798
rect 545205 599795 545271 599798
rect 478505 599722 478571 599725
rect 499573 599722 499639 599725
rect 478505 599720 499639 599722
rect 478505 599664 478510 599720
rect 478566 599664 499578 599720
rect 499634 599664 499639 599720
rect 478505 599662 499639 599664
rect 478505 599659 478571 599662
rect 499573 599659 499639 599662
rect 522246 599660 522252 599724
rect 522316 599722 522322 599724
rect 543958 599722 543964 599724
rect 522316 599662 543964 599722
rect 522316 599660 522322 599662
rect 543958 599660 543964 599662
rect 544028 599660 544034 599724
rect 178953 599586 179019 599589
rect 294965 599586 295031 599589
rect 391197 599586 391263 599589
rect 403617 599586 403683 599589
rect 54753 599584 60076 599586
rect 54753 599528 54758 599584
rect 54814 599528 60076 599584
rect 54753 599526 60076 599528
rect 171090 599584 180044 599586
rect 171090 599528 178958 599584
rect 179014 599528 180044 599584
rect 171090 599526 180044 599528
rect 294965 599584 300196 599586
rect 294965 599528 294970 599584
rect 295026 599528 300196 599584
rect 294965 599526 300196 599528
rect 391197 599584 403683 599586
rect 391197 599528 391202 599584
rect 391258 599528 403622 599584
rect 403678 599528 403683 599584
rect 391197 599526 403683 599528
rect 54753 599523 54819 599526
rect 178953 599523 179019 599526
rect 294965 599523 295031 599526
rect 391197 599523 391263 599526
rect 403617 599523 403683 599526
rect 462313 599586 462379 599589
rect 495709 599586 495775 599589
rect 462313 599584 495775 599586
rect 462313 599528 462318 599584
rect 462374 599528 495714 599584
rect 495770 599528 495775 599584
rect 462313 599526 495775 599528
rect 462313 599523 462379 599526
rect 495709 599523 495775 599526
rect 522430 599524 522436 599588
rect 522500 599586 522506 599588
rect 545062 599586 545068 599588
rect 522500 599526 545068 599586
rect 522500 599524 522506 599526
rect 545062 599524 545068 599526
rect 545132 599524 545138 599588
rect 537518 599388 537524 599452
rect 537588 599450 537594 599452
rect 545246 599450 545252 599452
rect 537588 599390 545252 599450
rect 537588 599388 537594 599390
rect 545246 599388 545252 599390
rect 545316 599388 545322 599452
rect 374637 599178 374703 599181
rect 134934 599118 142170 599178
rect 134934 599012 134994 599118
rect 142110 599042 142170 599118
rect 374637 599176 374746 599178
rect 374637 599120 374642 599176
rect 374698 599120 374746 599176
rect 374637 599115 374746 599120
rect 533286 599116 533292 599180
rect 533356 599178 533362 599180
rect 535729 599178 535795 599181
rect 533356 599176 535795 599178
rect 533356 599120 535734 599176
rect 535790 599120 535795 599176
rect 533356 599118 535795 599120
rect 533356 599116 533362 599118
rect 535729 599115 535795 599118
rect 175917 599042 175983 599045
rect 295742 599042 295748 599044
rect 142110 599040 175983 599042
rect 142110 598984 175922 599040
rect 175978 598984 175983 599040
rect 142110 598982 175983 598984
rect 254932 598982 295748 599042
rect 175917 598979 175983 598982
rect 295742 598980 295748 598982
rect 295812 598980 295818 599044
rect 374686 599012 374746 599115
rect 511901 599042 511967 599045
rect 536833 599042 536899 599045
rect 511901 599040 536899 599042
rect 511901 598984 511906 599040
rect 511962 598984 536838 599040
rect 536894 598984 536899 599040
rect 511901 598982 536899 598984
rect 511901 598979 511967 598982
rect 536833 598979 536899 598982
rect 56225 598498 56291 598501
rect 179137 598498 179203 598501
rect 294781 598498 294847 598501
rect 56225 598496 60076 598498
rect 56225 598440 56230 598496
rect 56286 598440 60076 598496
rect 56225 598438 60076 598440
rect 161430 598496 180044 598498
rect 161430 598440 179142 598496
rect 179198 598440 180044 598496
rect 161430 598438 180044 598440
rect 294781 598496 300196 598498
rect 294781 598440 294786 598496
rect 294842 598440 300196 598496
rect 294781 598438 300196 598440
rect 56225 598435 56291 598438
rect 137461 598362 137527 598365
rect 161430 598362 161490 598438
rect 179137 598435 179203 598438
rect 294781 598435 294847 598438
rect 137461 598360 161490 598362
rect 137461 598304 137466 598360
rect 137522 598304 161490 598360
rect 137461 598302 161490 598304
rect 523677 598362 523743 598365
rect 532141 598362 532207 598365
rect 523677 598360 532207 598362
rect 523677 598304 523682 598360
rect 523738 598304 532146 598360
rect 532202 598304 532207 598360
rect 523677 598302 532207 598304
rect 137461 598299 137527 598302
rect 523677 598299 523743 598302
rect 532141 598299 532207 598302
rect 536046 598300 536052 598364
rect 536116 598362 536122 598364
rect 542353 598362 542419 598365
rect 536116 598360 542419 598362
rect 536116 598304 542358 598360
rect 542414 598304 542419 598360
rect 536116 598302 542419 598304
rect 536116 598300 536122 598302
rect 542353 598299 542419 598302
rect 275134 598226 275140 598228
rect 134934 597682 134994 598196
rect 254932 598166 275140 598226
rect 275134 598164 275140 598166
rect 275204 598164 275210 598228
rect 376845 598226 376911 598229
rect 374900 598224 376911 598226
rect 374900 598168 376850 598224
rect 376906 598168 376911 598224
rect 374900 598166 376911 598168
rect 376845 598163 376911 598166
rect 490414 598164 490420 598228
rect 490484 598226 490490 598228
rect 492121 598226 492187 598229
rect 490484 598224 492187 598226
rect 490484 598168 492126 598224
rect 492182 598168 492187 598224
rect 490484 598166 492187 598168
rect 490484 598164 490490 598166
rect 492121 598163 492187 598166
rect 492990 598164 492996 598228
rect 493060 598226 493066 598228
rect 493501 598226 493567 598229
rect 493060 598224 493567 598226
rect 493060 598168 493506 598224
rect 493562 598168 493567 598224
rect 493060 598166 493567 598168
rect 493060 598164 493066 598166
rect 493501 598163 493567 598166
rect 494094 598164 494100 598228
rect 494164 598226 494170 598228
rect 494881 598226 494947 598229
rect 494164 598224 494947 598226
rect 494164 598168 494886 598224
rect 494942 598168 494947 598224
rect 494164 598166 494947 598168
rect 494164 598164 494170 598166
rect 494881 598163 494947 598166
rect 496854 598164 496860 598228
rect 496924 598226 496930 598228
rect 497641 598226 497707 598229
rect 496924 598224 497707 598226
rect 496924 598168 497646 598224
rect 497702 598168 497707 598224
rect 496924 598166 497707 598168
rect 496924 598164 496930 598166
rect 497641 598163 497707 598166
rect 530526 598164 530532 598228
rect 530596 598226 530602 598228
rect 542445 598226 542511 598229
rect 530596 598224 542511 598226
rect 530596 598168 542450 598224
rect 542506 598168 542511 598224
rect 530596 598166 542511 598168
rect 530596 598164 530602 598166
rect 542445 598163 542511 598166
rect 529197 598090 529263 598093
rect 537661 598090 537727 598093
rect 529197 598088 537727 598090
rect 529197 598032 529202 598088
rect 529258 598032 537666 598088
rect 537722 598032 537727 598088
rect 529197 598030 537727 598032
rect 529197 598027 529263 598030
rect 537661 598027 537727 598030
rect 137645 597682 137711 597685
rect 134934 597680 137711 597682
rect 134934 597624 137650 597680
rect 137706 597624 137711 597680
rect 134934 597622 137711 597624
rect 137645 597619 137711 597622
rect 294822 597484 294828 597548
rect 294892 597546 294898 597548
rect 295057 597546 295123 597549
rect 294892 597544 295123 597546
rect 294892 597488 295062 597544
rect 295118 597488 295123 597544
rect 294892 597486 295123 597488
rect 294892 597484 294898 597486
rect 295057 597483 295123 597486
rect 48037 597410 48103 597413
rect 167913 597410 167979 597413
rect 48037 597408 60076 597410
rect 48037 597352 48042 597408
rect 48098 597352 60076 597408
rect 142110 597408 167979 597410
rect 48037 597350 60076 597352
rect 48037 597347 48103 597350
rect 134934 597274 134994 597380
rect 142110 597352 167918 597408
rect 167974 597352 167979 597408
rect 142110 597350 167979 597352
rect 142110 597274 142170 597350
rect 167913 597347 167979 597350
rect 170673 597410 170739 597413
rect 179229 597410 179295 597413
rect 294689 597410 294755 597413
rect 375557 597410 375623 597413
rect 170673 597408 180044 597410
rect 170673 597352 170678 597408
rect 170734 597352 179234 597408
rect 179290 597352 180044 597408
rect 294689 597408 300196 597410
rect 170673 597350 180044 597352
rect 170673 597347 170739 597350
rect 179229 597347 179295 597350
rect 134934 597214 142170 597274
rect 254902 597274 254962 597380
rect 294689 597352 294694 597408
rect 294750 597352 300196 597408
rect 294689 597350 300196 597352
rect 374900 597408 375623 597410
rect 374900 597352 375562 597408
rect 375618 597352 375623 597408
rect 374900 597350 375623 597352
rect 294689 597347 294755 597350
rect 375557 597347 375623 597350
rect 295006 597274 295012 597276
rect 254902 597214 295012 597274
rect 295006 597212 295012 597214
rect 295076 597212 295082 597276
rect 501454 596804 501460 596868
rect 501524 596866 501530 596868
rect 542537 596866 542603 596869
rect 501524 596864 542603 596866
rect 501524 596808 542542 596864
rect 542598 596808 542603 596864
rect 501524 596806 542603 596808
rect 501524 596804 501530 596806
rect 542537 596803 542603 596806
rect 166441 596594 166507 596597
rect 256918 596594 256924 596596
rect 142110 596592 166507 596594
rect 134934 596458 134994 596564
rect 142110 596536 166446 596592
rect 166502 596536 166507 596592
rect 142110 596534 166507 596536
rect 254932 596534 256924 596594
rect 142110 596458 142170 596534
rect 166441 596531 166507 596534
rect 256918 596532 256924 596534
rect 256988 596532 256994 596596
rect 375833 596594 375899 596597
rect 374900 596592 375899 596594
rect 374900 596536 375838 596592
rect 375894 596536 375899 596592
rect 374900 596534 375899 596536
rect 375833 596531 375899 596534
rect 134934 596398 142170 596458
rect 54937 596322 55003 596325
rect 179321 596322 179387 596325
rect 294873 596322 294939 596325
rect 54937 596320 60076 596322
rect 54937 596264 54942 596320
rect 54998 596264 60076 596320
rect 54937 596262 60076 596264
rect 179321 596320 180044 596322
rect 179321 596264 179326 596320
rect 179382 596264 180044 596320
rect 179321 596262 180044 596264
rect 294873 596320 300196 596322
rect 294873 596264 294878 596320
rect 294934 596264 300196 596320
rect 294873 596262 300196 596264
rect 54937 596259 55003 596262
rect 179321 596259 179387 596262
rect 294873 596259 294939 596262
rect 134934 595854 142170 595914
rect 134934 595748 134994 595854
rect 142110 595778 142170 595854
rect 167821 595778 167887 595781
rect 257102 595778 257108 595780
rect 142110 595776 167887 595778
rect 142110 595720 167826 595776
rect 167882 595720 167887 595776
rect 142110 595718 167887 595720
rect 254932 595718 257108 595778
rect 167821 595715 167887 595718
rect 257102 595716 257108 595718
rect 257172 595716 257178 595780
rect 378501 595778 378567 595781
rect 374900 595776 378567 595778
rect 374900 595720 378506 595776
rect 378562 595720 378567 595776
rect 374900 595718 378567 595720
rect 378501 595715 378567 595718
rect 508446 595444 508452 595508
rect 508516 595506 508522 595508
rect 542854 595506 542860 595508
rect 508516 595446 542860 595506
rect 508516 595444 508522 595446
rect 542854 595444 542860 595446
rect 542924 595444 542930 595508
rect 56961 595234 57027 595237
rect 172329 595234 172395 595237
rect 298001 595234 298067 595237
rect 56961 595232 60076 595234
rect 56961 595176 56966 595232
rect 57022 595176 60076 595232
rect 56961 595174 60076 595176
rect 171090 595232 180044 595234
rect 171090 595176 172334 595232
rect 172390 595176 180044 595232
rect 171090 595174 180044 595176
rect 298001 595232 300196 595234
rect 298001 595176 298006 595232
rect 298062 595176 300196 595232
rect 298001 595174 300196 595176
rect 56961 595171 57027 595174
rect 134934 595038 142170 595098
rect 134934 594932 134994 595038
rect 142110 594962 142170 595038
rect 170397 594962 170463 594965
rect 142110 594960 170463 594962
rect 142110 594904 170402 594960
rect 170458 594904 170463 594960
rect 142110 594902 170463 594904
rect 170397 594899 170463 594902
rect 160829 594826 160895 594829
rect 171090 594826 171150 595174
rect 172329 595171 172395 595174
rect 298001 595171 298067 595174
rect 268142 594962 268148 594964
rect 254932 594902 268148 594962
rect 268142 594900 268148 594902
rect 268212 594900 268218 594964
rect 378041 594962 378107 594965
rect 374900 594960 378107 594962
rect 374900 594904 378046 594960
rect 378102 594904 378107 594960
rect 374900 594902 378107 594904
rect 378041 594899 378107 594902
rect 160829 594824 171150 594826
rect 160829 594768 160834 594824
rect 160890 594768 171150 594824
rect 160829 594766 171150 594768
rect 160829 594763 160895 594766
rect 256734 594764 256740 594828
rect 256804 594826 256810 594828
rect 257981 594826 258047 594829
rect 256804 594824 258047 594826
rect 256804 594768 257986 594824
rect 258042 594768 258047 594824
rect 256804 594766 258047 594768
rect 256804 594764 256810 594766
rect 257981 594763 258047 594766
rect 542997 594826 543063 594829
rect 543590 594826 543596 594828
rect 542997 594824 543596 594826
rect 542997 594768 543002 594824
rect 543058 594768 543596 594824
rect 542997 594766 543596 594768
rect 542997 594763 543063 594766
rect 543590 594764 543596 594766
rect 543660 594764 543666 594828
rect 50705 594146 50771 594149
rect 269614 594146 269620 594148
rect 50705 594144 60076 594146
rect 50705 594088 50710 594144
rect 50766 594088 60076 594144
rect 50705 594086 60076 594088
rect 50705 594083 50771 594086
rect 134934 594010 134994 594116
rect 175230 594086 180044 594146
rect 254932 594086 269620 594146
rect 175089 594010 175155 594013
rect 134934 594008 175155 594010
rect 134934 593952 175094 594008
rect 175150 593952 175155 594008
rect 134934 593950 175155 593952
rect 175089 593947 175155 593950
rect 160737 593466 160803 593469
rect 174353 593466 174419 593469
rect 175230 593466 175290 594086
rect 269614 594084 269620 594086
rect 269684 594084 269690 594148
rect 285213 594146 285279 594149
rect 375741 594146 375807 594149
rect 285213 594144 300196 594146
rect 285213 594088 285218 594144
rect 285274 594088 300196 594144
rect 285213 594086 300196 594088
rect 374900 594144 375807 594146
rect 374900 594088 375746 594144
rect 375802 594088 375807 594144
rect 374900 594086 375807 594088
rect 285213 594083 285279 594086
rect 375741 594083 375807 594086
rect 506974 593948 506980 594012
rect 507044 594010 507050 594012
rect 543222 594010 543228 594012
rect 507044 593950 543228 594010
rect 507044 593948 507050 593950
rect 543222 593948 543228 593950
rect 543292 593948 543298 594012
rect 543365 593468 543431 593469
rect 543365 593466 543412 593468
rect 160737 593464 175290 593466
rect 160737 593408 160742 593464
rect 160798 593408 174358 593464
rect 174414 593408 175290 593464
rect 160737 593406 175290 593408
rect 543320 593464 543412 593466
rect 543320 593408 543370 593464
rect 543320 593406 543412 593408
rect 160737 593403 160803 593406
rect 174353 593403 174419 593406
rect 543365 593404 543412 593406
rect 543476 593404 543482 593468
rect 543365 593403 543431 593404
rect 170949 593330 171015 593333
rect 296294 593330 296300 593332
rect 142110 593328 171015 593330
rect 134934 593194 134994 593300
rect 142110 593272 170954 593328
rect 171010 593272 171015 593328
rect 142110 593270 171015 593272
rect 254932 593270 296300 593330
rect 142110 593194 142170 593270
rect 170949 593267 171015 593270
rect 296294 593268 296300 593270
rect 296364 593268 296370 593332
rect 377949 593330 378015 593333
rect 374900 593328 378015 593330
rect 374900 593272 377954 593328
rect 378010 593272 378015 593328
rect 374900 593270 378015 593272
rect 377949 593267 378015 593270
rect -960 592908 480 593148
rect 134934 593134 142170 593194
rect 50521 593058 50587 593061
rect 169753 593058 169819 593061
rect 171041 593058 171107 593061
rect 285121 593058 285187 593061
rect 50521 593056 60076 593058
rect 50521 593000 50526 593056
rect 50582 593000 60076 593056
rect 50521 592998 60076 593000
rect 169753 593056 180044 593058
rect 169753 593000 169758 593056
rect 169814 593000 171046 593056
rect 171102 593000 180044 593056
rect 169753 592998 180044 593000
rect 285121 593056 300196 593058
rect 285121 593000 285126 593056
rect 285182 593000 300196 593056
rect 285121 592998 300196 593000
rect 50521 592995 50587 592998
rect 169753 592995 169819 592998
rect 171041 592995 171107 592998
rect 285121 592995 285187 592998
rect 134934 592590 142170 592650
rect 134934 592484 134994 592590
rect 142110 592514 142170 592590
rect 518014 592588 518020 592652
rect 518084 592650 518090 592652
rect 543038 592650 543044 592652
rect 518084 592590 543044 592650
rect 518084 592588 518090 592590
rect 543038 592588 543044 592590
rect 543108 592588 543114 592652
rect 179229 592514 179295 592517
rect 294822 592514 294828 592516
rect 142110 592512 179295 592514
rect 142110 592456 179234 592512
rect 179290 592456 179295 592512
rect 142110 592454 179295 592456
rect 254932 592454 294828 592514
rect 179229 592451 179295 592454
rect 294822 592452 294828 592454
rect 294892 592452 294898 592516
rect 378041 592514 378107 592517
rect 374900 592512 378107 592514
rect 374900 592456 378046 592512
rect 378102 592456 378107 592512
rect 374900 592454 378107 592456
rect 378041 592451 378107 592454
rect 160921 592106 160987 592109
rect 169753 592106 169819 592109
rect 160921 592104 169819 592106
rect 160921 592048 160926 592104
rect 160982 592048 169758 592104
rect 169814 592048 169819 592104
rect 160921 592046 169819 592048
rect 160921 592043 160987 592046
rect 169753 592043 169819 592046
rect 294454 592044 294460 592108
rect 294524 592106 294530 592108
rect 295241 592106 295307 592109
rect 294524 592104 295307 592106
rect 294524 592048 295246 592104
rect 295302 592048 295307 592104
rect 294524 592046 295307 592048
rect 294524 592044 294530 592046
rect 295241 592043 295307 592046
rect 54845 591970 54911 591973
rect 173801 591970 173867 591973
rect 285397 591970 285463 591973
rect 54845 591968 60076 591970
rect 54845 591912 54850 591968
rect 54906 591912 60076 591968
rect 54845 591910 60076 591912
rect 173801 591968 180044 591970
rect 173801 591912 173806 591968
rect 173862 591912 180044 591968
rect 173801 591910 180044 591912
rect 285397 591968 300196 591970
rect 285397 591912 285402 591968
rect 285458 591912 300196 591968
rect 285397 591910 300196 591912
rect 54845 591907 54911 591910
rect 173801 591907 173867 591910
rect 285397 591907 285463 591910
rect 134934 591774 142170 591834
rect 134934 591668 134994 591774
rect 142110 591698 142170 591774
rect 172053 591698 172119 591701
rect 298870 591698 298876 591700
rect 142110 591696 172119 591698
rect 142110 591640 172058 591696
rect 172114 591640 172119 591696
rect 142110 591638 172119 591640
rect 254932 591638 298876 591698
rect 172053 591635 172119 591638
rect 298870 591636 298876 591638
rect 298940 591636 298946 591700
rect 383837 591698 383903 591701
rect 374900 591696 383903 591698
rect 374900 591640 383842 591696
rect 383898 591640 383903 591696
rect 374900 591638 383903 591640
rect 383837 591635 383903 591638
rect 298318 591364 298324 591428
rect 298388 591426 298394 591428
rect 299197 591426 299263 591429
rect 298388 591424 299263 591426
rect 298388 591368 299202 591424
rect 299258 591368 299263 591424
rect 298388 591366 299263 591368
rect 298388 591364 298394 591366
rect 299197 591363 299263 591366
rect 163773 591018 163839 591021
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 134934 590958 142170 591018
rect 56961 590882 57027 590885
rect 56961 590880 60076 590882
rect 56961 590824 56966 590880
rect 57022 590824 60076 590880
rect 134934 590852 134994 590958
rect 142110 590882 142170 590958
rect 163773 591016 176578 591018
rect 163773 590960 163778 591016
rect 163834 590960 176578 591016
rect 163773 590958 176578 590960
rect 163773 590955 163839 590958
rect 174905 590882 174971 590885
rect 142110 590880 174971 590882
rect 56961 590822 60076 590824
rect 142110 590824 174910 590880
rect 174966 590824 174971 590880
rect 142110 590822 174971 590824
rect 176518 590882 176578 590958
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 178585 590882 178651 590885
rect 265750 590882 265756 590884
rect 176518 590880 180044 590882
rect 176518 590824 178590 590880
rect 178646 590824 180044 590880
rect 176518 590822 180044 590824
rect 254932 590822 265756 590882
rect 56961 590819 57027 590822
rect 174905 590819 174971 590822
rect 178585 590819 178651 590822
rect 265750 590820 265756 590822
rect 265820 590820 265826 590884
rect 298001 590882 298067 590885
rect 378041 590882 378107 590885
rect 298001 590880 300196 590882
rect 298001 590824 298006 590880
rect 298062 590824 300196 590880
rect 298001 590822 300196 590824
rect 374900 590880 378107 590882
rect 374900 590824 378046 590880
rect 378102 590824 378107 590880
rect 583520 590868 584960 590958
rect 374900 590822 378107 590824
rect 298001 590819 298067 590822
rect 378041 590819 378107 590822
rect 161105 590746 161171 590749
rect 173801 590746 173867 590749
rect 161105 590744 173867 590746
rect 161105 590688 161110 590744
rect 161166 590688 173806 590744
rect 173862 590688 173867 590744
rect 161105 590686 173867 590688
rect 161105 590683 161171 590686
rect 173801 590683 173867 590686
rect 141417 590610 141483 590613
rect 144177 590610 144243 590613
rect 141417 590608 144243 590610
rect 141417 590552 141422 590608
rect 141478 590552 144182 590608
rect 144238 590552 144243 590608
rect 141417 590550 144243 590552
rect 141417 590547 141483 590550
rect 144177 590547 144243 590550
rect 295558 590548 295564 590612
rect 295628 590610 295634 590612
rect 296621 590610 296687 590613
rect 295628 590608 296687 590610
rect 295628 590552 296626 590608
rect 296682 590552 296687 590608
rect 295628 590550 296687 590552
rect 295628 590548 295634 590550
rect 296621 590547 296687 590550
rect 134934 590142 142170 590202
rect 134934 590036 134994 590142
rect 142110 590066 142170 590142
rect 173433 590066 173499 590069
rect 296110 590066 296116 590068
rect 142110 590064 173499 590066
rect 142110 590008 173438 590064
rect 173494 590008 173499 590064
rect 142110 590006 173499 590008
rect 254932 590006 296116 590066
rect 173433 590003 173499 590006
rect 296110 590004 296116 590006
rect 296180 590004 296186 590068
rect 378041 590066 378107 590069
rect 374900 590064 378107 590066
rect 374900 590008 378046 590064
rect 378102 590008 378107 590064
rect 374900 590006 378107 590008
rect 378041 590003 378107 590006
rect 56961 589794 57027 589797
rect 176561 589794 176627 589797
rect 285489 589794 285555 589797
rect 56961 589792 60076 589794
rect 56961 589736 56966 589792
rect 57022 589736 60076 589792
rect 56961 589734 60076 589736
rect 176561 589792 180044 589794
rect 176561 589736 176566 589792
rect 176622 589736 180044 589792
rect 176561 589734 180044 589736
rect 285489 589792 300196 589794
rect 285489 589736 285494 589792
rect 285550 589736 300196 589792
rect 285489 589734 300196 589736
rect 56961 589731 57027 589734
rect 176561 589731 176627 589734
rect 285489 589731 285555 589734
rect 163865 589386 163931 589389
rect 176561 589386 176627 589389
rect 163865 589384 176627 589386
rect 163865 589328 163870 589384
rect 163926 589328 176566 589384
rect 176622 589328 176627 589384
rect 163865 589326 176627 589328
rect 163865 589323 163931 589326
rect 176561 589323 176627 589326
rect 170857 589250 170923 589253
rect 268326 589250 268332 589252
rect 142110 589248 170923 589250
rect 134934 589114 134994 589220
rect 142110 589192 170862 589248
rect 170918 589192 170923 589248
rect 142110 589190 170923 589192
rect 254932 589190 268332 589250
rect 142110 589114 142170 589190
rect 170857 589187 170923 589190
rect 268326 589188 268332 589190
rect 268396 589188 268402 589252
rect 378041 589250 378107 589253
rect 374900 589248 378107 589250
rect 374900 589192 378046 589248
rect 378102 589192 378107 589248
rect 374900 589190 378107 589192
rect 378041 589187 378107 589190
rect 134934 589054 142170 589114
rect 54937 588706 55003 588709
rect 179321 588706 179387 588709
rect 287973 588706 288039 588709
rect 54937 588704 60076 588706
rect 54937 588648 54942 588704
rect 54998 588648 60076 588704
rect 54937 588646 60076 588648
rect 176886 588704 180044 588706
rect 176886 588648 179326 588704
rect 179382 588648 180044 588704
rect 176886 588646 180044 588648
rect 287973 588704 300196 588706
rect 287973 588648 287978 588704
rect 288034 588648 300196 588704
rect 287973 588646 300196 588648
rect 54937 588643 55003 588646
rect 134934 588510 142170 588570
rect 134934 588404 134994 588510
rect 142110 588434 142170 588510
rect 173341 588434 173407 588437
rect 142110 588432 173407 588434
rect 142110 588376 173346 588432
rect 173402 588376 173407 588432
rect 142110 588374 173407 588376
rect 173341 588371 173407 588374
rect 163957 588298 164023 588301
rect 176886 588298 176946 588646
rect 179321 588643 179387 588646
rect 287973 588643 288039 588646
rect 277158 588434 277164 588436
rect 254932 588374 277164 588434
rect 277158 588372 277164 588374
rect 277228 588372 277234 588436
rect 377029 588434 377095 588437
rect 374900 588432 377095 588434
rect 374900 588376 377034 588432
rect 377090 588376 377095 588432
rect 374900 588374 377095 588376
rect 377029 588371 377095 588374
rect 163957 588296 176946 588298
rect 163957 588240 163962 588296
rect 164018 588240 176946 588296
rect 163957 588238 176946 588240
rect 163957 588235 164023 588238
rect 53189 587618 53255 587621
rect 173801 587618 173867 587621
rect 284886 587618 284892 587620
rect 53189 587616 60076 587618
rect 53189 587560 53194 587616
rect 53250 587560 60076 587616
rect 173801 587616 180044 587618
rect 53189 587558 60076 587560
rect 53189 587555 53255 587558
rect 134934 587482 134994 587588
rect 173801 587560 173806 587616
rect 173862 587560 180044 587616
rect 173801 587558 180044 587560
rect 254932 587558 284892 587618
rect 173801 587555 173867 587558
rect 284886 587556 284892 587558
rect 284956 587556 284962 587620
rect 288065 587618 288131 587621
rect 377857 587618 377923 587621
rect 288065 587616 300196 587618
rect 288065 587560 288070 587616
rect 288126 587560 300196 587616
rect 288065 587558 300196 587560
rect 374900 587616 377923 587618
rect 374900 587560 377862 587616
rect 377918 587560 377923 587616
rect 374900 587558 377923 587560
rect 288065 587555 288131 587558
rect 377857 587555 377923 587558
rect 174721 587482 174787 587485
rect 134934 587480 174787 587482
rect 134934 587424 174726 587480
rect 174782 587424 174787 587480
rect 134934 587422 174787 587424
rect 174721 587419 174787 587422
rect 134934 586878 142170 586938
rect 134934 586772 134994 586878
rect 142110 586802 142170 586878
rect 172421 586802 172487 586805
rect 291510 586802 291516 586804
rect 142110 586800 172487 586802
rect 142110 586744 172426 586800
rect 172482 586744 172487 586800
rect 142110 586742 172487 586744
rect 254932 586742 291516 586802
rect 172421 586739 172487 586742
rect 291510 586740 291516 586742
rect 291580 586740 291586 586804
rect 377857 586802 377923 586805
rect 374900 586800 377923 586802
rect 374900 586744 377862 586800
rect 377918 586744 377923 586800
rect 374900 586742 377923 586744
rect 377857 586739 377923 586742
rect 59494 586470 60076 586530
rect 179462 586470 180044 586530
rect 299614 586470 300196 586530
rect 54753 586394 54819 586397
rect 59494 586394 59554 586470
rect 54753 586392 59554 586394
rect 54753 586336 54758 586392
rect 54814 586336 59554 586392
rect 54753 586334 59554 586336
rect 172237 586394 172303 586397
rect 179462 586394 179522 586470
rect 172237 586392 179522 586394
rect 172237 586336 172242 586392
rect 172298 586336 179522 586392
rect 172237 586334 179522 586336
rect 287881 586394 287947 586397
rect 299614 586394 299674 586470
rect 287881 586392 299674 586394
rect 287881 586336 287886 586392
rect 287942 586336 299674 586392
rect 287881 586334 299674 586336
rect 54753 586331 54819 586334
rect 172237 586331 172303 586334
rect 287881 586331 287947 586334
rect 176469 585986 176535 585989
rect 295926 585986 295932 585988
rect 142110 585984 176535 585986
rect 134934 585850 134994 585956
rect 142110 585928 176474 585984
rect 176530 585928 176535 585984
rect 142110 585926 176535 585928
rect 254932 585926 295932 585986
rect 142110 585850 142170 585926
rect 176469 585923 176535 585926
rect 295926 585924 295932 585926
rect 295996 585924 296002 585988
rect 377029 585986 377095 585989
rect 374900 585984 377095 585986
rect 374900 585928 377034 585984
rect 377090 585928 377095 585984
rect 374900 585926 377095 585928
rect 377029 585923 377095 585926
rect 134934 585790 142170 585850
rect 54661 585442 54727 585445
rect 166533 585442 166599 585445
rect 175825 585442 175891 585445
rect 288249 585442 288315 585445
rect 54661 585440 60076 585442
rect 54661 585384 54666 585440
rect 54722 585384 60076 585440
rect 54661 585382 60076 585384
rect 166533 585440 180044 585442
rect 166533 585384 166538 585440
rect 166594 585384 175830 585440
rect 175886 585384 180044 585440
rect 166533 585382 180044 585384
rect 288249 585440 300196 585442
rect 288249 585384 288254 585440
rect 288310 585384 300196 585440
rect 288249 585382 300196 585384
rect 54661 585379 54727 585382
rect 166533 585379 166599 585382
rect 175825 585379 175891 585382
rect 288249 585379 288315 585382
rect 144177 585306 144243 585309
rect 145557 585306 145623 585309
rect 134934 585246 142170 585306
rect 134934 585140 134994 585246
rect 142110 585170 142170 585246
rect 144177 585304 145623 585306
rect 144177 585248 144182 585304
rect 144238 585248 145562 585304
rect 145618 585248 145623 585304
rect 144177 585246 145623 585248
rect 144177 585243 144243 585246
rect 145557 585243 145623 585246
rect 179137 585170 179203 585173
rect 289118 585170 289124 585172
rect 142110 585168 179203 585170
rect 142110 585112 179142 585168
rect 179198 585112 179203 585168
rect 142110 585110 179203 585112
rect 254932 585110 289124 585170
rect 179137 585107 179203 585110
rect 289118 585108 289124 585110
rect 289188 585108 289194 585172
rect 295374 585108 295380 585172
rect 295444 585170 295450 585172
rect 296529 585170 296595 585173
rect 377213 585170 377279 585173
rect 295444 585168 296595 585170
rect 295444 585112 296534 585168
rect 296590 585112 296595 585168
rect 295444 585110 296595 585112
rect 374900 585168 377279 585170
rect 374900 585112 377218 585168
rect 377274 585112 377279 585168
rect 374900 585110 377279 585112
rect 295444 585108 295450 585110
rect 296529 585107 296595 585110
rect 377213 585107 377279 585110
rect 54477 584354 54543 584357
rect 286542 584354 286548 584356
rect 54477 584352 60076 584354
rect 54477 584296 54482 584352
rect 54538 584296 60076 584352
rect 54477 584294 60076 584296
rect 54477 584291 54543 584294
rect 134934 584218 134994 584324
rect 176150 584294 180044 584354
rect 254932 584294 286548 584354
rect 176009 584218 176075 584221
rect 134934 584216 176075 584218
rect 134934 584160 176014 584216
rect 176070 584160 176075 584216
rect 134934 584158 176075 584160
rect 176009 584155 176075 584158
rect 169109 583810 169175 583813
rect 174445 583810 174511 583813
rect 176150 583810 176210 584294
rect 286542 584292 286548 584294
rect 286612 584292 286618 584356
rect 290549 584354 290615 584357
rect 377765 584354 377831 584357
rect 290549 584352 300196 584354
rect 290549 584296 290554 584352
rect 290610 584296 300196 584352
rect 290549 584294 300196 584296
rect 374900 584352 377831 584354
rect 374900 584296 377770 584352
rect 377826 584296 377831 584352
rect 374900 584294 377831 584296
rect 290549 584291 290615 584294
rect 377765 584291 377831 584294
rect 169109 583808 176210 583810
rect 169109 583752 169114 583808
rect 169170 583752 174450 583808
rect 174506 583752 176210 583808
rect 169109 583750 176210 583752
rect 169109 583747 169175 583750
rect 174445 583747 174511 583750
rect 285806 583748 285812 583812
rect 285876 583810 285882 583812
rect 286961 583810 287027 583813
rect 285876 583808 287027 583810
rect 285876 583752 286966 583808
rect 287022 583752 287027 583808
rect 285876 583750 287027 583752
rect 285876 583748 285882 583750
rect 286961 583747 287027 583750
rect 178861 583538 178927 583541
rect 283598 583538 283604 583540
rect 142110 583536 178927 583538
rect 134934 583402 134994 583508
rect 142110 583480 178866 583536
rect 178922 583480 178927 583536
rect 142110 583478 178927 583480
rect 254932 583478 283604 583538
rect 142110 583402 142170 583478
rect 178861 583475 178927 583478
rect 283598 583476 283604 583478
rect 283668 583476 283674 583540
rect 378041 583538 378107 583541
rect 374900 583536 378107 583538
rect 374900 583480 378046 583536
rect 378102 583480 378107 583536
rect 374900 583478 378107 583480
rect 378041 583475 378107 583478
rect 134934 583342 142170 583402
rect 55121 583266 55187 583269
rect 290641 583266 290707 583269
rect 55121 583264 60076 583266
rect 55121 583208 55126 583264
rect 55182 583208 60076 583264
rect 55121 583206 60076 583208
rect 176334 583206 180044 583266
rect 290641 583264 300196 583266
rect 290641 583208 290646 583264
rect 290702 583208 300196 583264
rect 290641 583206 300196 583208
rect 55121 583203 55187 583206
rect 176101 582722 176167 582725
rect 142110 582720 176167 582722
rect 134934 582586 134994 582692
rect 142110 582664 176106 582720
rect 176162 582664 176167 582720
rect 142110 582662 176167 582664
rect 142110 582586 142170 582662
rect 176101 582659 176167 582662
rect 134934 582526 142170 582586
rect 169385 582450 169451 582453
rect 176334 582450 176394 583206
rect 290641 583203 290707 583206
rect 403617 582994 403683 582997
rect 427077 582994 427143 582997
rect 403617 582992 427143 582994
rect 403617 582936 403622 582992
rect 403678 582936 427082 582992
rect 427138 582936 427143 582992
rect 403617 582934 427143 582936
rect 403617 582931 403683 582934
rect 427077 582931 427143 582934
rect 271454 582722 271460 582724
rect 254932 582662 271460 582722
rect 271454 582660 271460 582662
rect 271524 582660 271530 582724
rect 378041 582722 378107 582725
rect 374900 582720 378107 582722
rect 374900 582664 378046 582720
rect 378102 582664 378107 582720
rect 374900 582662 378107 582664
rect 378041 582659 378107 582662
rect 169385 582448 176394 582450
rect 169385 582392 169390 582448
rect 169446 582392 176394 582448
rect 169385 582390 176394 582392
rect 169385 582387 169451 582390
rect 51901 582178 51967 582181
rect 166993 582178 167059 582181
rect 168281 582178 168347 582181
rect 279877 582178 279943 582181
rect 51901 582176 60076 582178
rect 51901 582120 51906 582176
rect 51962 582120 60076 582176
rect 51901 582118 60076 582120
rect 166993 582176 180044 582178
rect 166993 582120 166998 582176
rect 167054 582120 168286 582176
rect 168342 582120 180044 582176
rect 166993 582118 180044 582120
rect 279877 582176 300196 582178
rect 279877 582120 279882 582176
rect 279938 582120 300196 582176
rect 279877 582118 300196 582120
rect 51901 582115 51967 582118
rect 166993 582115 167059 582118
rect 168281 582115 168347 582118
rect 279877 582115 279943 582118
rect 173525 581906 173591 581909
rect 290590 581906 290596 581908
rect 142110 581904 173591 581906
rect 134934 581770 134994 581876
rect 142110 581848 173530 581904
rect 173586 581848 173591 581904
rect 142110 581846 173591 581848
rect 254932 581846 290596 581906
rect 142110 581770 142170 581846
rect 173525 581843 173591 581846
rect 290590 581844 290596 581846
rect 290660 581844 290666 581908
rect 382273 581906 382339 581909
rect 374900 581904 382339 581906
rect 374900 581848 382278 581904
rect 382334 581848 382339 581904
rect 374900 581846 382339 581848
rect 382273 581843 382339 581846
rect 134934 581710 142170 581770
rect 174997 581362 175063 581365
rect 134934 581360 175063 581362
rect 134934 581304 175002 581360
rect 175058 581304 175063 581360
rect 134934 581302 175063 581304
rect 54569 581090 54635 581093
rect 54569 581088 60076 581090
rect 54569 581032 54574 581088
rect 54630 581032 60076 581088
rect 134934 581060 134994 581302
rect 174997 581299 175063 581302
rect 157977 581226 158043 581229
rect 166993 581226 167059 581229
rect 157977 581224 167059 581226
rect 157977 581168 157982 581224
rect 158038 581168 166998 581224
rect 167054 581168 167059 581224
rect 157977 581166 167059 581168
rect 157977 581163 158043 581166
rect 166993 581163 167059 581166
rect 159541 581090 159607 581093
rect 179873 581090 179939 581093
rect 274030 581090 274036 581092
rect 159541 581088 180044 581090
rect 54569 581030 60076 581032
rect 159541 581032 159546 581088
rect 159602 581032 179878 581088
rect 179934 581032 180044 581088
rect 159541 581030 180044 581032
rect 254932 581030 274036 581090
rect 54569 581027 54635 581030
rect 159541 581027 159607 581030
rect 179873 581027 179939 581030
rect 274030 581028 274036 581030
rect 274100 581028 274106 581092
rect 282545 581090 282611 581093
rect 378041 581090 378107 581093
rect 282545 581088 300196 581090
rect 282545 581032 282550 581088
rect 282606 581032 300196 581088
rect 282545 581030 300196 581032
rect 374900 581088 378107 581090
rect 374900 581032 378046 581088
rect 378102 581032 378107 581088
rect 374900 581030 378107 581032
rect 282545 581027 282611 581030
rect 378041 581027 378107 581030
rect 179045 580274 179111 580277
rect 292246 580274 292252 580276
rect 142110 580272 179111 580274
rect 134934 580138 134994 580244
rect 142110 580216 179050 580272
rect 179106 580216 179111 580272
rect 142110 580214 179111 580216
rect 254932 580214 292252 580274
rect 142110 580138 142170 580214
rect 179045 580211 179111 580214
rect 292246 580212 292252 580214
rect 292316 580212 292322 580276
rect 378041 580274 378107 580277
rect 374900 580272 378107 580274
rect 374900 580216 378046 580272
rect 378102 580216 378107 580272
rect 374900 580214 378107 580216
rect 378041 580211 378107 580214
rect -960 580002 480 580092
rect 134934 580078 142170 580138
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 49417 580002 49483 580005
rect 282453 580002 282519 580005
rect 49417 580000 60076 580002
rect 49417 579944 49422 580000
rect 49478 579944 60076 580000
rect 49417 579942 60076 579944
rect 171090 579942 180044 580002
rect 282453 580000 300196 580002
rect 282453 579944 282458 580000
rect 282514 579944 300196 580000
rect 282453 579942 300196 579944
rect 49417 579939 49483 579942
rect 158161 579730 158227 579733
rect 168189 579730 168255 579733
rect 171090 579730 171150 579942
rect 282453 579939 282519 579942
rect 158161 579728 171150 579730
rect 158161 579672 158166 579728
rect 158222 579672 168194 579728
rect 168250 579672 171150 579728
rect 158161 579670 171150 579672
rect 158161 579667 158227 579670
rect 168189 579667 168255 579670
rect 291326 579532 291332 579596
rect 291396 579594 291402 579596
rect 292389 579594 292455 579597
rect 291396 579592 292455 579594
rect 291396 579536 292394 579592
rect 292450 579536 292455 579592
rect 291396 579534 292455 579536
rect 291396 579532 291402 579534
rect 292389 579531 292455 579534
rect 176285 579458 176351 579461
rect 290958 579458 290964 579460
rect 142110 579456 176351 579458
rect 134934 579322 134994 579428
rect 142110 579400 176290 579456
rect 176346 579400 176351 579456
rect 142110 579398 176351 579400
rect 254932 579398 290964 579458
rect 142110 579322 142170 579398
rect 176285 579395 176351 579398
rect 290958 579396 290964 579398
rect 291028 579396 291034 579460
rect 377029 579458 377095 579461
rect 374900 579456 377095 579458
rect 374900 579400 377034 579456
rect 377090 579400 377095 579456
rect 374900 579398 377095 579400
rect 377029 579395 377095 579398
rect 134934 579262 142170 579322
rect 51809 578914 51875 578917
rect 169753 578914 169819 578917
rect 170305 578914 170371 578917
rect 282269 578914 282335 578917
rect 51809 578912 60076 578914
rect 51809 578856 51814 578912
rect 51870 578856 60076 578912
rect 51809 578854 60076 578856
rect 169753 578912 180044 578914
rect 169753 578856 169758 578912
rect 169814 578856 170310 578912
rect 170366 578856 180044 578912
rect 169753 578854 180044 578856
rect 282269 578912 300196 578914
rect 282269 578856 282274 578912
rect 282330 578856 300196 578912
rect 282269 578854 300196 578856
rect 51809 578851 51875 578854
rect 169753 578851 169819 578854
rect 170305 578851 170371 578854
rect 282269 578851 282335 578854
rect 178953 578642 179019 578645
rect 291878 578642 291884 578644
rect 142110 578640 179019 578642
rect 134934 578506 134994 578612
rect 142110 578584 178958 578640
rect 179014 578584 179019 578640
rect 142110 578582 179019 578584
rect 254932 578582 291884 578642
rect 142110 578506 142170 578582
rect 178953 578579 179019 578582
rect 291878 578580 291884 578582
rect 291948 578580 291954 578644
rect 378041 578642 378107 578645
rect 374900 578640 378107 578642
rect 374900 578584 378046 578640
rect 378102 578584 378107 578640
rect 374900 578582 378107 578584
rect 378041 578579 378107 578582
rect 134934 578446 142170 578506
rect 158069 578370 158135 578373
rect 169753 578370 169819 578373
rect 158069 578368 169819 578370
rect 158069 578312 158074 578368
rect 158130 578312 169758 578368
rect 169814 578312 169819 578368
rect 158069 578310 169819 578312
rect 158069 578307 158135 578310
rect 169753 578307 169819 578310
rect 427077 578370 427143 578373
rect 431953 578370 432019 578373
rect 427077 578368 432019 578370
rect 427077 578312 427082 578368
rect 427138 578312 431958 578368
rect 432014 578312 432019 578368
rect 427077 578310 432019 578312
rect 427077 578307 427143 578310
rect 431953 578307 432019 578310
rect 290590 578172 290596 578236
rect 290660 578234 290666 578236
rect 291009 578234 291075 578237
rect 290660 578232 291075 578234
rect 290660 578176 291014 578232
rect 291070 578176 291075 578232
rect 290660 578174 291075 578176
rect 290660 578172 290666 578174
rect 291009 578171 291075 578174
rect 291142 578172 291148 578236
rect 291212 578234 291218 578236
rect 292481 578234 292547 578237
rect 291212 578232 292547 578234
rect 291212 578176 292486 578232
rect 292542 578176 292547 578232
rect 291212 578174 292547 578176
rect 291212 578172 291218 578174
rect 292481 578171 292547 578174
rect 49509 577826 49575 577829
rect 172513 577826 172579 577829
rect 282729 577826 282795 577829
rect 379605 577826 379671 577829
rect 49509 577824 60076 577826
rect 49509 577768 49514 577824
rect 49570 577768 60076 577824
rect 172513 577824 180044 577826
rect 49509 577766 60076 577768
rect 49509 577763 49575 577766
rect 134934 577690 134994 577796
rect 172513 577768 172518 577824
rect 172574 577768 180044 577824
rect 282729 577824 300196 577826
rect 172513 577766 180044 577768
rect 172513 577763 172579 577766
rect 178769 577690 178835 577693
rect 134934 577688 178835 577690
rect 134934 577632 178774 577688
rect 178830 577632 178835 577688
rect 134934 577630 178835 577632
rect 254902 577690 254962 577796
rect 282729 577768 282734 577824
rect 282790 577768 300196 577824
rect 282729 577766 300196 577768
rect 374900 577824 379671 577826
rect 374900 577768 379610 577824
rect 379666 577768 379671 577824
rect 374900 577766 379671 577768
rect 282729 577763 282795 577766
rect 379605 577763 379671 577766
rect 291694 577690 291700 577692
rect 254902 577630 291700 577690
rect 178769 577627 178835 577630
rect 291694 577628 291700 577630
rect 291764 577628 291770 577692
rect 548374 577628 548380 577692
rect 548444 577690 548450 577692
rect 583520 577690 584960 577780
rect 548444 577630 584960 577690
rect 548444 577628 548450 577630
rect 583520 577540 584960 577630
rect 290774 577010 290780 577012
rect 134934 576874 134994 576980
rect 254932 576950 290780 577010
rect 290774 576948 290780 576950
rect 290844 576948 290850 577012
rect 381302 577010 381308 577012
rect 374900 576950 381308 577010
rect 381302 576948 381308 576950
rect 381372 576948 381378 577012
rect 137369 576874 137435 576877
rect 134934 576872 137435 576874
rect 134934 576816 137374 576872
rect 137430 576816 137435 576872
rect 134934 576814 137435 576816
rect 137369 576811 137435 576814
rect 158345 576874 158411 576877
rect 172513 576874 172579 576877
rect 158345 576872 172579 576874
rect 158345 576816 158350 576872
rect 158406 576816 172518 576872
rect 172574 576816 172579 576872
rect 158345 576814 172579 576816
rect 158345 576811 158411 576814
rect 172513 576811 172579 576814
rect 47853 576738 47919 576741
rect 175733 576738 175799 576741
rect 282361 576738 282427 576741
rect 47853 576736 60076 576738
rect 47853 576680 47858 576736
rect 47914 576680 60076 576736
rect 47853 576678 60076 576680
rect 175733 576736 180044 576738
rect 175733 576680 175738 576736
rect 175794 576680 180044 576736
rect 175733 576678 180044 576680
rect 282361 576736 300196 576738
rect 282361 576680 282366 576736
rect 282422 576680 300196 576736
rect 282361 576678 300196 576680
rect 47853 576675 47919 576678
rect 175733 576675 175799 576678
rect 282361 576675 282427 576678
rect 173617 576194 173683 576197
rect 295558 576194 295564 576196
rect 142110 576192 173683 576194
rect 134934 576058 134994 576164
rect 142110 576136 173622 576192
rect 173678 576136 173683 576192
rect 142110 576134 173683 576136
rect 254932 576134 295564 576194
rect 142110 576058 142170 576134
rect 173617 576131 173683 576134
rect 295558 576132 295564 576134
rect 295628 576132 295634 576196
rect 377029 576194 377095 576197
rect 374900 576192 377095 576194
rect 374900 576136 377034 576192
rect 377090 576136 377095 576192
rect 374900 576134 377095 576136
rect 377029 576131 377095 576134
rect 134934 575998 142170 576058
rect 50429 575650 50495 575653
rect 161013 575650 161079 575653
rect 170213 575650 170279 575653
rect 282637 575650 282703 575653
rect 50429 575648 60076 575650
rect 50429 575592 50434 575648
rect 50490 575592 60076 575648
rect 50429 575590 60076 575592
rect 161013 575648 180044 575650
rect 161013 575592 161018 575648
rect 161074 575592 170218 575648
rect 170274 575592 180044 575648
rect 161013 575590 180044 575592
rect 282637 575648 300196 575650
rect 282637 575592 282642 575648
rect 282698 575592 300196 575648
rect 282637 575590 300196 575592
rect 50429 575587 50495 575590
rect 161013 575587 161079 575590
rect 170213 575587 170279 575590
rect 282637 575587 282703 575590
rect 158529 575514 158595 575517
rect 175733 575514 175799 575517
rect 176377 575514 176443 575517
rect 158529 575512 176443 575514
rect 158529 575456 158534 575512
rect 158590 575456 175738 575512
rect 175794 575456 176382 575512
rect 176438 575456 176443 575512
rect 158529 575454 176443 575456
rect 158529 575451 158595 575454
rect 175733 575451 175799 575454
rect 176377 575451 176443 575454
rect 295742 575452 295748 575516
rect 295812 575514 295818 575516
rect 296345 575514 296411 575517
rect 295812 575512 296411 575514
rect 295812 575456 296350 575512
rect 296406 575456 296411 575512
rect 295812 575454 296411 575456
rect 295812 575452 295818 575454
rect 296345 575451 296411 575454
rect 166901 575378 166967 575381
rect 256734 575378 256740 575380
rect 142110 575376 166967 575378
rect 134934 575242 134994 575348
rect 142110 575320 166906 575376
rect 166962 575320 166967 575376
rect 142110 575318 166967 575320
rect 254932 575318 256740 575378
rect 142110 575242 142170 575318
rect 166901 575315 166967 575318
rect 256734 575316 256740 575318
rect 256804 575316 256810 575380
rect 376109 575378 376175 575381
rect 374900 575376 376175 575378
rect 374900 575320 376114 575376
rect 376170 575320 376175 575376
rect 374900 575318 376175 575320
rect 376109 575315 376175 575318
rect 134934 575182 142170 575242
rect 51717 574562 51783 574565
rect 164049 574562 164115 574565
rect 179873 574562 179939 574565
rect 285581 574562 285647 574565
rect 378041 574562 378107 574565
rect 51717 574560 60076 574562
rect 51717 574504 51722 574560
rect 51778 574504 60076 574560
rect 164049 574560 180044 574562
rect 51717 574502 60076 574504
rect 51717 574499 51783 574502
rect 134934 574426 134994 574532
rect 164049 574504 164054 574560
rect 164110 574504 179878 574560
rect 179934 574504 180044 574560
rect 285581 574560 300196 574562
rect 164049 574502 180044 574504
rect 164049 574499 164115 574502
rect 179873 574499 179939 574502
rect 168005 574426 168071 574429
rect 134934 574424 168071 574426
rect 134934 574368 168010 574424
rect 168066 574368 168071 574424
rect 134934 574366 168071 574368
rect 254902 574426 254962 574532
rect 285581 574504 285586 574560
rect 285642 574504 300196 574560
rect 285581 574502 300196 574504
rect 374900 574560 378107 574562
rect 374900 574504 378046 574560
rect 378102 574504 378107 574560
rect 374900 574502 378107 574504
rect 285581 574499 285647 574502
rect 378041 574499 378107 574502
rect 292982 574426 292988 574428
rect 254902 574366 292988 574426
rect 168005 574363 168071 574366
rect 292982 574364 292988 574366
rect 293052 574364 293058 574428
rect 256918 574092 256924 574156
rect 256988 574154 256994 574156
rect 257889 574154 257955 574157
rect 256988 574152 257955 574154
rect 256988 574096 257894 574152
rect 257950 574096 257955 574152
rect 256988 574094 257955 574096
rect 256988 574092 256994 574094
rect 257889 574091 257955 574094
rect 292614 574092 292620 574156
rect 292684 574154 292690 574156
rect 293677 574154 293743 574157
rect 292684 574152 293743 574154
rect 292684 574096 293682 574152
rect 293738 574096 293743 574152
rect 292684 574094 293743 574096
rect 292684 574092 292690 574094
rect 293677 574091 293743 574094
rect 292062 573746 292068 573748
rect 53097 573474 53163 573477
rect 53097 573472 60076 573474
rect 53097 573416 53102 573472
rect 53158 573416 60076 573472
rect 53097 573414 60076 573416
rect 53097 573411 53163 573414
rect 134934 573066 134994 573716
rect 254932 573686 292068 573746
rect 292062 573684 292068 573686
rect 292132 573684 292138 573748
rect 376017 573746 376083 573749
rect 374900 573744 376083 573746
rect 374900 573688 376022 573744
rect 376078 573688 376083 573744
rect 374900 573686 376083 573688
rect 376017 573683 376083 573686
rect 166717 573474 166783 573477
rect 179781 573474 179847 573477
rect 288341 573474 288407 573477
rect 166717 573472 180044 573474
rect 166717 573416 166722 573472
rect 166778 573416 179786 573472
rect 179842 573416 180044 573472
rect 166717 573414 180044 573416
rect 288341 573472 300196 573474
rect 288341 573416 288346 573472
rect 288402 573416 300196 573472
rect 288341 573414 300196 573416
rect 166717 573411 166783 573414
rect 179781 573411 179847 573414
rect 288341 573411 288407 573414
rect 134934 573006 135730 573066
rect 135670 572930 135730 573006
rect 277350 573006 292498 573066
rect 137553 572930 137619 572933
rect 169477 572930 169543 572933
rect 277350 572930 277410 573006
rect 135670 572928 137619 572930
rect 134934 572794 134994 572900
rect 135670 572872 137558 572928
rect 137614 572872 137619 572928
rect 135670 572870 137619 572872
rect 137553 572867 137619 572870
rect 142110 572928 169543 572930
rect 142110 572872 169482 572928
rect 169538 572872 169543 572928
rect 142110 572870 169543 572872
rect 254932 572870 277410 572930
rect 142110 572794 142170 572870
rect 169477 572867 169543 572870
rect 291510 572868 291516 572932
rect 291580 572930 291586 572932
rect 292297 572930 292363 572933
rect 292438 572932 292498 573006
rect 291580 572928 292363 572930
rect 291580 572872 292302 572928
rect 292358 572872 292363 572928
rect 291580 572870 292363 572872
rect 291580 572868 291586 572870
rect 292297 572867 292363 572870
rect 292430 572868 292436 572932
rect 292500 572868 292506 572932
rect 377581 572930 377647 572933
rect 374900 572928 377647 572930
rect 374900 572872 377586 572928
rect 377642 572872 377647 572928
rect 374900 572870 377647 572872
rect 377581 572867 377647 572870
rect 292205 572796 292271 572797
rect 292205 572794 292252 572796
rect 134934 572734 142170 572794
rect 292160 572792 292252 572794
rect 292160 572736 292210 572792
rect 292160 572734 292252 572736
rect 292205 572732 292252 572734
rect 292316 572732 292322 572796
rect 431953 572794 432019 572797
rect 435357 572794 435423 572797
rect 431953 572792 435423 572794
rect 431953 572736 431958 572792
rect 432014 572736 435362 572792
rect 435418 572736 435423 572792
rect 431953 572734 435423 572736
rect 292205 572731 292271 572732
rect 431953 572731 432019 572734
rect 435357 572731 435423 572734
rect 54886 572324 54892 572388
rect 54956 572386 54962 572388
rect 178401 572386 178467 572389
rect 290733 572386 290799 572389
rect 54956 572326 60076 572386
rect 178401 572384 180044 572386
rect 178401 572328 178406 572384
rect 178462 572328 180044 572384
rect 178401 572326 180044 572328
rect 290733 572384 300196 572386
rect 290733 572328 290738 572384
rect 290794 572328 300196 572384
rect 290733 572326 300196 572328
rect 54956 572324 54962 572326
rect 178401 572323 178467 572326
rect 290733 572323 290799 572326
rect 172145 572114 172211 572117
rect 294454 572114 294460 572116
rect 142110 572112 172211 572114
rect 134934 571978 134994 572084
rect 142110 572056 172150 572112
rect 172206 572056 172211 572112
rect 142110 572054 172211 572056
rect 254932 572054 294460 572114
rect 142110 571978 142170 572054
rect 172145 572051 172211 572054
rect 294454 572052 294460 572054
rect 294524 572052 294530 572116
rect 383694 572114 383700 572116
rect 374900 572054 383700 572114
rect 383694 572052 383700 572054
rect 383764 572052 383770 572116
rect 134934 571918 142170 571978
rect 294638 571372 294644 571436
rect 294708 571434 294714 571436
rect 295149 571434 295215 571437
rect 294708 571432 295215 571434
rect 294708 571376 295154 571432
rect 295210 571376 295215 571432
rect 294708 571374 295215 571376
rect 294708 571372 294714 571374
rect 295149 571371 295215 571374
rect 58617 571298 58683 571301
rect 175457 571298 175523 571301
rect 277301 571298 277367 571301
rect 379462 571298 379468 571300
rect 58617 571296 60076 571298
rect 58617 571240 58622 571296
rect 58678 571240 60076 571296
rect 142110 571296 175523 571298
rect 58617 571238 60076 571240
rect 58617 571235 58683 571238
rect 134934 571162 134994 571268
rect 142110 571240 175462 571296
rect 175518 571240 175523 571296
rect 142110 571238 175523 571240
rect 142110 571162 142170 571238
rect 175457 571235 175523 571238
rect 175598 571238 180044 571298
rect 277301 571296 300196 571298
rect 134934 571102 142170 571162
rect 169518 571100 169524 571164
rect 169588 571162 169594 571164
rect 175598 571162 175658 571238
rect 169588 571102 175658 571162
rect 254902 571162 254962 571268
rect 277301 571240 277306 571296
rect 277362 571240 300196 571296
rect 277301 571238 300196 571240
rect 374900 571238 379468 571298
rect 277301 571235 277367 571238
rect 379462 571236 379468 571238
rect 379532 571236 379538 571300
rect 299790 571162 299796 571164
rect 254902 571102 299796 571162
rect 169588 571100 169594 571102
rect 299790 571100 299796 571102
rect 299860 571100 299866 571164
rect 161197 570482 161263 570485
rect 299422 570482 299428 570484
rect 142110 570480 161263 570482
rect 134934 570346 134994 570452
rect 142110 570424 161202 570480
rect 161258 570424 161263 570480
rect 142110 570422 161263 570424
rect 254932 570422 299428 570482
rect 142110 570346 142170 570422
rect 161197 570419 161263 570422
rect 299422 570420 299428 570422
rect 299492 570420 299498 570484
rect 382222 570482 382228 570484
rect 374900 570422 382228 570482
rect 382222 570420 382228 570422
rect 382292 570420 382298 570484
rect 134934 570286 142170 570346
rect 55949 570210 56015 570213
rect 55949 570208 60076 570210
rect 55949 570152 55954 570208
rect 56010 570152 60076 570208
rect 55949 570150 60076 570152
rect 55949 570147 56015 570150
rect 171542 570148 171548 570212
rect 171612 570210 171618 570212
rect 171612 570150 180044 570210
rect 171612 570148 171618 570150
rect 281022 570148 281028 570212
rect 281092 570210 281098 570212
rect 281092 570150 300196 570210
rect 281092 570148 281098 570150
rect 299105 570074 299171 570077
rect 299238 570074 299244 570076
rect 299105 570072 299244 570074
rect 299105 570016 299110 570072
rect 299166 570016 299244 570072
rect 299105 570014 299244 570016
rect 299105 570011 299171 570014
rect 299238 570012 299244 570014
rect 299308 570012 299314 570076
rect 299606 570012 299612 570076
rect 299676 570074 299682 570076
rect 299841 570074 299907 570077
rect 299676 570072 299907 570074
rect 299676 570016 299846 570072
rect 299902 570016 299907 570072
rect 299676 570014 299907 570016
rect 299676 570012 299682 570014
rect 299841 570011 299907 570014
rect 142153 569938 142219 569941
rect 144177 569938 144243 569941
rect 142153 569936 144243 569938
rect 142153 569880 142158 569936
rect 142214 569880 144182 569936
rect 144238 569880 144243 569936
rect 142153 569878 144243 569880
rect 142153 569875 142219 569878
rect 144177 569875 144243 569878
rect 177113 569938 177179 569941
rect 177246 569938 177252 569940
rect 177113 569936 177252 569938
rect 177113 569880 177118 569936
rect 177174 569880 177252 569936
rect 177113 569878 177252 569880
rect 177113 569875 177179 569878
rect 177246 569876 177252 569878
rect 177316 569876 177322 569940
rect 170765 569666 170831 569669
rect 295558 569666 295564 569668
rect 142110 569664 170831 569666
rect 134934 569530 134994 569636
rect 142110 569608 170770 569664
rect 170826 569608 170831 569664
rect 142110 569606 170831 569608
rect 254932 569606 295564 569666
rect 142110 569530 142170 569606
rect 170765 569603 170831 569606
rect 295558 569604 295564 569606
rect 295628 569604 295634 569668
rect 377949 569666 378015 569669
rect 374900 569664 378015 569666
rect 374900 569608 377954 569664
rect 378010 569608 378015 569664
rect 374900 569606 378015 569608
rect 377949 569603 378015 569606
rect 134934 569470 142170 569530
rect 59537 569122 59603 569125
rect 59537 569120 60076 569122
rect 59537 569064 59542 569120
rect 59598 569064 60076 569120
rect 59537 569062 60076 569064
rect 59537 569059 59603 569062
rect 177798 569060 177804 569124
rect 177868 569122 177874 569124
rect 297909 569122 297975 569125
rect 177868 569062 180044 569122
rect 297909 569120 300196 569122
rect 297909 569064 297914 569120
rect 297970 569064 300196 569120
rect 297909 569062 300196 569064
rect 177868 569060 177874 569062
rect 297909 569059 297975 569062
rect 134934 568926 142170 568986
rect 134934 568820 134994 568926
rect 142110 568850 142170 568926
rect 163681 568850 163747 568853
rect 288934 568850 288940 568852
rect 142110 568848 163747 568850
rect 142110 568792 163686 568848
rect 163742 568792 163747 568848
rect 142110 568790 163747 568792
rect 254932 568790 288940 568850
rect 163681 568787 163747 568790
rect 288934 568788 288940 568790
rect 289004 568788 289010 568852
rect 379646 568850 379652 568852
rect 374900 568790 379652 568850
rect 379646 568788 379652 568790
rect 379716 568788 379722 568852
rect 296294 568652 296300 568716
rect 296364 568714 296370 568716
rect 296437 568714 296503 568717
rect 296364 568712 296503 568714
rect 296364 568656 296442 568712
rect 296498 568656 296503 568712
rect 296364 568654 296503 568656
rect 296364 568652 296370 568654
rect 296437 568651 296503 568654
rect 56041 568034 56107 568037
rect 56041 568032 60076 568034
rect 56041 567976 56046 568032
rect 56102 567976 60076 568032
rect 56041 567974 60076 567976
rect 56041 567971 56107 567974
rect 173566 567972 173572 568036
rect 173636 568034 173642 568036
rect 296713 568034 296779 568037
rect 173636 567974 180044 568034
rect 296713 568032 300196 568034
rect 296713 567976 296718 568032
rect 296774 567976 300196 568032
rect 296713 567974 300196 567976
rect 173636 567972 173642 567974
rect 296713 567971 296779 567974
rect -960 566946 480 567036
rect 29494 566946 29500 566948
rect -960 566886 29500 566946
rect -960 566796 480 566886
rect 29494 566884 29500 566886
rect 29564 566884 29570 566948
rect 179270 566884 179276 566948
rect 179340 566946 179346 566948
rect 179340 566886 180044 566946
rect 179340 566884 179346 566886
rect 285254 566884 285260 566948
rect 285324 566946 285330 566948
rect 285324 566886 299674 566946
rect 285324 566884 285330 566886
rect 299614 566878 299674 566886
rect 59540 566818 60076 566878
rect 299614 566818 300196 566878
rect 59261 566810 59327 566813
rect 59540 566810 59600 566818
rect 59261 566808 59600 566810
rect 59261 566752 59266 566808
rect 59322 566752 59600 566808
rect 59261 566750 59600 566752
rect 59261 566747 59327 566750
rect 58341 565858 58407 565861
rect 139577 565858 139643 565861
rect 141417 565858 141483 565861
rect 58341 565856 59922 565858
rect 58341 565800 58346 565856
rect 58402 565800 59922 565856
rect 58341 565798 59922 565800
rect 58341 565795 58407 565798
rect 59862 565790 59922 565798
rect 139577 565856 141483 565858
rect 139577 565800 139582 565856
rect 139638 565800 141422 565856
rect 141478 565800 141483 565856
rect 139577 565798 141483 565800
rect 139577 565795 139643 565798
rect 141417 565795 141483 565798
rect 174854 565796 174860 565860
rect 174924 565858 174930 565860
rect 174924 565798 180044 565858
rect 174924 565796 174930 565798
rect 277158 565796 277164 565860
rect 277228 565858 277234 565860
rect 277228 565798 300042 565858
rect 277228 565796 277234 565798
rect 299982 565790 300042 565798
rect 59862 565730 60076 565790
rect 299982 565730 300196 565790
rect 175038 564708 175044 564772
rect 175108 564770 175114 564772
rect 175108 564710 180044 564770
rect 175108 564708 175114 564710
rect 279366 564708 279372 564772
rect 279436 564770 279442 564772
rect 279436 564710 299674 564770
rect 279436 564708 279442 564710
rect 60406 564640 60412 564704
rect 60476 564640 60482 564704
rect 299614 564702 299674 564710
rect 299614 564642 300196 564702
rect 54518 564300 54524 564364
rect 54588 564362 54594 564364
rect 55213 564362 55279 564365
rect 54588 564360 55279 564362
rect 54588 564304 55218 564360
rect 55274 564304 55279 564360
rect 54588 564302 55279 564304
rect 54588 564300 54594 564302
rect 55213 564299 55279 564302
rect 504173 564362 504239 564365
rect 583520 564362 584960 564452
rect 504173 564360 584960 564362
rect 504173 564304 504178 564360
rect 504234 564304 584960 564360
rect 504173 564302 584960 564304
rect 504173 564299 504239 564302
rect 583520 564212 584960 564302
rect 179094 563622 180044 563682
rect 59494 563554 60076 563614
rect 55673 563546 55739 563549
rect 59494 563546 59554 563554
rect 179094 563548 179154 563622
rect 285070 563620 285076 563684
rect 285140 563682 285146 563684
rect 285140 563622 299674 563682
rect 285140 563620 285146 563622
rect 299614 563614 299674 563622
rect 299614 563554 300196 563614
rect 55673 563544 59554 563546
rect 55673 563488 55678 563544
rect 55734 563488 59554 563544
rect 55673 563486 59554 563488
rect 55673 563483 55739 563486
rect 179086 563484 179092 563548
rect 179156 563484 179162 563548
rect 295742 563212 295748 563276
rect 295812 563274 295818 563276
rect 296478 563274 296484 563276
rect 295812 563214 296484 563274
rect 295812 563212 295818 563214
rect 296478 563212 296484 563214
rect 296548 563212 296554 563276
rect 484209 563002 484275 563005
rect 503805 563002 503871 563005
rect 504173 563002 504239 563005
rect 484209 563000 504239 563002
rect 484209 562944 484214 563000
rect 484270 562944 503810 563000
rect 503866 562944 504178 563000
rect 504234 562944 504239 563000
rect 484209 562942 504239 562944
rect 484209 562939 484275 562942
rect 503805 562939 503871 562942
rect 504173 562939 504239 562942
rect 287830 562532 287836 562596
rect 287900 562594 287906 562596
rect 287900 562534 299674 562594
rect 287900 562532 287906 562534
rect 60590 562464 60596 562528
rect 60660 562464 60666 562528
rect 180558 562464 180564 562528
rect 180628 562464 180634 562528
rect 299614 562526 299674 562534
rect 299614 562466 300196 562526
rect 179270 562124 179276 562188
rect 179340 562186 179346 562188
rect 179597 562186 179663 562189
rect 179340 562184 179663 562186
rect 179340 562128 179602 562184
rect 179658 562128 179663 562184
rect 179340 562126 179663 562128
rect 179340 562124 179346 562126
rect 179597 562123 179663 562126
rect 142153 561778 142219 561781
rect 139350 561776 142219 561778
rect 139350 561720 142158 561776
rect 142214 561720 142219 561776
rect 139350 561718 142219 561720
rect 135161 561642 135227 561645
rect 139350 561642 139410 561718
rect 142153 561715 142219 561718
rect 135161 561640 139410 561642
rect 135161 561584 135166 561640
rect 135222 561584 139410 561640
rect 135161 561582 139410 561584
rect 172329 561642 172395 561645
rect 179413 561642 179479 561645
rect 172329 561640 179479 561642
rect 172329 561584 172334 561640
rect 172390 561584 179418 561640
rect 179474 561584 179479 561640
rect 172329 561582 179479 561584
rect 135161 561579 135227 561582
rect 172329 561579 172395 561582
rect 179413 561579 179479 561582
rect 254577 561642 254643 561645
rect 299749 561642 299815 561645
rect 254577 561640 299815 561642
rect 254577 561584 254582 561640
rect 254638 561584 299754 561640
rect 299810 561584 299815 561640
rect 254577 561582 299815 561584
rect 254577 561579 254643 561582
rect 299749 561579 299815 561582
rect 59862 561378 60076 561438
rect 59118 560356 59124 560420
rect 59188 560418 59194 560420
rect 59862 560418 59922 561378
rect 179822 561376 179828 561440
rect 179892 561438 179898 561440
rect 179892 561378 180044 561438
rect 299614 561378 300196 561438
rect 179892 561376 179898 561378
rect 298001 561370 298067 561373
rect 299614 561370 299674 561378
rect 298001 561368 299674 561370
rect 298001 561312 298006 561368
rect 298062 561312 299674 561368
rect 298001 561310 299674 561312
rect 298001 561307 298067 561310
rect 152641 561234 152707 561237
rect 178493 561234 178559 561237
rect 152641 561232 178559 561234
rect 152641 561176 152646 561232
rect 152702 561176 178498 561232
rect 178554 561176 178559 561232
rect 152641 561174 178559 561176
rect 152641 561171 152707 561174
rect 178493 561171 178559 561174
rect 146937 561098 147003 561101
rect 175365 561098 175431 561101
rect 146937 561096 175431 561098
rect 146937 561040 146942 561096
rect 146998 561040 175370 561096
rect 175426 561040 175431 561096
rect 146937 561038 175431 561040
rect 146937 561035 147003 561038
rect 175365 561035 175431 561038
rect 137645 560962 137711 560965
rect 179689 560962 179755 560965
rect 137645 560960 179755 560962
rect 137645 560904 137650 560960
rect 137706 560904 179694 560960
rect 179750 560904 179755 560960
rect 137645 560902 179755 560904
rect 137645 560899 137711 560902
rect 179689 560899 179755 560902
rect 276974 560764 276980 560828
rect 277044 560764 277050 560828
rect 176377 560554 176443 560557
rect 229737 560554 229803 560557
rect 176377 560552 229803 560554
rect 176377 560496 176382 560552
rect 176438 560496 229742 560552
rect 229798 560496 229803 560552
rect 176377 560494 229803 560496
rect 276982 560554 277042 560764
rect 476614 560554 476620 560556
rect 276982 560494 476620 560554
rect 176377 560491 176443 560494
rect 229737 560491 229803 560494
rect 476614 560492 476620 560494
rect 476684 560492 476690 560556
rect 60733 560418 60799 560421
rect 59188 560358 59738 560418
rect 59862 560416 60799 560418
rect 59862 560360 60738 560416
rect 60794 560360 60799 560416
rect 59862 560358 60799 560360
rect 59188 560356 59194 560358
rect 57513 560282 57579 560285
rect 59678 560282 59738 560358
rect 60733 560355 60799 560358
rect 277158 560356 277164 560420
rect 277228 560418 277234 560420
rect 277301 560418 277367 560421
rect 277228 560416 277367 560418
rect 277228 560360 277306 560416
rect 277362 560360 277367 560416
rect 277228 560358 277367 560360
rect 277228 560356 277234 560358
rect 277301 560355 277367 560358
rect 59997 560282 60063 560285
rect 57513 560280 57714 560282
rect 57513 560224 57518 560280
rect 57574 560224 57714 560280
rect 57513 560222 57714 560224
rect 59678 560280 60063 560282
rect 59678 560224 60002 560280
rect 60058 560224 60063 560280
rect 59678 560222 60063 560224
rect 57513 560219 57579 560222
rect 57654 560146 57714 560222
rect 59997 560219 60063 560222
rect 96521 560282 96587 560285
rect 160921 560282 160987 560285
rect 96521 560280 160987 560282
rect 96521 560224 96526 560280
rect 96582 560224 160926 560280
rect 160982 560224 160987 560280
rect 96521 560222 160987 560224
rect 96521 560219 96587 560222
rect 160921 560219 160987 560222
rect 173934 560220 173940 560284
rect 174004 560282 174010 560284
rect 175181 560282 175247 560285
rect 174004 560280 175247 560282
rect 174004 560224 175186 560280
rect 175242 560224 175247 560280
rect 174004 560222 175247 560224
rect 174004 560220 174010 560222
rect 175181 560219 175247 560222
rect 177982 560220 177988 560284
rect 178052 560282 178058 560284
rect 179229 560282 179295 560285
rect 178052 560280 179295 560282
rect 178052 560224 179234 560280
rect 179290 560224 179295 560280
rect 178052 560222 179295 560224
rect 178052 560220 178058 560222
rect 179229 560219 179295 560222
rect 435357 560282 435423 560285
rect 437657 560282 437723 560285
rect 435357 560280 437723 560282
rect 435357 560224 435362 560280
rect 435418 560224 437662 560280
rect 437718 560224 437723 560280
rect 435357 560222 437723 560224
rect 435357 560219 435423 560222
rect 437657 560219 437723 560222
rect 63769 560146 63835 560149
rect 57654 560144 63835 560146
rect 57654 560088 63774 560144
rect 63830 560088 63835 560144
rect 57654 560086 63835 560088
rect 63769 560083 63835 560086
rect 94589 560146 94655 560149
rect 161105 560146 161171 560149
rect 94589 560144 161171 560146
rect 94589 560088 94594 560144
rect 94650 560088 161110 560144
rect 161166 560088 161171 560144
rect 94589 560086 161171 560088
rect 94589 560083 94655 560086
rect 161105 560083 161171 560086
rect 173709 560146 173775 560149
rect 285397 560146 285463 560149
rect 173709 560144 285463 560146
rect 173709 560088 173714 560144
rect 173770 560088 285402 560144
rect 285458 560088 285463 560144
rect 173709 560086 285463 560088
rect 173709 560083 173775 560086
rect 285397 560083 285463 560086
rect 57237 560010 57303 560013
rect 253197 560010 253263 560013
rect 57237 560008 253263 560010
rect 57237 559952 57242 560008
rect 57298 559952 253202 560008
rect 253258 559952 253263 560008
rect 57237 559950 253263 559952
rect 57237 559947 57303 559950
rect 253197 559947 253263 559950
rect 296478 559948 296484 560012
rect 296548 560010 296554 560012
rect 514150 560010 514156 560012
rect 296548 559950 514156 560010
rect 296548 559948 296554 559950
rect 514150 559948 514156 559950
rect 514220 559948 514226 560012
rect 57053 559874 57119 559877
rect 258717 559874 258783 559877
rect 57053 559872 258783 559874
rect 57053 559816 57058 559872
rect 57114 559816 258722 559872
rect 258778 559816 258783 559872
rect 57053 559814 258783 559816
rect 57053 559811 57119 559814
rect 258717 559811 258783 559814
rect 277894 559812 277900 559876
rect 277964 559874 277970 559876
rect 498510 559874 498516 559876
rect 277964 559814 498516 559874
rect 277964 559812 277970 559814
rect 498510 559812 498516 559814
rect 498580 559812 498586 559876
rect 31569 559738 31635 559741
rect 57605 559738 57671 559741
rect 31569 559736 57671 559738
rect 31569 559680 31574 559736
rect 31630 559680 57610 559736
rect 57666 559680 57671 559736
rect 31569 559678 57671 559680
rect 31569 559675 31635 559678
rect 57605 559675 57671 559678
rect 64321 559738 64387 559741
rect 140957 559738 141023 559741
rect 64321 559736 141023 559738
rect 64321 559680 64326 559736
rect 64382 559680 140962 559736
rect 141018 559680 141023 559736
rect 64321 559678 141023 559680
rect 64321 559675 64387 559678
rect 140957 559675 141023 559678
rect 176469 559738 176535 559741
rect 408401 559738 408467 559741
rect 176469 559736 408467 559738
rect 176469 559680 176474 559736
rect 176530 559680 408406 559736
rect 408462 559680 408467 559736
rect 176469 559678 408467 559680
rect 176469 559675 176535 559678
rect 408401 559675 408467 559678
rect 53189 559602 53255 559605
rect 87781 559602 87847 559605
rect 166809 559602 166875 559605
rect 53189 559600 166875 559602
rect 53189 559544 53194 559600
rect 53250 559544 87786 559600
rect 87842 559544 166814 559600
rect 166870 559544 166875 559600
rect 53189 559542 166875 559544
rect 53189 559539 53255 559542
rect 87781 559539 87847 559542
rect 166809 559539 166875 559542
rect 179505 559602 179571 559605
rect 420821 559602 420887 559605
rect 179505 559600 420887 559602
rect 179505 559544 179510 559600
rect 179566 559544 420826 559600
rect 420882 559544 420887 559600
rect 179505 559542 420887 559544
rect 179505 559539 179571 559542
rect 420821 559539 420887 559542
rect 54845 559466 54911 559469
rect 94221 559466 94287 559469
rect 94589 559466 94655 559469
rect 54845 559464 94655 559466
rect 54845 559408 54850 559464
rect 54906 559408 94226 559464
rect 94282 559408 94594 559464
rect 94650 559408 94655 559464
rect 54845 559406 94655 559408
rect 54845 559403 54911 559406
rect 94221 559403 94287 559406
rect 94589 559403 94655 559406
rect 97717 559466 97783 559469
rect 160737 559466 160803 559469
rect 97717 559464 160803 559466
rect 97717 559408 97722 559464
rect 97778 559408 160742 559464
rect 160798 559408 160803 559464
rect 97717 559406 160803 559408
rect 97717 559403 97783 559406
rect 160737 559403 160803 559406
rect 174353 559466 174419 559469
rect 285213 559466 285279 559469
rect 174353 559464 285279 559466
rect 174353 559408 174358 559464
rect 174414 559408 285218 559464
rect 285274 559408 285279 559464
rect 174353 559406 285279 559408
rect 174353 559403 174419 559406
rect 285213 559403 285279 559406
rect 47894 559268 47900 559332
rect 47964 559330 47970 559332
rect 57329 559330 57395 559333
rect 47964 559328 57395 559330
rect 47964 559272 57334 559328
rect 57390 559272 57395 559328
rect 47964 559270 57395 559272
rect 47964 559268 47970 559270
rect 57329 559267 57395 559270
rect 58065 559330 58131 559333
rect 97809 559330 97875 559333
rect 58065 559328 97875 559330
rect 58065 559272 58070 559328
rect 58126 559272 97814 559328
rect 97870 559272 97875 559328
rect 58065 559270 97875 559272
rect 58065 559267 58131 559270
rect 97809 559267 97875 559270
rect 268142 559268 268148 559332
rect 268212 559330 268218 559332
rect 474406 559330 474412 559332
rect 268212 559270 474412 559330
rect 268212 559268 268218 559270
rect 474406 559268 474412 559270
rect 474476 559268 474482 559332
rect 47710 559132 47716 559196
rect 47780 559194 47786 559196
rect 57513 559194 57579 559197
rect 47780 559192 57579 559194
rect 47780 559136 57518 559192
rect 57574 559136 57579 559192
rect 47780 559134 57579 559136
rect 47780 559132 47786 559134
rect 57513 559131 57579 559134
rect 175825 559194 175891 559197
rect 288249 559194 288315 559197
rect 175825 559192 288315 559194
rect 175825 559136 175830 559192
rect 175886 559136 288254 559192
rect 288310 559136 288315 559192
rect 175825 559134 288315 559136
rect 175825 559131 175891 559134
rect 288249 559131 288315 559134
rect 50521 559058 50587 559061
rect 95601 559058 95667 559061
rect 96521 559058 96587 559061
rect 50521 559056 96587 559058
rect 50521 559000 50526 559056
rect 50582 559000 95606 559056
rect 95662 559000 96526 559056
rect 96582 559000 96587 559056
rect 50521 558998 96587 559000
rect 50521 558995 50587 558998
rect 95601 558995 95667 558998
rect 96521 558995 96587 558998
rect 282678 558996 282684 559060
rect 282748 558996 282754 559060
rect 487153 559058 487219 559061
rect 487286 559058 487292 559060
rect 487153 559056 487292 559058
rect 487153 559000 487158 559056
rect 487214 559000 487292 559056
rect 487153 558998 487292 559000
rect 55765 558922 55831 558925
rect 55990 558922 55996 558924
rect 55765 558920 55996 558922
rect 55765 558864 55770 558920
rect 55826 558864 55996 558920
rect 55765 558862 55996 558864
rect 55765 558859 55831 558862
rect 55990 558860 55996 558862
rect 56060 558860 56066 558924
rect 60590 558860 60596 558924
rect 60660 558922 60666 558924
rect 119061 558922 119127 558925
rect 124213 558922 124279 558925
rect 126329 558922 126395 558925
rect 60660 558862 118250 558922
rect 60660 558860 60666 558862
rect 60406 558724 60412 558788
rect 60476 558786 60482 558788
rect 117773 558786 117839 558789
rect 60476 558784 117839 558786
rect 60476 558728 117778 558784
rect 117834 558728 117839 558784
rect 60476 558726 117839 558728
rect 60476 558724 60482 558726
rect 117773 558723 117839 558726
rect 57053 558650 57119 558653
rect 117957 558650 118023 558653
rect 57053 558648 118023 558650
rect 57053 558592 57058 558648
rect 57114 558592 117962 558648
rect 118018 558592 118023 558648
rect 57053 558590 118023 558592
rect 118190 558650 118250 558862
rect 119061 558920 122850 558922
rect 119061 558864 119066 558920
rect 119122 558864 122850 558920
rect 119061 558862 122850 558864
rect 119061 558859 119127 558862
rect 120165 558786 120231 558789
rect 122097 558786 122163 558789
rect 120165 558784 122163 558786
rect 120165 558728 120170 558784
rect 120226 558728 122102 558784
rect 122158 558728 122163 558784
rect 120165 558726 122163 558728
rect 122790 558786 122850 558862
rect 124213 558920 126395 558922
rect 124213 558864 124218 558920
rect 124274 558864 126334 558920
rect 126390 558864 126395 558920
rect 124213 558862 126395 558864
rect 124213 558859 124279 558862
rect 126329 558859 126395 558862
rect 280838 558860 280844 558924
rect 280908 558922 280914 558924
rect 281390 558922 281396 558924
rect 280908 558862 281396 558922
rect 280908 558860 280914 558862
rect 281390 558860 281396 558862
rect 281460 558860 281466 558924
rect 282686 558922 282746 558996
rect 487153 558995 487219 558998
rect 487286 558996 487292 558998
rect 487356 558996 487362 559060
rect 284201 558922 284267 558925
rect 282686 558920 284267 558922
rect 282686 558864 284206 558920
rect 284262 558864 284267 558920
rect 282686 558862 284267 558864
rect 284201 558859 284267 558862
rect 135253 558786 135319 558789
rect 122790 558784 135319 558786
rect 122790 558728 135258 558784
rect 135314 558728 135319 558784
rect 122790 558726 135319 558728
rect 120165 558723 120231 558726
rect 122097 558723 122163 558726
rect 135253 558723 135319 558726
rect 171041 558786 171107 558789
rect 285121 558786 285187 558789
rect 171041 558784 285187 558786
rect 171041 558728 171046 558784
rect 171102 558728 285126 558784
rect 285182 558728 285187 558784
rect 171041 558726 285187 558728
rect 171041 558723 171107 558726
rect 285121 558723 285187 558726
rect 292205 558786 292271 558789
rect 494605 558786 494671 558789
rect 292205 558784 494671 558786
rect 292205 558728 292210 558784
rect 292266 558728 494610 558784
rect 494666 558728 494671 558784
rect 292205 558726 494671 558728
rect 292205 558723 292271 558726
rect 494605 558723 494671 558726
rect 120165 558650 120231 558653
rect 118190 558648 120231 558650
rect 118190 558592 120170 558648
rect 120226 558592 120231 558648
rect 118190 558590 120231 558592
rect 57053 558587 57119 558590
rect 117957 558587 118023 558590
rect 120165 558587 120231 558590
rect 120809 558650 120875 558653
rect 138105 558650 138171 558653
rect 120809 558648 138171 558650
rect 120809 558592 120814 558648
rect 120870 558592 138110 558648
rect 138166 558592 138171 558648
rect 120809 558590 138171 558592
rect 120809 558587 120875 558590
rect 138105 558587 138171 558590
rect 176561 558650 176627 558653
rect 285489 558650 285555 558653
rect 176561 558648 285555 558650
rect 176561 558592 176566 558648
rect 176622 558592 285494 558648
rect 285550 558592 285555 558648
rect 176561 558590 285555 558592
rect 176561 558587 176627 558590
rect 285489 558587 285555 558590
rect 53373 558514 53439 558517
rect 91001 558514 91067 558517
rect 53373 558512 91067 558514
rect 53373 558456 53378 558512
rect 53434 558456 91006 558512
rect 91062 558456 91067 558512
rect 53373 558454 91067 558456
rect 53373 558451 53439 558454
rect 91001 558451 91067 558454
rect 109677 558514 109743 558517
rect 136817 558514 136883 558517
rect 109677 558512 136883 558514
rect 109677 558456 109682 558512
rect 109738 558456 136822 558512
rect 136878 558456 136883 558512
rect 109677 558454 136883 558456
rect 109677 558451 109743 558454
rect 136817 558451 136883 558454
rect 228357 558514 228423 558517
rect 485129 558514 485195 558517
rect 228357 558512 485195 558514
rect 228357 558456 228362 558512
rect 228418 558456 485134 558512
rect 485190 558456 485195 558512
rect 228357 558454 485195 558456
rect 228357 558451 228423 558454
rect 485129 558451 485195 558454
rect 55121 558378 55187 558381
rect 81525 558378 81591 558381
rect 169385 558378 169451 558381
rect 55121 558376 169451 558378
rect 55121 558320 55126 558376
rect 55182 558320 81530 558376
rect 81586 558320 169390 558376
rect 169446 558320 169451 558376
rect 55121 558318 169451 558320
rect 55121 558315 55187 558318
rect 81525 558315 81591 558318
rect 169385 558315 169451 558318
rect 180558 558316 180564 558380
rect 180628 558378 180634 558380
rect 510838 558378 510844 558380
rect 180628 558318 510844 558378
rect 180628 558316 180634 558318
rect 510838 558316 510844 558318
rect 510908 558316 510914 558380
rect 54886 558180 54892 558244
rect 54956 558242 54962 558244
rect 65885 558242 65951 558245
rect 178401 558242 178467 558245
rect 54956 558240 178467 558242
rect 54956 558184 65890 558240
rect 65946 558184 178406 558240
rect 178462 558184 178467 558240
rect 54956 558182 178467 558184
rect 54956 558180 54962 558182
rect 65885 558179 65951 558182
rect 178401 558179 178467 558182
rect 179086 558180 179092 558244
rect 179156 558242 179162 558244
rect 511022 558242 511028 558244
rect 179156 558182 511028 558242
rect 179156 558180 179162 558182
rect 511022 558180 511028 558182
rect 511092 558180 511098 558244
rect 117497 558106 117563 558109
rect 139485 558106 139551 558109
rect 117497 558104 139551 558106
rect 117497 558048 117502 558104
rect 117558 558048 139490 558104
rect 139546 558048 139551 558104
rect 117497 558046 139551 558048
rect 117497 558043 117563 558046
rect 139485 558043 139551 558046
rect 173750 558044 173756 558108
rect 173820 558106 173826 558108
rect 280153 558106 280219 558109
rect 173820 558104 280219 558106
rect 173820 558048 280158 558104
rect 280214 558048 280219 558104
rect 173820 558046 280219 558048
rect 173820 558044 173826 558046
rect 280153 558043 280219 558046
rect 280838 558044 280844 558108
rect 280908 558106 280914 558108
rect 281441 558106 281507 558109
rect 280908 558104 281507 558106
rect 280908 558048 281446 558104
rect 281502 558048 281507 558104
rect 280908 558046 281507 558048
rect 280908 558044 280914 558046
rect 281441 558043 281507 558046
rect 57605 557970 57671 557973
rect 45510 557968 57671 557970
rect 45510 557912 57610 557968
rect 57666 557912 57671 557968
rect 45510 557910 57671 557912
rect 33726 557636 33732 557700
rect 33796 557698 33802 557700
rect 45510 557698 45570 557910
rect 57605 557907 57671 557910
rect 118141 557970 118207 557973
rect 119337 557970 119403 557973
rect 118141 557968 119403 557970
rect 118141 557912 118146 557968
rect 118202 557912 119342 557968
rect 119398 557912 119403 557968
rect 118141 557910 119403 557912
rect 118141 557907 118207 557910
rect 119337 557907 119403 557910
rect 281390 557772 281396 557836
rect 281460 557834 281466 557836
rect 501270 557834 501276 557836
rect 281460 557774 501276 557834
rect 281460 557772 281466 557774
rect 501270 557772 501276 557774
rect 501340 557772 501346 557836
rect 33796 557638 45570 557698
rect 50061 557698 50127 557701
rect 56501 557698 56567 557701
rect 50061 557696 56567 557698
rect 50061 557640 50066 557696
rect 50122 557640 56506 557696
rect 56562 557640 56567 557696
rect 50061 557638 56567 557640
rect 33796 557636 33802 557638
rect 50061 557635 50127 557638
rect 56501 557635 56567 557638
rect 91001 557698 91067 557701
rect 120073 557698 120139 557701
rect 91001 557696 120139 557698
rect 91001 557640 91006 557696
rect 91062 557640 120078 557696
rect 120134 557640 120139 557696
rect 91001 557638 120139 557640
rect 91001 557635 91067 557638
rect 120073 557635 120139 557638
rect 174445 557698 174511 557701
rect 290549 557698 290615 557701
rect 174445 557696 290615 557698
rect 174445 557640 174450 557696
rect 174506 557640 290554 557696
rect 290610 557640 290615 557696
rect 174445 557638 290615 557640
rect 174445 557635 174511 557638
rect 290549 557635 290615 557638
rect 31518 557500 31524 557564
rect 31588 557562 31594 557564
rect 109125 557562 109191 557565
rect 31588 557560 109191 557562
rect 31588 557504 109130 557560
rect 109186 557504 109191 557560
rect 31588 557502 109191 557504
rect 31588 557500 31594 557502
rect 109125 557499 109191 557502
rect 50705 557426 50771 557429
rect 97165 557426 97231 557429
rect 50705 557424 97231 557426
rect 50705 557368 50710 557424
rect 50766 557368 97170 557424
rect 97226 557368 97231 557424
rect 50705 557366 97231 557368
rect 50705 557363 50771 557366
rect 97165 557363 97231 557366
rect 112805 557426 112871 557429
rect 135345 557426 135411 557429
rect 112805 557424 135411 557426
rect 112805 557368 112810 557424
rect 112866 557368 135350 557424
rect 135406 557368 135411 557424
rect 112805 557366 135411 557368
rect 112805 557363 112871 557366
rect 135345 557363 135411 557366
rect 173065 557426 173131 557429
rect 290641 557426 290707 557429
rect 173065 557424 290707 557426
rect 173065 557368 173070 557424
rect 173126 557368 290646 557424
rect 290702 557368 290707 557424
rect 173065 557366 290707 557368
rect 173065 557363 173131 557366
rect 290641 557363 290707 557366
rect 56225 557290 56291 557293
rect 102133 557290 102199 557293
rect 56225 557288 102199 557290
rect 56225 557232 56230 557288
rect 56286 557232 102138 557288
rect 102194 557232 102199 557288
rect 56225 557230 102199 557232
rect 56225 557227 56291 557230
rect 102133 557227 102199 557230
rect 104985 557290 105051 557293
rect 138933 557290 138999 557293
rect 104985 557288 138999 557290
rect 104985 557232 104990 557288
rect 105046 557232 138938 557288
rect 138994 557232 138999 557288
rect 104985 557230 138999 557232
rect 104985 557227 105051 557230
rect 138933 557227 138999 557230
rect 172145 557290 172211 557293
rect 381813 557290 381879 557293
rect 172145 557288 381879 557290
rect 172145 557232 172150 557288
rect 172206 557232 381818 557288
rect 381874 557232 381879 557288
rect 172145 557230 381879 557232
rect 172145 557227 172211 557230
rect 381813 557227 381879 557230
rect 59537 557154 59603 557157
rect 250437 557154 250503 557157
rect 59537 557152 250503 557154
rect 59537 557096 59542 557152
rect 59598 557096 250442 557152
rect 250498 557096 250503 557152
rect 59537 557094 250503 557096
rect 59537 557091 59603 557094
rect 250437 557091 250503 557094
rect 265934 557092 265940 557156
rect 266004 557154 266010 557156
rect 478086 557154 478092 557156
rect 266004 557094 478092 557154
rect 266004 557092 266010 557094
rect 478086 557092 478092 557094
rect 478156 557092 478162 557156
rect 48037 557018 48103 557021
rect 100845 557018 100911 557021
rect 48037 557016 100911 557018
rect 48037 556960 48042 557016
rect 48098 556960 100850 557016
rect 100906 556960 100911 557016
rect 48037 556958 100911 556960
rect 48037 556955 48103 556958
rect 100845 556955 100911 556958
rect 102133 557018 102199 557021
rect 103421 557018 103487 557021
rect 137461 557018 137527 557021
rect 102133 557016 137527 557018
rect 102133 556960 102138 557016
rect 102194 556960 103426 557016
rect 103482 556960 137466 557016
rect 137522 556960 137527 557016
rect 102133 556958 137527 556960
rect 102133 556955 102199 556958
rect 103421 556955 103487 556958
rect 137461 556955 137527 556958
rect 169477 557018 169543 557021
rect 383377 557018 383443 557021
rect 169477 557016 383443 557018
rect 169477 556960 169482 557016
rect 169538 556960 383382 557016
rect 383438 556960 383443 557016
rect 169477 556958 383443 556960
rect 169477 556955 169543 556958
rect 383377 556955 383443 556958
rect 54937 556882 55003 556885
rect 89345 556882 89411 556885
rect 163957 556882 164023 556885
rect 54937 556880 164023 556882
rect 54937 556824 54942 556880
rect 54998 556824 89350 556880
rect 89406 556824 163962 556880
rect 164018 556824 164023 556880
rect 54937 556822 164023 556824
rect 54937 556819 55003 556822
rect 89345 556819 89411 556822
rect 163957 556819 164023 556822
rect 168005 556882 168071 556885
rect 386505 556882 386571 556885
rect 168005 556880 386571 556882
rect 168005 556824 168010 556880
rect 168066 556824 386510 556880
rect 386566 556824 386571 556880
rect 168005 556822 386571 556824
rect 168005 556819 168071 556822
rect 386505 556819 386571 556822
rect 54753 556746 54819 556749
rect 86217 556746 86283 556749
rect 166625 556746 166691 556749
rect 54753 556744 166691 556746
rect 54753 556688 54758 556744
rect 54814 556688 86222 556744
rect 86278 556688 166630 556744
rect 166686 556688 166691 556744
rect 54753 556686 166691 556688
rect 54753 556683 54819 556686
rect 86217 556683 86283 556686
rect 166625 556683 166691 556686
rect 166901 556746 166967 556749
rect 388069 556746 388135 556749
rect 166901 556744 388135 556746
rect 166901 556688 166906 556744
rect 166962 556688 388074 556744
rect 388130 556688 388135 556744
rect 166901 556686 388135 556688
rect 166901 556683 166967 556686
rect 388069 556683 388135 556686
rect 55438 556548 55444 556612
rect 55508 556610 55514 556612
rect 55857 556610 55923 556613
rect 55508 556608 55923 556610
rect 55508 556552 55862 556608
rect 55918 556552 55923 556608
rect 55508 556550 55923 556552
rect 55508 556548 55514 556550
rect 55857 556547 55923 556550
rect 94129 556610 94195 556613
rect 134977 556610 135043 556613
rect 94129 556608 135043 556610
rect 94129 556552 94134 556608
rect 94190 556552 134982 556608
rect 135038 556552 135043 556608
rect 94129 556550 135043 556552
rect 94129 556547 94195 556550
rect 134977 556547 135043 556550
rect 170949 556610 171015 556613
rect 178033 556610 178099 556613
rect 170949 556608 178099 556610
rect 170949 556552 170954 556608
rect 171010 556552 178038 556608
rect 178094 556552 178099 556608
rect 170949 556550 178099 556552
rect 170949 556547 171015 556550
rect 178033 556547 178099 556550
rect 179321 556610 179387 556613
rect 287973 556610 288039 556613
rect 179321 556608 288039 556610
rect 179321 556552 179326 556608
rect 179382 556552 287978 556608
rect 288034 556552 288039 556608
rect 179321 556550 288039 556552
rect 179321 556547 179387 556550
rect 287973 556547 288039 556550
rect 53598 556412 53604 556476
rect 53668 556474 53674 556476
rect 95141 556474 95207 556477
rect 53668 556472 95207 556474
rect 53668 556416 95146 556472
rect 95202 556416 95207 556472
rect 53668 556414 95207 556416
rect 53668 556412 53674 556414
rect 95141 556411 95207 556414
rect 33910 556276 33916 556340
rect 33980 556338 33986 556340
rect 60089 556338 60155 556341
rect 33980 556336 60155 556338
rect 33980 556280 60094 556336
rect 60150 556280 60155 556336
rect 33980 556278 60155 556280
rect 33980 556276 33986 556278
rect 60089 556275 60155 556278
rect 43529 556202 43595 556205
rect 56501 556202 56567 556205
rect 43529 556200 56567 556202
rect 43529 556144 43534 556200
rect 43590 556144 56506 556200
rect 56562 556144 56567 556200
rect 43529 556142 56567 556144
rect 43529 556139 43595 556142
rect 56501 556139 56567 556142
rect 100845 556066 100911 556069
rect 101857 556066 101923 556069
rect 170673 556066 170739 556069
rect 100845 556064 170739 556066
rect 100845 556008 100850 556064
rect 100906 556008 101862 556064
rect 101918 556008 170678 556064
rect 170734 556008 170739 556064
rect 100845 556006 170739 556008
rect 100845 556003 100911 556006
rect 101857 556003 101923 556006
rect 170673 556003 170739 556006
rect 173801 556066 173867 556069
rect 288065 556066 288131 556069
rect 173801 556064 288131 556066
rect 173801 556008 173806 556064
rect 173862 556008 288070 556064
rect 288126 556008 288131 556064
rect 173801 556006 288131 556008
rect 173801 556003 173867 556006
rect 288065 556003 288131 556006
rect 57145 555930 57211 555933
rect 124121 555930 124187 555933
rect 57145 555928 124187 555930
rect 57145 555872 57150 555928
rect 57206 555872 124126 555928
rect 124182 555872 124187 555928
rect 57145 555870 124187 555872
rect 57145 555867 57211 555870
rect 124121 555867 124187 555870
rect 124397 555930 124463 555933
rect 139669 555930 139735 555933
rect 124397 555928 139735 555930
rect 124397 555872 124402 555928
rect 124458 555872 139674 555928
rect 139730 555872 139735 555928
rect 124397 555870 139735 555872
rect 124397 555867 124463 555870
rect 139669 555867 139735 555870
rect 178401 555930 178467 555933
rect 290733 555930 290799 555933
rect 178401 555928 290799 555930
rect 178401 555872 178406 555928
rect 178462 555872 290738 555928
rect 290794 555872 290799 555928
rect 178401 555870 290799 555872
rect 178401 555867 178467 555870
rect 290733 555867 290799 555870
rect 296345 555930 296411 555933
rect 505461 555930 505527 555933
rect 296345 555928 505527 555930
rect 296345 555872 296350 555928
rect 296406 555872 505466 555928
rect 505522 555872 505527 555928
rect 296345 555870 505527 555872
rect 296345 555867 296411 555870
rect 505461 555867 505527 555870
rect 54661 555794 54727 555797
rect 84653 555794 84719 555797
rect 166533 555794 166599 555797
rect 54661 555792 166599 555794
rect 54661 555736 54666 555792
rect 54722 555736 84658 555792
rect 84714 555736 166538 555792
rect 166594 555736 166599 555792
rect 54661 555734 166599 555736
rect 54661 555731 54727 555734
rect 84653 555731 84719 555734
rect 166533 555731 166599 555734
rect 179965 555794 180031 555797
rect 282545 555794 282611 555797
rect 179965 555792 282611 555794
rect 179965 555736 179970 555792
rect 180026 555736 282550 555792
rect 282606 555736 282611 555792
rect 179965 555734 282611 555736
rect 179965 555731 180031 555734
rect 282545 555731 282611 555734
rect 54477 555658 54543 555661
rect 83089 555658 83155 555661
rect 169109 555658 169175 555661
rect 54477 555656 169175 555658
rect 54477 555600 54482 555656
rect 54538 555600 83094 555656
rect 83150 555600 169114 555656
rect 169170 555600 169175 555656
rect 54477 555598 169175 555600
rect 54477 555595 54543 555598
rect 83089 555595 83155 555598
rect 169109 555595 169175 555598
rect 174813 555658 174879 555661
rect 453757 555658 453823 555661
rect 174813 555656 453823 555658
rect 174813 555600 174818 555656
rect 174874 555600 453762 555656
rect 453818 555600 453823 555656
rect 174813 555598 453823 555600
rect 174813 555595 174879 555598
rect 453757 555595 453823 555598
rect 49417 555522 49483 555525
rect 76833 555522 76899 555525
rect 158161 555522 158227 555525
rect 49417 555520 158227 555522
rect 49417 555464 49422 555520
rect 49478 555464 76838 555520
rect 76894 555464 158166 555520
rect 158222 555464 158227 555520
rect 49417 555462 158227 555464
rect 49417 555459 49483 555462
rect 76833 555459 76899 555462
rect 158161 555459 158227 555462
rect 166349 555522 166415 555525
rect 467741 555522 467807 555525
rect 166349 555520 467807 555522
rect 166349 555464 166354 555520
rect 166410 555464 467746 555520
rect 467802 555464 467807 555520
rect 166349 555462 467807 555464
rect 166349 555459 166415 555462
rect 467741 555459 467807 555462
rect 53097 555386 53163 555389
rect 67449 555386 67515 555389
rect 166717 555386 166783 555389
rect 53097 555384 166783 555386
rect 53097 555328 53102 555384
rect 53158 555328 67454 555384
rect 67510 555328 166722 555384
rect 166778 555328 166783 555384
rect 53097 555326 166783 555328
rect 53097 555323 53163 555326
rect 67449 555323 67515 555326
rect 166717 555323 166783 555326
rect 177798 555324 177804 555388
rect 177868 555386 177874 555388
rect 494278 555386 494284 555388
rect 177868 555326 494284 555386
rect 177868 555324 177874 555326
rect 494278 555324 494284 555326
rect 494348 555324 494354 555388
rect 122189 555250 122255 555253
rect 140865 555250 140931 555253
rect 122189 555248 140931 555250
rect 122189 555192 122194 555248
rect 122250 555192 140870 555248
rect 140926 555192 140931 555248
rect 122189 555190 140931 555192
rect 122189 555187 122255 555190
rect 140865 555187 140931 555190
rect 177430 555188 177436 555252
rect 177500 555250 177506 555252
rect 275921 555250 275987 555253
rect 177500 555248 275987 555250
rect 177500 555192 275926 555248
rect 275982 555192 275987 555248
rect 177500 555190 275987 555192
rect 177500 555188 177506 555190
rect 275921 555187 275987 555190
rect 275134 555052 275140 555116
rect 275204 555114 275210 555116
rect 502742 555114 502748 555116
rect 275204 555054 502748 555114
rect 275204 555052 275210 555054
rect 502742 555052 502748 555054
rect 502812 555052 502818 555116
rect 57605 554978 57671 554981
rect 100753 554978 100819 554981
rect 57605 554976 100819 554978
rect 57605 554920 57610 554976
rect 57666 554920 100758 554976
rect 100814 554920 100819 554976
rect 57605 554918 100819 554920
rect 57605 554915 57671 554918
rect 100753 554915 100819 554918
rect 56225 554842 56291 554845
rect 121453 554842 121519 554845
rect 56225 554840 121519 554842
rect 56225 554784 56230 554840
rect 56286 554784 121458 554840
rect 121514 554784 121519 554840
rect 56225 554782 121519 554784
rect 56225 554779 56291 554782
rect 121453 554779 121519 554782
rect 59261 554706 59327 554709
rect 115841 554706 115907 554709
rect 59261 554704 115907 554706
rect 59261 554648 59266 554704
rect 59322 554648 115846 554704
rect 115902 554648 115907 554704
rect 59261 554646 115907 554648
rect 59261 554643 59327 554646
rect 115841 554643 115907 554646
rect 176878 554644 176884 554708
rect 176948 554706 176954 554708
rect 293953 554706 294019 554709
rect 176948 554704 294019 554706
rect 176948 554648 293958 554704
rect 294014 554648 294019 554704
rect 176948 554646 294019 554648
rect 176948 554644 176954 554646
rect 293953 554643 294019 554646
rect 55673 554570 55739 554573
rect 108297 554570 108363 554573
rect 55673 554568 108363 554570
rect 55673 554512 55678 554568
rect 55734 554512 108302 554568
rect 108358 554512 108363 554568
rect 55673 554510 108363 554512
rect 55673 554507 55739 554510
rect 108297 554507 108363 554510
rect 115749 554570 115815 554573
rect 140773 554570 140839 554573
rect 115749 554568 140839 554570
rect 115749 554512 115754 554568
rect 115810 554512 140778 554568
rect 140834 554512 140839 554568
rect 115749 554510 140839 554512
rect 115749 554507 115815 554510
rect 140773 554507 140839 554510
rect 172237 554570 172303 554573
rect 287881 554570 287947 554573
rect 172237 554568 287947 554570
rect 172237 554512 172242 554568
rect 172298 554512 287886 554568
rect 287942 554512 287947 554568
rect 172237 554510 287947 554512
rect 172237 554507 172303 554510
rect 287881 554507 287947 554510
rect 299197 554570 299263 554573
rect 482277 554570 482343 554573
rect 299197 554568 482343 554570
rect 299197 554512 299202 554568
rect 299258 554512 482282 554568
rect 482338 554512 482343 554568
rect 299197 554510 482343 554512
rect 299197 554507 299263 554510
rect 482277 554507 482343 554510
rect 73613 554434 73679 554437
rect 144085 554434 144151 554437
rect 73613 554432 144151 554434
rect 73613 554376 73618 554432
rect 73674 554376 144090 554432
rect 144146 554376 144151 554432
rect 73613 554374 144151 554376
rect 73613 554371 73679 554374
rect 144085 554371 144151 554374
rect 172973 554434 173039 554437
rect 282729 554434 282795 554437
rect 172973 554432 282795 554434
rect 172973 554376 172978 554432
rect 173034 554376 282734 554432
rect 282790 554376 282795 554432
rect 172973 554374 282795 554376
rect 172973 554371 173039 554374
rect 282729 554371 282795 554374
rect 294822 554372 294828 554436
rect 294892 554434 294898 554436
rect 501086 554434 501092 554436
rect 294892 554374 501092 554434
rect 294892 554372 294898 554374
rect 501086 554372 501092 554374
rect 501156 554372 501162 554436
rect 157977 554298 158043 554301
rect 84150 554296 158043 554298
rect 84150 554240 157982 554296
rect 158038 554240 158043 554296
rect 84150 554238 158043 554240
rect 51901 554162 51967 554165
rect 79961 554162 80027 554165
rect 84150 554162 84210 554238
rect 157977 554235 158043 554238
rect 290774 554236 290780 554300
rect 290844 554298 290850 554300
rect 499798 554298 499804 554300
rect 290844 554238 499804 554298
rect 290844 554236 290850 554238
rect 499798 554236 499804 554238
rect 499868 554236 499874 554300
rect 51901 554160 84210 554162
rect 51901 554104 51906 554160
rect 51962 554104 79966 554160
rect 80022 554104 84210 554160
rect 51901 554102 84210 554104
rect 88793 554162 88859 554165
rect 167545 554162 167611 554165
rect 88793 554160 167611 554162
rect 88793 554104 88798 554160
rect 88854 554104 167550 554160
rect 167606 554104 167611 554160
rect 88793 554102 167611 554104
rect 51901 554099 51967 554102
rect 79961 554099 80027 554102
rect 88793 554099 88859 554102
rect 167545 554099 167611 554102
rect 252461 554162 252527 554165
rect 483749 554162 483815 554165
rect 252461 554160 483815 554162
rect 252461 554104 252466 554160
rect 252522 554104 483754 554160
rect 483810 554104 483815 554160
rect 252461 554102 483815 554104
rect 252461 554099 252527 554102
rect 483749 554099 483815 554102
rect 51717 554026 51783 554029
rect 68921 554026 68987 554029
rect 164049 554026 164115 554029
rect 51717 554024 164115 554026
rect -960 553890 480 553980
rect 51717 553968 51722 554024
rect 51778 553968 68926 554024
rect 68982 553968 164054 554024
rect 164110 553968 164115 554024
rect 51717 553966 164115 553968
rect 51717 553963 51783 553966
rect 68921 553963 68987 553966
rect 164049 553963 164115 553966
rect 174854 553964 174860 554028
rect 174924 554026 174930 554028
rect 499614 554026 499620 554028
rect 174924 553966 499620 554026
rect 174924 553964 174930 553966
rect 499614 553964 499620 553966
rect 499684 553964 499690 554028
rect 2814 553890 2820 553892
rect -960 553830 2820 553890
rect -960 553740 480 553830
rect 2814 553828 2820 553830
rect 2884 553828 2890 553892
rect 106549 553890 106615 553893
rect 140037 553890 140103 553893
rect 106549 553888 140103 553890
rect 106549 553832 106554 553888
rect 106610 553832 140042 553888
rect 140098 553832 140103 553888
rect 106549 553830 140103 553832
rect 106549 553827 106615 553830
rect 140037 553827 140103 553830
rect 142797 553890 142863 553893
rect 183185 553890 183251 553893
rect 142797 553888 183251 553890
rect 142797 553832 142802 553888
rect 142858 553832 183190 553888
rect 183246 553832 183251 553888
rect 142797 553830 183251 553832
rect 142797 553827 142863 553830
rect 183185 553827 183251 553830
rect 190913 553890 190979 553893
rect 299289 553890 299355 553893
rect 190913 553888 299355 553890
rect 190913 553832 190918 553888
rect 190974 553832 299294 553888
rect 299350 553832 299355 553888
rect 190913 553830 299355 553832
rect 190913 553827 190979 553830
rect 299289 553827 299355 553830
rect 47393 553754 47459 553757
rect 73153 553754 73219 553757
rect 47393 553752 73219 553754
rect 47393 553696 47398 553752
rect 47454 553696 73158 553752
rect 73214 553696 73219 553752
rect 47393 553694 73219 553696
rect 47393 553691 47459 553694
rect 73153 553691 73219 553694
rect 108113 553754 108179 553757
rect 138841 553754 138907 553757
rect 108113 553752 138907 553754
rect 108113 553696 108118 553752
rect 108174 553696 138846 553752
rect 138902 553696 138907 553752
rect 108113 553694 138907 553696
rect 108113 553691 108179 553694
rect 138841 553691 138907 553694
rect 282177 553754 282243 553757
rect 361481 553754 361547 553757
rect 282177 553752 361547 553754
rect 282177 553696 282182 553752
rect 282238 553696 361486 553752
rect 361542 553696 361547 553752
rect 282177 553694 361547 553696
rect 282177 553691 282243 553694
rect 361481 553691 361547 553694
rect 51901 553618 51967 553621
rect 88977 553618 89043 553621
rect 51901 553616 89043 553618
rect 51901 553560 51906 553616
rect 51962 553560 88982 553616
rect 89038 553560 89043 553616
rect 51901 553558 89043 553560
rect 51901 553555 51967 553558
rect 88977 553555 89043 553558
rect 275461 553618 275527 553621
rect 353661 553618 353727 553621
rect 275461 553616 353727 553618
rect 275461 553560 275466 553616
rect 275522 553560 353666 553616
rect 353722 553560 353727 553616
rect 275461 553558 353727 553560
rect 275461 553555 275527 553558
rect 353661 553555 353727 553558
rect 47526 553420 47532 553484
rect 47596 553482 47602 553484
rect 107561 553482 107627 553485
rect 47596 553480 107627 553482
rect 47596 553424 107566 553480
rect 107622 553424 107627 553480
rect 47596 553422 107627 553424
rect 47596 553420 47602 553422
rect 107561 553419 107627 553422
rect 57646 553284 57652 553348
rect 57716 553346 57722 553348
rect 299289 553346 299355 553349
rect 57716 553344 299355 553346
rect 57716 553288 299294 553344
rect 299350 553288 299355 553344
rect 57716 553286 299355 553288
rect 57716 553284 57722 553286
rect 299289 553283 299355 553286
rect 437657 553346 437723 553349
rect 462221 553346 462287 553349
rect 437657 553344 462287 553346
rect 437657 553288 437662 553344
rect 437718 553288 462226 553344
rect 462282 553288 462287 553344
rect 437657 553286 462287 553288
rect 437657 553283 437723 553286
rect 462221 553283 462287 553286
rect 81709 553210 81775 553213
rect 156597 553210 156663 553213
rect 81709 553208 156663 553210
rect 81709 553152 81714 553208
rect 81770 553152 156602 553208
rect 156658 553152 156663 553208
rect 81709 553150 156663 553152
rect 81709 553147 81775 553150
rect 156597 553147 156663 553150
rect 169753 553210 169819 553213
rect 170990 553210 170996 553212
rect 169753 553208 170996 553210
rect 169753 553152 169758 553208
rect 169814 553152 170996 553208
rect 169753 553150 170996 553152
rect 169753 553147 169819 553150
rect 170990 553148 170996 553150
rect 171060 553148 171066 553212
rect 173566 553148 173572 553212
rect 173636 553210 173642 553212
rect 175825 553210 175891 553213
rect 173636 553208 175891 553210
rect 173636 553152 175830 553208
rect 175886 553152 175891 553208
rect 173636 553150 175891 553152
rect 173636 553148 173642 553150
rect 175825 553147 175891 553150
rect 176193 553210 176259 553213
rect 291745 553210 291811 553213
rect 176193 553208 291811 553210
rect 176193 553152 176198 553208
rect 176254 553152 291750 553208
rect 291806 553152 291811 553208
rect 176193 553150 291811 553152
rect 176193 553147 176259 553150
rect 291745 553147 291811 553150
rect 299289 553210 299355 553213
rect 481766 553210 481772 553212
rect 299289 553208 481772 553210
rect 299289 553152 299294 553208
rect 299350 553152 481772 553208
rect 299289 553150 481772 553152
rect 299289 553147 299355 553150
rect 481766 553148 481772 553150
rect 481836 553148 481842 553212
rect 78397 553074 78463 553077
rect 159541 553074 159607 553077
rect 64830 553072 159607 553074
rect 64830 553016 78402 553072
rect 78458 553016 159546 553072
rect 159602 553016 159607 553072
rect 64830 553014 159607 553016
rect 54569 552938 54635 552941
rect 64830 552938 64890 553014
rect 78397 553011 78463 553014
rect 159541 553011 159607 553014
rect 168189 553074 168255 553077
rect 282453 553074 282519 553077
rect 168189 553072 282519 553074
rect 168189 553016 168194 553072
rect 168250 553016 282458 553072
rect 282514 553016 282519 553072
rect 168189 553014 282519 553016
rect 168189 553011 168255 553014
rect 282453 553011 282519 553014
rect 291878 553012 291884 553076
rect 291948 553074 291954 553076
rect 498326 553074 498332 553076
rect 291948 553014 498332 553074
rect 291948 553012 291954 553014
rect 498326 553012 498332 553014
rect 498396 553012 498402 553076
rect 54569 552936 64890 552938
rect 54569 552880 54574 552936
rect 54630 552880 64890 552936
rect 54569 552878 64890 552880
rect 98913 552938 98979 552941
rect 192569 552938 192635 552941
rect 98913 552936 192635 552938
rect 98913 552880 98918 552936
rect 98974 552880 192574 552936
rect 192630 552880 192635 552936
rect 98913 552878 192635 552880
rect 54569 552875 54635 552878
rect 98913 552875 98979 552878
rect 192569 552875 192635 552878
rect 262806 552876 262812 552940
rect 262876 552938 262882 552940
rect 476062 552938 476068 552940
rect 262876 552878 476068 552938
rect 262876 552876 262882 552878
rect 476062 552876 476068 552878
rect 476132 552876 476138 552940
rect 51809 552802 51875 552805
rect 75269 552802 75335 552805
rect 158069 552802 158135 552805
rect 51809 552800 158135 552802
rect 51809 552744 51814 552800
rect 51870 552744 75274 552800
rect 75330 552744 158074 552800
rect 158130 552744 158135 552800
rect 51809 552742 158135 552744
rect 51809 552739 51875 552742
rect 75269 552739 75335 552742
rect 158069 552739 158135 552742
rect 166758 552740 166764 552804
rect 166828 552802 166834 552804
rect 173801 552802 173867 552805
rect 166828 552800 173867 552802
rect 166828 552744 173806 552800
rect 173862 552744 173867 552800
rect 166828 552742 173867 552744
rect 166828 552740 166834 552742
rect 173801 552739 173867 552742
rect 179781 552802 179847 552805
rect 288341 552802 288407 552805
rect 179781 552800 288407 552802
rect 179781 552744 179786 552800
rect 179842 552744 288346 552800
rect 288402 552744 288407 552800
rect 179781 552742 288407 552744
rect 179781 552739 179847 552742
rect 288341 552739 288407 552742
rect 292430 552740 292436 552804
rect 292500 552802 292506 552804
rect 510654 552802 510660 552804
rect 292500 552742 510660 552802
rect 292500 552740 292506 552742
rect 510654 552740 510660 552742
rect 510724 552740 510730 552804
rect 55949 552666 56015 552669
rect 252001 552666 252067 552669
rect 55949 552664 252067 552666
rect 55949 552608 55954 552664
rect 56010 552608 252006 552664
rect 252062 552608 252067 552664
rect 55949 552606 252067 552608
rect 55949 552603 56015 552606
rect 252001 552603 252067 552606
rect 292062 552604 292068 552668
rect 292132 552666 292138 552668
rect 512126 552666 512132 552668
rect 292132 552606 512132 552666
rect 292132 552604 292138 552606
rect 512126 552604 512132 552606
rect 512196 552604 512202 552668
rect 35433 552530 35499 552533
rect 57789 552530 57855 552533
rect 35433 552528 57855 552530
rect 35433 552472 35438 552528
rect 35494 552472 57794 552528
rect 57850 552472 57855 552528
rect 35433 552470 57855 552472
rect 35433 552467 35499 552470
rect 57789 552467 57855 552470
rect 229369 552530 229435 552533
rect 278681 552530 278747 552533
rect 229369 552528 278747 552530
rect 229369 552472 229374 552528
rect 229430 552472 278686 552528
rect 278742 552472 278747 552528
rect 229369 552470 278747 552472
rect 229369 552467 229435 552470
rect 278681 552467 278747 552470
rect 296110 552468 296116 552532
rect 296180 552530 296186 552532
rect 476798 552530 476804 552532
rect 296180 552470 476804 552530
rect 296180 552468 296186 552470
rect 476798 552468 476804 552470
rect 476868 552468 476874 552532
rect 47945 552394 48011 552397
rect 81433 552394 81499 552397
rect 47945 552392 81499 552394
rect 47945 552336 47950 552392
rect 48006 552336 81438 552392
rect 81494 552336 81499 552392
rect 47945 552334 81499 552336
rect 47945 552331 48011 552334
rect 81433 552331 81499 552334
rect 163589 552394 163655 552397
rect 308305 552394 308371 552397
rect 163589 552392 308371 552394
rect 163589 552336 163594 552392
rect 163650 552336 308310 552392
rect 308366 552336 308371 552392
rect 163589 552334 308371 552336
rect 163589 552331 163655 552334
rect 308305 552331 308371 552334
rect 48037 552258 48103 552261
rect 98637 552258 98703 552261
rect 48037 552256 98703 552258
rect 48037 552200 48042 552256
rect 48098 552200 98642 552256
rect 98698 552200 98703 552256
rect 48037 552198 98703 552200
rect 48037 552195 48103 552198
rect 98637 552195 98703 552198
rect 278313 552258 278379 552261
rect 295333 552258 295399 552261
rect 278313 552256 295399 552258
rect 278313 552200 278318 552256
rect 278374 552200 295338 552256
rect 295394 552200 295399 552256
rect 278313 552198 295399 552200
rect 278313 552195 278379 552198
rect 295333 552195 295399 552198
rect 46606 552060 46612 552124
rect 46676 552122 46682 552124
rect 179413 552122 179479 552125
rect 46676 552120 179479 552122
rect 46676 552064 179418 552120
rect 179474 552064 179479 552120
rect 46676 552062 179479 552064
rect 46676 552060 46682 552062
rect 179413 552059 179479 552062
rect 49509 551986 49575 551989
rect 73705 551986 73771 551989
rect 158345 551986 158411 551989
rect 49509 551984 158411 551986
rect 49509 551928 49514 551984
rect 49570 551928 73710 551984
rect 73766 551928 158350 551984
rect 158406 551928 158411 551984
rect 49509 551926 158411 551928
rect 49509 551923 49575 551926
rect 73705 551923 73771 551926
rect 158345 551923 158411 551926
rect 170213 551986 170279 551989
rect 282637 551986 282703 551989
rect 170213 551984 282703 551986
rect 170213 551928 170218 551984
rect 170274 551928 282642 551984
rect 282698 551928 282703 551984
rect 170213 551926 282703 551928
rect 170213 551923 170279 551926
rect 282637 551923 282703 551926
rect 58525 551850 58591 551853
rect 270769 551850 270835 551853
rect 58525 551848 270835 551850
rect 58525 551792 58530 551848
rect 58586 551792 270774 551848
rect 270830 551792 270835 551848
rect 58525 551790 270835 551792
rect 58525 551787 58591 551790
rect 270769 551787 270835 551790
rect 286317 551850 286383 551853
rect 350441 551850 350507 551853
rect 286317 551848 350507 551850
rect 286317 551792 286322 551848
rect 286378 551792 350446 551848
rect 350502 551792 350507 551848
rect 286317 551790 350507 551792
rect 286317 551787 286383 551790
rect 350441 551787 350507 551790
rect 71773 551714 71839 551717
rect 158529 551714 158595 551717
rect 71773 551712 158595 551714
rect 71773 551656 71778 551712
rect 71834 551656 158534 551712
rect 158590 551656 158595 551712
rect 71773 551654 158595 551656
rect 71773 551651 71839 551654
rect 158529 551651 158595 551654
rect 179137 551714 179203 551717
rect 406837 551714 406903 551717
rect 179137 551712 406903 551714
rect 179137 551656 179142 551712
rect 179198 551656 406842 551712
rect 406898 551656 406903 551712
rect 179137 551654 406903 551656
rect 179137 551651 179203 551654
rect 406837 551651 406903 551654
rect 50429 551578 50495 551581
rect 70577 551578 70643 551581
rect 161013 551578 161079 551581
rect 50429 551576 161079 551578
rect 50429 551520 50434 551576
rect 50490 551520 70582 551576
rect 70638 551520 161018 551576
rect 161074 551520 161079 551576
rect 50429 551518 161079 551520
rect 50429 551515 50495 551518
rect 70577 551515 70643 551518
rect 161013 551515 161079 551518
rect 169518 551516 169524 551580
rect 169588 551578 169594 551580
rect 241421 551578 241487 551581
rect 169588 551576 241487 551578
rect 169588 551520 241426 551576
rect 241482 551520 241487 551576
rect 169588 551518 241487 551520
rect 169588 551516 169594 551518
rect 241421 551515 241487 551518
rect 241605 551578 241671 551581
rect 484393 551578 484459 551581
rect 241605 551576 484459 551578
rect 241605 551520 241610 551576
rect 241666 551520 484398 551576
rect 484454 551520 484459 551576
rect 241605 551518 484459 551520
rect 241605 551515 241671 551518
rect 484393 551515 484459 551518
rect 39757 551442 39823 551445
rect 303245 551442 303311 551445
rect 39757 551440 303311 551442
rect 39757 551384 39762 551440
rect 39818 551384 303250 551440
rect 303306 551384 303311 551440
rect 39757 551382 303311 551384
rect 39757 551379 39823 551382
rect 303245 551379 303311 551382
rect 47853 551306 47919 551309
rect 71773 551306 71839 551309
rect 47853 551304 71839 551306
rect 47853 551248 47858 551304
rect 47914 551248 71778 551304
rect 71834 551248 71839 551304
rect 47853 551246 71839 551248
rect 47853 551243 47919 551246
rect 71773 551243 71839 551246
rect 99925 551306 99991 551309
rect 194133 551306 194199 551309
rect 99925 551304 194199 551306
rect 99925 551248 99930 551304
rect 99986 551248 194138 551304
rect 194194 551248 194199 551304
rect 99925 551246 194199 551248
rect 99925 551243 99991 551246
rect 194133 551243 194199 551246
rect 206093 551306 206159 551309
rect 487705 551306 487771 551309
rect 206093 551304 487771 551306
rect 206093 551248 206098 551304
rect 206154 551248 487710 551304
rect 487766 551248 487771 551304
rect 206093 551246 487771 551248
rect 206093 551243 206159 551246
rect 487705 551243 487771 551246
rect 34329 551170 34395 551173
rect 52453 551170 52519 551173
rect 34329 551168 52519 551170
rect 34329 551112 34334 551168
rect 34390 551112 52458 551168
rect 52514 551112 52519 551168
rect 34329 551110 52519 551112
rect 34329 551107 34395 551110
rect 52453 551107 52519 551110
rect 82721 551170 82787 551173
rect 158161 551170 158227 551173
rect 82721 551168 158227 551170
rect 82721 551112 82726 551168
rect 82782 551112 158166 551168
rect 158222 551112 158227 551168
rect 82721 551110 158227 551112
rect 82721 551107 82787 551110
rect 158161 551107 158227 551110
rect 173249 551170 173315 551173
rect 269113 551170 269179 551173
rect 173249 551168 269179 551170
rect 173249 551112 173254 551168
rect 173310 551112 269118 551168
rect 269174 551112 269179 551168
rect 173249 551110 269179 551112
rect 173249 551107 173315 551110
rect 269113 551107 269179 551110
rect 47761 551034 47827 551037
rect 59261 551034 59327 551037
rect 47761 551032 59327 551034
rect 47761 550976 47766 551032
rect 47822 550976 59266 551032
rect 59322 550976 59327 551032
rect 47761 550974 59327 550976
rect 47761 550971 47827 550974
rect 59261 550971 59327 550974
rect 163998 550972 164004 551036
rect 164068 551034 164074 551036
rect 178033 551034 178099 551037
rect 164068 551032 178099 551034
rect 164068 550976 178038 551032
rect 178094 550976 178099 551032
rect 164068 550974 178099 550976
rect 164068 550972 164074 550974
rect 178033 550971 178099 550974
rect 269798 550972 269804 551036
rect 269868 551034 269874 551036
rect 478270 551034 478276 551036
rect 269868 550974 478276 551034
rect 269868 550972 269874 550974
rect 478270 550972 478276 550974
rect 478340 550972 478346 551036
rect 583520 551020 584960 551260
rect 53097 550898 53163 550901
rect 81433 550898 81499 550901
rect 53097 550896 81499 550898
rect 53097 550840 53102 550896
rect 53158 550840 81438 550896
rect 81494 550840 81499 550896
rect 53097 550838 81499 550840
rect 53097 550835 53163 550838
rect 81433 550835 81499 550838
rect 41086 550700 41092 550764
rect 41156 550762 41162 550764
rect 99373 550762 99439 550765
rect 41156 550760 99439 550762
rect 41156 550704 99378 550760
rect 99434 550704 99439 550760
rect 41156 550702 99439 550704
rect 41156 550700 41162 550702
rect 99373 550699 99439 550702
rect 168281 550626 168347 550629
rect 279877 550626 279943 550629
rect 168281 550624 279943 550626
rect 168281 550568 168286 550624
rect 168342 550568 279882 550624
rect 279938 550568 279943 550624
rect 168281 550566 279943 550568
rect 168281 550563 168347 550566
rect 279877 550563 279943 550566
rect 57513 550490 57579 550493
rect 275553 550490 275619 550493
rect 57513 550488 275619 550490
rect 57513 550432 57518 550488
rect 57574 550432 275558 550488
rect 275614 550432 275619 550488
rect 57513 550430 275619 550432
rect 57513 550427 57579 550430
rect 275553 550427 275619 550430
rect 295057 550490 295123 550493
rect 481725 550490 481791 550493
rect 295057 550488 481791 550490
rect 295057 550432 295062 550488
rect 295118 550432 481730 550488
rect 481786 550432 481791 550488
rect 295057 550430 481791 550432
rect 295057 550427 295123 550430
rect 481725 550427 481791 550430
rect 32990 550292 32996 550356
rect 33060 550354 33066 550356
rect 271270 550354 271276 550356
rect 33060 550294 271276 550354
rect 33060 550292 33066 550294
rect 271270 550292 271276 550294
rect 271340 550292 271346 550356
rect 286542 550292 286548 550356
rect 286612 550354 286618 550356
rect 500902 550354 500908 550356
rect 286612 550294 500908 550354
rect 286612 550292 286618 550294
rect 500902 550292 500908 550294
rect 500972 550292 500978 550356
rect 204805 550218 204871 550221
rect 224953 550218 225019 550221
rect 204805 550216 225019 550218
rect 204805 550160 204810 550216
rect 204866 550160 224958 550216
rect 225014 550160 225019 550216
rect 204805 550158 225019 550160
rect 204805 550155 204871 550158
rect 224953 550155 225019 550158
rect 233049 550218 233115 550221
rect 483197 550218 483263 550221
rect 233049 550216 483263 550218
rect 233049 550160 233054 550216
rect 233110 550160 483202 550216
rect 483258 550160 483263 550216
rect 233049 550158 483263 550160
rect 233049 550155 233115 550158
rect 483197 550155 483263 550158
rect 84745 550082 84811 550085
rect 161289 550082 161355 550085
rect 84745 550080 161355 550082
rect 84745 550024 84750 550080
rect 84806 550024 161294 550080
rect 161350 550024 161355 550080
rect 84745 550022 161355 550024
rect 84745 550019 84811 550022
rect 161289 550019 161355 550022
rect 170581 550082 170647 550085
rect 434989 550082 435055 550085
rect 170581 550080 435055 550082
rect 170581 550024 170586 550080
rect 170642 550024 434994 550080
rect 435050 550024 435055 550080
rect 170581 550022 435055 550024
rect 170581 550019 170647 550022
rect 434989 550019 435055 550022
rect 462221 550082 462287 550085
rect 471605 550082 471671 550085
rect 462221 550080 471671 550082
rect 462221 550024 462226 550080
rect 462282 550024 471610 550080
rect 471666 550024 471671 550080
rect 462221 550022 471671 550024
rect 462221 550019 462287 550022
rect 471605 550019 471671 550022
rect 49509 549946 49575 549949
rect 85481 549946 85547 549949
rect 49509 549944 85547 549946
rect 49509 549888 49514 549944
rect 49570 549888 85486 549944
rect 85542 549888 85547 549944
rect 49509 549886 85547 549888
rect 49509 549883 49575 549886
rect 85481 549883 85547 549886
rect 100937 549946 101003 549949
rect 195697 549946 195763 549949
rect 100937 549944 195763 549946
rect 100937 549888 100942 549944
rect 100998 549888 195702 549944
rect 195758 549888 195763 549944
rect 100937 549886 195763 549888
rect 100937 549883 101003 549886
rect 195697 549883 195763 549886
rect 225045 549946 225111 549949
rect 492121 549946 492187 549949
rect 225045 549944 492187 549946
rect 225045 549888 225050 549944
rect 225106 549888 492126 549944
rect 492182 549888 492187 549944
rect 225045 549886 492187 549888
rect 225045 549883 225111 549886
rect 492121 549883 492187 549886
rect 42425 549810 42491 549813
rect 100753 549810 100819 549813
rect 42425 549808 100819 549810
rect 42425 549752 42430 549808
rect 42486 549752 100758 549808
rect 100814 549752 100819 549808
rect 42425 549750 100819 549752
rect 42425 549747 42491 549750
rect 100753 549747 100819 549750
rect 179873 549810 179939 549813
rect 285581 549810 285647 549813
rect 179873 549808 285647 549810
rect 179873 549752 179878 549808
rect 179934 549752 285586 549808
rect 285642 549752 285647 549808
rect 179873 549750 285647 549752
rect 179873 549747 179939 549750
rect 285581 549747 285647 549750
rect 53189 549674 53255 549677
rect 169753 549674 169819 549677
rect 53189 549672 169819 549674
rect 53189 549616 53194 549672
rect 53250 549616 169758 549672
rect 169814 549616 169819 549672
rect 53189 549614 169819 549616
rect 53189 549611 53255 549614
rect 169753 549611 169819 549614
rect 39430 549476 39436 549540
rect 39500 549538 39506 549540
rect 179413 549538 179479 549541
rect 39500 549536 179479 549538
rect 39500 549480 179418 549536
rect 179474 549480 179479 549536
rect 39500 549478 179479 549480
rect 39500 549476 39506 549478
rect 179413 549475 179479 549478
rect 31150 549340 31156 549404
rect 31220 549402 31226 549404
rect 233141 549402 233207 549405
rect 31220 549400 233207 549402
rect 31220 549344 233146 549400
rect 233202 549344 233207 549400
rect 31220 549342 233207 549344
rect 31220 549340 31226 549342
rect 233141 549339 233207 549342
rect 75637 549266 75703 549269
rect 147213 549266 147279 549269
rect 75637 549264 147279 549266
rect 75637 549208 75642 549264
rect 75698 549208 147218 549264
rect 147274 549208 147279 549264
rect 75637 549206 147279 549208
rect 75637 549203 75703 549206
rect 147213 549203 147279 549206
rect 170305 549266 170371 549269
rect 282269 549266 282335 549269
rect 296294 549266 296300 549268
rect 170305 549264 282335 549266
rect 170305 549208 170310 549264
rect 170366 549208 282274 549264
rect 282330 549208 282335 549264
rect 170305 549206 282335 549208
rect 170305 549203 170371 549206
rect 282269 549203 282335 549206
rect 287010 549206 296300 549266
rect 58341 549130 58407 549133
rect 261385 549130 261451 549133
rect 58341 549128 261451 549130
rect 58341 549072 58346 549128
rect 58402 549072 261390 549128
rect 261446 549072 261451 549128
rect 58341 549070 261451 549072
rect 58341 549067 58407 549070
rect 261385 549067 261451 549070
rect 262857 549130 262923 549133
rect 278681 549130 278747 549133
rect 262857 549128 278747 549130
rect 262857 549072 262862 549128
rect 262918 549072 278686 549128
rect 278742 549072 278747 549128
rect 262857 549070 278747 549072
rect 262857 549067 262923 549070
rect 278681 549067 278747 549070
rect 59118 548932 59124 548996
rect 59188 548994 59194 548996
rect 287010 548994 287070 549206
rect 296294 549204 296300 549206
rect 296364 549204 296370 549268
rect 295742 549068 295748 549132
rect 295812 549130 295818 549132
rect 505134 549130 505140 549132
rect 295812 549070 505140 549130
rect 295812 549068 295818 549070
rect 505134 549068 505140 549070
rect 505204 549068 505210 549132
rect 59188 548934 287070 548994
rect 59188 548932 59194 548934
rect 299054 548932 299060 548996
rect 299124 548994 299130 548996
rect 500166 548994 500172 548996
rect 299124 548934 500172 548994
rect 299124 548932 299130 548934
rect 500166 548932 500172 548934
rect 500236 548932 500242 548996
rect 34278 548796 34284 548860
rect 34348 548858 34354 548860
rect 273846 548858 273852 548860
rect 34348 548798 273852 548858
rect 34348 548796 34354 548798
rect 273846 548796 273852 548798
rect 273916 548796 273922 548860
rect 274030 548796 274036 548860
rect 274100 548858 274106 548860
rect 502374 548858 502380 548860
rect 274100 548798 502380 548858
rect 274100 548796 274106 548798
rect 502374 548796 502380 548798
rect 502444 548796 502450 548860
rect 126329 548722 126395 548725
rect 231669 548722 231735 548725
rect 126329 548720 231735 548722
rect 126329 548664 126334 548720
rect 126390 548664 231674 548720
rect 231730 548664 231735 548720
rect 126329 548662 231735 548664
rect 126329 548659 126395 548662
rect 231669 548659 231735 548662
rect 238201 548722 238267 548725
rect 484485 548722 484551 548725
rect 238201 548720 484551 548722
rect 238201 548664 238206 548720
rect 238262 548664 484490 548720
rect 484546 548664 484551 548720
rect 238201 548662 484551 548664
rect 238201 548659 238267 548662
rect 484485 548659 484551 548662
rect 85757 548586 85823 548589
rect 162761 548586 162827 548589
rect 85757 548584 162827 548586
rect 85757 548528 85762 548584
rect 85818 548528 162766 548584
rect 162822 548528 162827 548584
rect 85757 548526 162827 548528
rect 85757 548523 85823 548526
rect 162761 548523 162827 548526
rect 167913 548586 167979 548589
rect 430297 548586 430363 548589
rect 167913 548584 430363 548586
rect 167913 548528 167918 548584
rect 167974 548528 430302 548584
rect 430358 548528 430363 548584
rect 167913 548526 430363 548528
rect 167913 548523 167979 548526
rect 430297 548523 430363 548526
rect 45001 548450 45067 548453
rect 59261 548450 59327 548453
rect 45001 548448 59327 548450
rect 45001 548392 45006 548448
rect 45062 548392 59266 548448
rect 59322 548392 59327 548448
rect 45001 548390 59327 548392
rect 45001 548387 45067 548390
rect 59261 548387 59327 548390
rect 278221 548450 278287 548453
rect 347405 548450 347471 548453
rect 278221 548448 347471 548450
rect 278221 548392 278226 548448
rect 278282 548392 347410 548448
rect 347466 548392 347471 548448
rect 278221 548390 347471 548392
rect 278221 548387 278287 548390
rect 347405 548387 347471 548390
rect 50705 548314 50771 548317
rect 86861 548314 86927 548317
rect 50705 548312 86927 548314
rect 50705 548256 50710 548312
rect 50766 548256 86866 548312
rect 86922 548256 86927 548312
rect 50705 548254 86927 548256
rect 50705 548251 50771 548254
rect 86861 548251 86927 548254
rect 279601 548314 279667 548317
rect 342713 548314 342779 548317
rect 279601 548312 342779 548314
rect 279601 548256 279606 548312
rect 279662 548256 342718 548312
rect 342774 548256 342779 548312
rect 279601 548254 342779 548256
rect 279601 548251 279667 548254
rect 342713 548251 342779 548254
rect 36629 548178 36695 548181
rect 75821 548178 75887 548181
rect 36629 548176 75887 548178
rect 36629 548120 36634 548176
rect 36690 548120 75826 548176
rect 75882 548120 75887 548176
rect 36629 548118 75887 548120
rect 36629 548115 36695 548118
rect 75821 548115 75887 548118
rect 54753 548042 54819 548045
rect 126881 548042 126947 548045
rect 54753 548040 126947 548042
rect 54753 547984 54758 548040
rect 54814 547984 126886 548040
rect 126942 547984 126947 548040
rect 54753 547982 126947 547984
rect 54753 547979 54819 547982
rect 126881 547979 126947 547982
rect 44081 547906 44147 547909
rect 280061 547906 280127 547909
rect 44081 547904 280127 547906
rect 44081 547848 44086 547904
rect 44142 547848 280066 547904
rect 280122 547848 280127 547904
rect 44081 547846 280127 547848
rect 44081 547843 44147 547846
rect 280061 547843 280127 547846
rect 170254 547708 170260 547772
rect 170324 547770 170330 547772
rect 173801 547770 173867 547773
rect 170324 547768 173867 547770
rect 170324 547712 173806 547768
rect 173862 547712 173867 547768
rect 170324 547710 173867 547712
rect 170324 547708 170330 547710
rect 173801 547707 173867 547710
rect 57830 547572 57836 547636
rect 57900 547634 57906 547636
rect 230381 547634 230447 547637
rect 57900 547632 230447 547634
rect 57900 547576 230386 547632
rect 230442 547576 230447 547632
rect 57900 547574 230447 547576
rect 57900 547572 57906 547574
rect 230381 547571 230447 547574
rect 256734 547572 256740 547636
rect 256804 547634 256810 547636
rect 487470 547634 487476 547636
rect 256804 547574 487476 547634
rect 256804 547572 256810 547574
rect 487470 547572 487476 547574
rect 487540 547572 487546 547636
rect 56041 547498 56107 547501
rect 248873 547498 248939 547501
rect 56041 547496 248939 547498
rect 56041 547440 56046 547496
rect 56102 547440 248878 547496
rect 248934 547440 248939 547496
rect 56041 547438 248939 547440
rect 56041 547435 56107 547438
rect 248873 547435 248939 547438
rect 271454 547436 271460 547500
rect 271524 547498 271530 547500
rect 502558 547498 502564 547500
rect 271524 547438 502564 547498
rect 271524 547436 271530 547438
rect 502558 547436 502564 547438
rect 502628 547436 502634 547500
rect 77661 547362 77727 547365
rect 150341 547362 150407 547365
rect 77661 547360 150407 547362
rect 77661 547304 77666 547360
rect 77722 547304 150346 547360
rect 150402 547304 150407 547360
rect 77661 547302 150407 547304
rect 77661 547299 77727 547302
rect 150341 547299 150407 547302
rect 173433 547362 173499 547365
rect 416221 547362 416287 547365
rect 173433 547360 416287 547362
rect 173433 547304 173438 547360
rect 173494 547304 416226 547360
rect 416282 547304 416287 547360
rect 173433 547302 416287 547304
rect 173433 547299 173499 547302
rect 416221 547299 416287 547302
rect 57421 547226 57487 547229
rect 246389 547226 246455 547229
rect 57421 547224 246455 547226
rect 57421 547168 57426 547224
rect 57482 547168 246394 547224
rect 246450 547168 246455 547224
rect 57421 547166 246455 547168
rect 57421 547163 57487 547166
rect 246389 547163 246455 547166
rect 247401 547226 247467 547229
rect 490373 547226 490439 547229
rect 247401 547224 490439 547226
rect 247401 547168 247406 547224
rect 247462 547168 490378 547224
rect 490434 547168 490439 547224
rect 247401 547166 490439 547168
rect 247401 547163 247467 547166
rect 490373 547163 490439 547166
rect 89805 547090 89871 547093
rect 169109 547090 169175 547093
rect 89805 547088 169175 547090
rect 89805 547032 89810 547088
rect 89866 547032 169114 547088
rect 169170 547032 169175 547088
rect 89805 547030 169175 547032
rect 89805 547027 89871 547030
rect 169109 547027 169175 547030
rect 216949 547090 217015 547093
rect 476941 547090 477007 547093
rect 216949 547088 477007 547090
rect 216949 547032 216954 547088
rect 217010 547032 476946 547088
rect 477002 547032 477007 547088
rect 216949 547030 477007 547032
rect 216949 547027 217015 547030
rect 476941 547027 477007 547030
rect 57329 546954 57395 546957
rect 78581 546954 78647 546957
rect 57329 546952 78647 546954
rect 57329 546896 57334 546952
rect 57390 546896 78586 546952
rect 78642 546896 78647 546952
rect 57329 546894 78647 546896
rect 57329 546891 57395 546894
rect 78581 546891 78647 546894
rect 126237 546954 126303 546957
rect 233877 546954 233943 546957
rect 126237 546952 233943 546954
rect 126237 546896 126242 546952
rect 126298 546896 233882 546952
rect 233938 546896 233943 546952
rect 126237 546894 233943 546896
rect 126237 546891 126303 546894
rect 233877 546891 233943 546894
rect 50521 546818 50587 546821
rect 89713 546818 89779 546821
rect 50521 546816 89779 546818
rect 50521 546760 50526 546816
rect 50582 546760 89718 546816
rect 89774 546760 89779 546816
rect 50521 546758 89779 546760
rect 50521 546755 50587 546758
rect 89713 546755 89779 546758
rect 229737 546818 229803 546821
rect 282361 546818 282427 546821
rect 229737 546816 282427 546818
rect 229737 546760 229742 546816
rect 229798 546760 282366 546816
rect 282422 546760 282427 546816
rect 229737 546758 282427 546760
rect 229737 546755 229803 546758
rect 282361 546755 282427 546758
rect 54845 546682 54911 546685
rect 126881 546682 126947 546685
rect 54845 546680 126947 546682
rect 54845 546624 54850 546680
rect 54906 546624 126886 546680
rect 126942 546624 126947 546680
rect 54845 546622 126947 546624
rect 54845 546619 54911 546622
rect 126881 546619 126947 546622
rect 161197 546682 161263 546685
rect 372245 546682 372311 546685
rect 161197 546680 372311 546682
rect 161197 546624 161202 546680
rect 161258 546624 372250 546680
rect 372306 546624 372311 546680
rect 161197 546622 372311 546624
rect 161197 546619 161263 546622
rect 372245 546619 372311 546622
rect 38469 546546 38535 546549
rect 216673 546546 216739 546549
rect 38469 546544 216739 546546
rect 38469 546488 38474 546544
rect 38530 546488 216678 546544
rect 216734 546488 216739 546544
rect 38469 546486 216739 546488
rect 38469 546483 38535 546486
rect 216673 546483 216739 546486
rect 59670 546348 59676 546412
rect 59740 546410 59746 546412
rect 298921 546410 298987 546413
rect 59740 546408 298987 546410
rect 59740 546352 298926 546408
rect 298982 546352 298987 546408
rect 59740 546350 298987 546352
rect 59740 546348 59746 546350
rect 298921 546347 298987 546350
rect 299105 546410 299171 546413
rect 491937 546410 492003 546413
rect 299105 546408 492003 546410
rect 299105 546352 299110 546408
rect 299166 546352 491942 546408
rect 491998 546352 492003 546408
rect 299105 546350 492003 546352
rect 299105 546347 299171 546350
rect 491937 546347 492003 546350
rect 170857 546274 170923 546277
rect 414657 546274 414723 546277
rect 170857 546272 414723 546274
rect 170857 546216 170862 546272
rect 170918 546216 414662 546272
rect 414718 546216 414723 546272
rect 170857 546214 414723 546216
rect 170857 546211 170923 546214
rect 414657 546211 414723 546214
rect 30230 546076 30236 546140
rect 30300 546138 30306 546140
rect 286358 546138 286364 546140
rect 30300 546078 286364 546138
rect 30300 546076 30306 546078
rect 286358 546076 286364 546078
rect 286428 546076 286434 546140
rect 292982 546076 292988 546140
rect 293052 546138 293058 546140
rect 511206 546138 511212 546140
rect 293052 546078 511212 546138
rect 293052 546076 293058 546078
rect 511206 546076 511212 546078
rect 511276 546076 511282 546140
rect 51809 546002 51875 546005
rect 309593 546002 309659 546005
rect 51809 546000 309659 546002
rect 51809 545944 51814 546000
rect 51870 545944 309598 546000
rect 309654 545944 309659 546000
rect 51809 545942 309659 545944
rect 51809 545939 51875 545942
rect 309593 545939 309659 545942
rect 59670 545804 59676 545868
rect 59740 545866 59746 545868
rect 60365 545866 60431 545869
rect 59740 545864 60431 545866
rect 59740 545808 60370 545864
rect 60426 545808 60431 545864
rect 59740 545806 60431 545808
rect 59740 545804 59746 545806
rect 60365 545803 60431 545806
rect 90817 545866 90883 545869
rect 170673 545866 170739 545869
rect 90817 545864 170739 545866
rect 90817 545808 90822 545864
rect 90878 545808 170678 545864
rect 170734 545808 170739 545864
rect 90817 545806 170739 545808
rect 90817 545803 90883 545806
rect 170673 545803 170739 545806
rect 223021 545866 223087 545869
rect 483841 545866 483907 545869
rect 223021 545864 483907 545866
rect 223021 545808 223026 545864
rect 223082 545808 483846 545864
rect 483902 545808 483907 545864
rect 223021 545806 483907 545808
rect 223021 545803 223087 545806
rect 483841 545803 483907 545806
rect 34237 545730 34303 545733
rect 60181 545730 60247 545733
rect 34237 545728 60247 545730
rect 34237 545672 34242 545728
rect 34298 545672 60186 545728
rect 60242 545672 60247 545728
rect 34237 545670 60247 545672
rect 34237 545667 34303 545670
rect 60181 545667 60247 545670
rect 78673 545730 78739 545733
rect 151905 545730 151971 545733
rect 78673 545728 151971 545730
rect 78673 545672 78678 545728
rect 78734 545672 151910 545728
rect 151966 545672 151971 545728
rect 78673 545670 151971 545672
rect 78673 545667 78739 545670
rect 151905 545667 151971 545670
rect 169293 545730 169359 545733
rect 452193 545730 452259 545733
rect 169293 545728 452259 545730
rect 169293 545672 169298 545728
rect 169354 545672 452198 545728
rect 452254 545672 452259 545728
rect 169293 545670 452259 545672
rect 169293 545667 169359 545670
rect 452193 545667 452259 545670
rect 49417 545594 49483 545597
rect 79317 545594 79383 545597
rect 49417 545592 79383 545594
rect 49417 545536 49422 545592
rect 49478 545536 79322 545592
rect 79378 545536 79383 545592
rect 49417 545534 79383 545536
rect 49417 545531 49483 545534
rect 79317 545531 79383 545534
rect 122281 545594 122347 545597
rect 228541 545594 228607 545597
rect 122281 545592 228607 545594
rect 122281 545536 122286 545592
rect 122342 545536 228546 545592
rect 228602 545536 228607 545592
rect 122281 545534 228607 545536
rect 122281 545531 122347 545534
rect 228541 545531 228607 545534
rect 289118 545532 289124 545596
rect 289188 545594 289194 545596
rect 498694 545594 498700 545596
rect 289188 545534 498700 545594
rect 289188 545532 289194 545534
rect 498694 545532 498700 545534
rect 498764 545532 498770 545596
rect 35341 545458 35407 545461
rect 89713 545458 89779 545461
rect 35341 545456 89779 545458
rect 35341 545400 35346 545456
rect 35402 545400 89718 545456
rect 89774 545400 89779 545456
rect 35341 545398 89779 545400
rect 35341 545395 35407 545398
rect 89713 545395 89779 545398
rect 41045 545322 41111 545325
rect 121453 545322 121519 545325
rect 41045 545320 121519 545322
rect 41045 545264 41050 545320
rect 41106 545264 121458 545320
rect 121514 545264 121519 545320
rect 41045 545262 121519 545264
rect 41045 545259 41111 545262
rect 121453 545259 121519 545262
rect 38193 545186 38259 545189
rect 223481 545186 223547 545189
rect 38193 545184 223547 545186
rect 38193 545128 38198 545184
rect 38254 545128 223486 545184
rect 223542 545128 223547 545184
rect 38193 545126 223547 545128
rect 38193 545123 38259 545126
rect 223481 545123 223547 545126
rect 485773 545186 485839 545189
rect 486366 545186 486372 545188
rect 485773 545184 486372 545186
rect 485773 545128 485778 545184
rect 485834 545128 486372 545184
rect 485773 545126 486372 545128
rect 485773 545123 485839 545126
rect 486366 545124 486372 545126
rect 486436 545124 486442 545188
rect 159449 545050 159515 545053
rect 323945 545050 324011 545053
rect 159449 545048 324011 545050
rect 159449 544992 159454 545048
rect 159510 544992 323950 545048
rect 324006 544992 324011 545048
rect 159449 544990 324011 544992
rect 159449 544987 159515 544990
rect 323945 544987 324011 544990
rect 79685 544914 79751 544917
rect 153469 544914 153535 544917
rect 79685 544912 153535 544914
rect 79685 544856 79690 544912
rect 79746 544856 153474 544912
rect 153530 544856 153535 544912
rect 79685 544854 153535 544856
rect 79685 544851 79751 544854
rect 153469 544851 153535 544854
rect 171961 544914 172027 544917
rect 175273 544914 175339 544917
rect 171961 544912 175339 544914
rect 171961 544856 171966 544912
rect 172022 544856 175278 544912
rect 175334 544856 175339 544912
rect 171961 544854 175339 544856
rect 171961 544851 172027 544854
rect 175273 544851 175339 544854
rect 175733 544914 175799 544917
rect 380249 544914 380315 544917
rect 175733 544912 380315 544914
rect 175733 544856 175738 544912
rect 175794 544856 380254 544912
rect 380310 544856 380315 544912
rect 175733 544854 380315 544856
rect 175733 544851 175799 544854
rect 380249 544851 380315 544854
rect 58709 544778 58775 544781
rect 273897 544778 273963 544781
rect 58709 544776 273963 544778
rect 58709 544720 58714 544776
rect 58770 544720 273902 544776
rect 273958 544720 273963 544776
rect 58709 544718 273963 544720
rect 58709 544715 58775 544718
rect 273897 544715 273963 544718
rect 276749 544778 276815 544781
rect 345841 544778 345907 544781
rect 276749 544776 345907 544778
rect 276749 544720 276754 544776
rect 276810 544720 345846 544776
rect 345902 544720 345907 544776
rect 276749 544718 345907 544720
rect 276749 544715 276815 544718
rect 345841 544715 345907 544718
rect 128169 544642 128235 544645
rect 237925 544642 237991 544645
rect 128169 544640 237991 544642
rect 128169 544584 128174 544640
rect 128230 544584 237930 544640
rect 237986 544584 237991 544640
rect 128169 544582 237991 544584
rect 128169 544579 128235 544582
rect 237925 544579 237991 544582
rect 249333 544642 249399 544645
rect 486325 544642 486391 544645
rect 249333 544640 486391 544642
rect 249333 544584 249338 544640
rect 249394 544584 486330 544640
rect 486386 544584 486391 544640
rect 249333 544582 486391 544584
rect 249333 544579 249399 544582
rect 486325 544579 486391 544582
rect 92841 544506 92907 544509
rect 173709 544506 173775 544509
rect 92841 544504 173775 544506
rect 92841 544448 92846 544504
rect 92902 544448 173714 544504
rect 173770 544448 173775 544504
rect 92841 544446 173775 544448
rect 92841 544443 92907 544446
rect 173709 544443 173775 544446
rect 174905 544506 174971 544509
rect 417785 544506 417851 544509
rect 174905 544504 417851 544506
rect 174905 544448 174910 544504
rect 174966 544448 417790 544504
rect 417846 544448 417851 544504
rect 174905 544446 417851 544448
rect 174905 544443 174971 544446
rect 417785 544443 417851 544446
rect 31334 544308 31340 544372
rect 31404 544370 31410 544372
rect 277158 544370 277164 544372
rect 31404 544310 277164 544370
rect 31404 544308 31410 544310
rect 277158 544308 277164 544310
rect 277228 544308 277234 544372
rect 295006 544308 295012 544372
rect 295076 544370 295082 544372
rect 506606 544370 506612 544372
rect 295076 544310 506612 544370
rect 295076 544308 295082 544310
rect 506606 544308 506612 544310
rect 506676 544308 506682 544372
rect 43846 544172 43852 544236
rect 43916 544234 43922 544236
rect 92473 544234 92539 544237
rect 43916 544232 92539 544234
rect 43916 544176 92478 544232
rect 92534 544176 92539 544232
rect 43916 544174 92539 544176
rect 43916 544172 43922 544174
rect 92473 544171 92539 544174
rect 152549 544234 152615 544237
rect 293953 544234 294019 544237
rect 152549 544232 294019 544234
rect 152549 544176 152554 544232
rect 152610 544176 293958 544232
rect 294014 544176 294019 544232
rect 152549 544174 294019 544176
rect 152549 544171 152615 544174
rect 293953 544171 294019 544174
rect 49141 544098 49207 544101
rect 127617 544098 127683 544101
rect 49141 544096 127683 544098
rect 49141 544040 49146 544096
rect 49202 544040 127622 544096
rect 127678 544040 127683 544096
rect 49141 544038 127683 544040
rect 49141 544035 49207 544038
rect 127617 544035 127683 544038
rect 289261 544098 289327 544101
rect 344277 544098 344343 544101
rect 289261 544096 344343 544098
rect 289261 544040 289266 544096
rect 289322 544040 344282 544096
rect 344338 544040 344343 544096
rect 289261 544038 344343 544040
rect 289261 544035 289327 544038
rect 344277 544035 344343 544038
rect 41229 543962 41295 543965
rect 153101 543962 153167 543965
rect 41229 543960 153167 543962
rect 41229 543904 41234 543960
rect 41290 543904 153106 543960
rect 153162 543904 153167 543960
rect 41229 543902 153167 543904
rect 41229 543899 41295 543902
rect 153101 543899 153167 543902
rect 54937 543826 55003 543829
rect 172421 543826 172487 543829
rect 54937 543824 172487 543826
rect 54937 543768 54942 543824
rect 54998 543768 172426 543824
rect 172482 543768 172487 543824
rect 54937 543766 172487 543768
rect 54937 543763 55003 543766
rect 172421 543763 172487 543766
rect 57697 543690 57763 543693
rect 269757 543690 269823 543693
rect 57697 543688 269823 543690
rect 57697 543632 57702 543688
rect 57758 543632 269762 543688
rect 269818 543632 269823 543688
rect 57697 543630 269823 543632
rect 57697 543627 57763 543630
rect 269757 543627 269823 543630
rect 72601 543554 72667 543557
rect 142521 543554 142587 543557
rect 72601 543552 142587 543554
rect 72601 543496 72606 543552
rect 72662 543496 142526 543552
rect 142582 543496 142587 543552
rect 72601 543494 142587 543496
rect 72601 543491 72667 543494
rect 142521 543491 142587 543494
rect 173525 543554 173591 543557
rect 400581 543554 400647 543557
rect 173525 543552 400647 543554
rect 173525 543496 173530 543552
rect 173586 543496 400586 543552
rect 400642 543496 400647 543552
rect 173525 543494 400647 543496
rect 173525 543491 173591 543494
rect 400581 543491 400647 543494
rect 58433 543418 58499 543421
rect 287973 543418 288039 543421
rect 58433 543416 288039 543418
rect 58433 543360 58438 543416
rect 58494 543360 287978 543416
rect 288034 543360 288039 543416
rect 58433 543358 288039 543360
rect 58433 543355 58499 543358
rect 287973 543355 288039 543358
rect 293166 543356 293172 543420
rect 293236 543418 293242 543420
rect 481950 543418 481956 543420
rect 293236 543358 481956 543418
rect 293236 543356 293242 543358
rect 481950 543356 481956 543358
rect 482020 543356 482026 543420
rect 125225 543282 125291 543285
rect 231209 543282 231275 543285
rect 125225 543280 231275 543282
rect 125225 543224 125230 543280
rect 125286 543224 231214 543280
rect 231270 543224 231275 543280
rect 125225 543222 231275 543224
rect 125225 543219 125291 543222
rect 231209 543219 231275 543222
rect 237189 543282 237255 543285
rect 484577 543282 484643 543285
rect 237189 543280 484643 543282
rect 237189 543224 237194 543280
rect 237250 543224 484582 543280
rect 484638 543224 484643 543280
rect 237189 543222 484643 543224
rect 237189 543219 237255 543222
rect 484577 543219 484643 543222
rect 94865 543146 94931 543149
rect 187877 543146 187943 543149
rect 94865 543144 187943 543146
rect 94865 543088 94870 543144
rect 94926 543088 187882 543144
rect 187938 543088 187943 543144
rect 94865 543086 187943 543088
rect 94865 543083 94931 543086
rect 187877 543083 187943 543086
rect 200757 543146 200823 543149
rect 230381 543146 230447 543149
rect 200757 543144 230447 543146
rect 200757 543088 200762 543144
rect 200818 543088 230386 543144
rect 230442 543088 230447 543144
rect 200757 543086 230447 543088
rect 200757 543083 200823 543086
rect 230381 543083 230447 543086
rect 230657 543146 230723 543149
rect 490281 543146 490347 543149
rect 230657 543144 490347 543146
rect 230657 543088 230662 543144
rect 230718 543088 490286 543144
rect 490342 543088 490347 543144
rect 230657 543086 490347 543088
rect 230657 543083 230723 543086
rect 490281 543083 490347 543086
rect 87873 543010 87939 543013
rect 165981 543010 166047 543013
rect 87873 543008 166047 543010
rect 87873 542952 87878 543008
rect 87934 542952 165986 543008
rect 166042 542952 166047 543008
rect 87873 542950 166047 542952
rect 87873 542947 87939 542950
rect 165981 542947 166047 542950
rect 167637 543010 167703 543013
rect 172513 543010 172579 543013
rect 167637 543008 172579 543010
rect 167637 542952 167642 543008
rect 167698 542952 172518 543008
rect 172574 542952 172579 543008
rect 167637 542950 172579 542952
rect 167637 542947 167703 542950
rect 172513 542947 172579 542950
rect 175958 542948 175964 543012
rect 176028 543010 176034 543012
rect 444281 543010 444347 543013
rect 176028 543008 444347 543010
rect 176028 542952 444286 543008
rect 444342 542952 444347 543008
rect 176028 542950 444347 542952
rect 176028 542948 176034 542950
rect 444281 542947 444347 542950
rect 155401 542874 155467 542877
rect 339585 542874 339651 542877
rect 155401 542872 339651 542874
rect 155401 542816 155406 542872
rect 155462 542816 339590 542872
rect 339646 542816 339651 542872
rect 155401 542814 339651 542816
rect 155401 542811 155467 542814
rect 339585 542811 339651 542814
rect 48865 542738 48931 542741
rect 95141 542738 95207 542741
rect 48865 542736 95207 542738
rect 48865 542680 48870 542736
rect 48926 542680 95146 542736
rect 95202 542680 95207 542736
rect 48865 542678 95207 542680
rect 48865 542675 48931 542678
rect 95141 542675 95207 542678
rect 54661 542602 54727 542605
rect 125501 542602 125567 542605
rect 54661 542600 125567 542602
rect 54661 542544 54666 542600
rect 54722 542544 125506 542600
rect 125562 542544 125567 542600
rect 54661 542542 125567 542544
rect 54661 542539 54727 542542
rect 125501 542539 125567 542542
rect 39665 542466 39731 542469
rect 175273 542466 175339 542469
rect 39665 542464 175339 542466
rect 39665 542408 39670 542464
rect 39726 542408 175278 542464
rect 175334 542408 175339 542464
rect 39665 542406 175339 542408
rect 39665 542403 39731 542406
rect 175273 542403 175339 542406
rect 49601 542330 49667 542333
rect 284845 542330 284911 542333
rect 49601 542328 284911 542330
rect 49601 542272 49606 542328
rect 49662 542272 284850 542328
rect 284906 542272 284911 542328
rect 49601 542270 284911 542272
rect 49601 542267 49667 542270
rect 284845 542267 284911 542270
rect 293677 542330 293743 542333
rect 481817 542330 481883 542333
rect 293677 542328 481883 542330
rect 293677 542272 293682 542328
rect 293738 542272 481822 542328
rect 481878 542272 481883 542328
rect 293677 542270 481883 542272
rect 293677 542267 293743 542270
rect 481817 542267 481883 542270
rect 173341 542194 173407 542197
rect 413093 542194 413159 542197
rect 173341 542192 413159 542194
rect 173341 542136 173346 542192
rect 173402 542136 413098 542192
rect 413154 542136 413159 542192
rect 173341 542134 413159 542136
rect 173341 542131 173407 542134
rect 413093 542131 413159 542134
rect 56317 542058 56383 542061
rect 302049 542058 302115 542061
rect 56317 542056 302115 542058
rect 56317 542000 56322 542056
rect 56378 542000 302054 542056
rect 302110 542000 302115 542056
rect 56317 541998 302115 542000
rect 56317 541995 56383 541998
rect 302049 541995 302115 541998
rect 232129 541922 232195 541925
rect 483289 541922 483355 541925
rect 232129 541920 483355 541922
rect 232129 541864 232134 541920
rect 232190 541864 483294 541920
rect 483350 541864 483355 541920
rect 232129 541862 483355 541864
rect 232129 541859 232195 541862
rect 483289 541859 483355 541862
rect 113081 541786 113147 541789
rect 214465 541786 214531 541789
rect 113081 541784 214531 541786
rect 113081 541728 113086 541784
rect 113142 541728 214470 541784
rect 214526 541728 214531 541784
rect 113081 541726 214531 541728
rect 113081 541723 113147 541726
rect 214465 541723 214531 541726
rect 224033 541786 224099 541789
rect 486233 541786 486299 541789
rect 224033 541784 486299 541786
rect 224033 541728 224038 541784
rect 224094 541728 486238 541784
rect 486294 541728 486299 541784
rect 224033 541726 486299 541728
rect 224033 541723 224099 541726
rect 486233 541723 486299 541726
rect 76649 541650 76715 541653
rect 148777 541650 148843 541653
rect 76649 541648 148843 541650
rect 76649 541592 76654 541648
rect 76710 541592 148782 541648
rect 148838 541592 148843 541648
rect 76649 541590 148843 541592
rect 76649 541587 76715 541590
rect 148777 541587 148843 541590
rect 166441 541650 166507 541653
rect 428733 541650 428799 541653
rect 166441 541648 428799 541650
rect 166441 541592 166446 541648
rect 166502 541592 428738 541648
rect 428794 541592 428799 541648
rect 166441 541590 428799 541592
rect 166441 541587 166507 541590
rect 428733 541587 428799 541590
rect 58617 541514 58683 541517
rect 253565 541514 253631 541517
rect 58617 541512 253631 541514
rect 58617 541456 58622 541512
rect 58678 541456 253570 541512
rect 253626 541456 253631 541512
rect 58617 541454 253631 541456
rect 58617 541451 58683 541454
rect 253565 541451 253631 541454
rect 287789 541514 287855 541517
rect 341149 541514 341215 541517
rect 287789 541512 341215 541514
rect 287789 541456 287794 541512
rect 287850 541456 341154 541512
rect 341210 541456 341215 541512
rect 287789 541454 341215 541456
rect 287789 541451 287855 541454
rect 341149 541451 341215 541454
rect 49233 541378 49299 541381
rect 111793 541378 111859 541381
rect 49233 541376 111859 541378
rect 49233 541320 49238 541376
rect 49294 541320 111798 541376
rect 111854 541320 111859 541376
rect 49233 541318 111859 541320
rect 49233 541315 49299 541318
rect 111793 541315 111859 541318
rect 213913 541378 213979 541381
rect 233141 541378 233207 541381
rect 213913 541376 233207 541378
rect 213913 541320 213918 541376
rect 213974 541320 233146 541376
rect 233202 541320 233207 541376
rect 213913 541318 233207 541320
rect 213913 541315 213979 541318
rect 233141 541315 233207 541318
rect 41137 541242 41203 541245
rect 172513 541242 172579 541245
rect 41137 541240 172579 541242
rect 41137 541184 41142 541240
rect 41198 541184 172518 541240
rect 172574 541184 172579 541240
rect 41137 541182 172579 541184
rect 41137 541179 41203 541182
rect 172513 541179 172579 541182
rect 31477 541106 31543 541109
rect 224217 541106 224283 541109
rect 31477 541104 224283 541106
rect 31477 541048 31482 541104
rect 31538 541048 224222 541104
rect 224278 541048 224283 541104
rect 31477 541046 224283 541048
rect 31477 541043 31543 541046
rect 224217 541043 224283 541046
rect 91829 540970 91895 540973
rect 172145 540970 172211 540973
rect 91829 540968 172211 540970
rect -960 540684 480 540924
rect 91829 540912 91834 540968
rect 91890 540912 172150 540968
rect 172206 540912 172211 540968
rect 91829 540910 172211 540912
rect 91829 540907 91895 540910
rect 172145 540907 172211 540910
rect 172329 540970 172395 540973
rect 409965 540970 410031 540973
rect 172329 540968 410031 540970
rect 172329 540912 172334 540968
rect 172390 540912 409970 540968
rect 410026 540912 410031 540968
rect 172329 540910 410031 540912
rect 172329 540907 172395 540910
rect 409965 540907 410031 540910
rect 56409 540834 56475 540837
rect 300485 540834 300551 540837
rect 56409 540832 300551 540834
rect 56409 540776 56414 540832
rect 56470 540776 300490 540832
rect 300546 540776 300551 540832
rect 56409 540774 300551 540776
rect 56409 540771 56475 540774
rect 300485 540771 300551 540774
rect 122097 540698 122163 540701
rect 225413 540698 225479 540701
rect 122097 540696 225479 540698
rect 122097 540640 122102 540696
rect 122158 540640 225418 540696
rect 225474 540640 225479 540696
rect 122097 540638 225479 540640
rect 122097 540635 122163 540638
rect 225413 540635 225479 540638
rect 239213 540698 239279 540701
rect 484669 540698 484735 540701
rect 239213 540696 484735 540698
rect 239213 540640 239218 540696
rect 239274 540640 484674 540696
rect 484730 540640 484735 540696
rect 239213 540638 484735 540640
rect 239213 540635 239279 540638
rect 484669 540635 484735 540638
rect 32806 540500 32812 540564
rect 32876 540562 32882 540564
rect 281022 540562 281028 540564
rect 32876 540502 281028 540562
rect 32876 540500 32882 540502
rect 281022 540500 281028 540502
rect 281092 540500 281098 540564
rect 292297 540562 292363 540565
rect 506933 540562 506999 540565
rect 292297 540560 506999 540562
rect 292297 540504 292302 540560
rect 292358 540504 506938 540560
rect 506994 540504 506999 540560
rect 292297 540502 506999 540504
rect 292297 540499 292363 540502
rect 506933 540499 506999 540502
rect 53373 540426 53439 540429
rect 304533 540426 304599 540429
rect 53373 540424 304599 540426
rect 53373 540368 53378 540424
rect 53434 540368 304538 540424
rect 304594 540368 304599 540424
rect 53373 540366 304599 540368
rect 53373 540363 53439 540366
rect 304533 540363 304599 540366
rect 74625 540290 74691 540293
rect 145649 540290 145715 540293
rect 74625 540288 145715 540290
rect 74625 540232 74630 540288
rect 74686 540232 145654 540288
rect 145710 540232 145715 540288
rect 74625 540230 145715 540232
rect 74625 540227 74691 540230
rect 145649 540227 145715 540230
rect 167729 540290 167795 540293
rect 442809 540290 442875 540293
rect 167729 540288 442875 540290
rect 167729 540232 167734 540288
rect 167790 540232 442814 540288
rect 442870 540232 442875 540288
rect 167729 540230 442875 540232
rect 167729 540227 167795 540230
rect 442809 540227 442875 540230
rect 272006 540092 272012 540156
rect 272076 540154 272082 540156
rect 494462 540154 494468 540156
rect 272076 540094 494468 540154
rect 272076 540092 272082 540094
rect 494462 540092 494468 540094
rect 494532 540092 494538 540156
rect 38377 540018 38443 540021
rect 75821 540018 75887 540021
rect 38377 540016 75887 540018
rect 38377 539960 38382 540016
rect 38438 539960 75826 540016
rect 75882 539960 75887 540016
rect 38377 539958 75887 539960
rect 38377 539955 38443 539958
rect 75821 539955 75887 539958
rect 35525 539882 35591 539885
rect 91093 539882 91159 539885
rect 35525 539880 91159 539882
rect 35525 539824 35530 539880
rect 35586 539824 91098 539880
rect 91154 539824 91159 539880
rect 35525 539822 91159 539824
rect 35525 539819 35591 539822
rect 91093 539819 91159 539822
rect 47669 539746 47735 539749
rect 121453 539746 121519 539749
rect 47669 539744 121519 539746
rect 47669 539688 47674 539744
rect 47730 539688 121458 539744
rect 121514 539688 121519 539744
rect 47669 539686 121519 539688
rect 47669 539683 47735 539686
rect 121453 539683 121519 539686
rect 54569 539610 54635 539613
rect 272517 539610 272583 539613
rect 54569 539608 272583 539610
rect 54569 539552 54574 539608
rect 54630 539552 272522 539608
rect 272578 539552 272583 539608
rect 54569 539550 272583 539552
rect 54569 539547 54635 539550
rect 272517 539547 272583 539550
rect 57881 539474 57947 539477
rect 264329 539474 264395 539477
rect 57881 539472 264395 539474
rect 57881 539416 57886 539472
rect 57942 539416 264334 539472
rect 264390 539416 264395 539472
rect 57881 539414 264395 539416
rect 57881 539411 57947 539414
rect 264329 539411 264395 539414
rect 86769 539338 86835 539341
rect 164417 539338 164483 539341
rect 86769 539336 164483 539338
rect 86769 539280 86774 539336
rect 86830 539280 164422 539336
rect 164478 539280 164483 539336
rect 86769 539278 164483 539280
rect 86769 539275 86835 539278
rect 164417 539275 164483 539278
rect 173617 539338 173683 539341
rect 389633 539338 389699 539341
rect 173617 539336 389699 539338
rect 173617 539280 173622 539336
rect 173678 539280 389638 539336
rect 389694 539280 389699 539336
rect 173617 539278 389699 539280
rect 173617 539275 173683 539278
rect 389633 539275 389699 539278
rect 56133 539202 56199 539205
rect 272333 539202 272399 539205
rect 56133 539200 272399 539202
rect 56133 539144 56138 539200
rect 56194 539144 272338 539200
rect 272394 539144 272399 539200
rect 56133 539142 272399 539144
rect 56133 539139 56199 539142
rect 272333 539139 272399 539142
rect 276657 539202 276723 539205
rect 338021 539202 338087 539205
rect 276657 539200 338087 539202
rect 276657 539144 276662 539200
rect 276718 539144 338026 539200
rect 338082 539144 338087 539200
rect 276657 539142 338087 539144
rect 276657 539139 276723 539142
rect 338021 539139 338087 539142
rect 131297 539066 131363 539069
rect 240777 539066 240843 539069
rect 131297 539064 240843 539066
rect 131297 539008 131302 539064
rect 131358 539008 240782 539064
rect 240838 539008 240843 539064
rect 131297 539006 240843 539008
rect 131297 539003 131363 539006
rect 240777 539003 240843 539006
rect 257889 539066 257955 539069
rect 479885 539066 479951 539069
rect 257889 539064 479951 539066
rect 257889 539008 257894 539064
rect 257950 539008 479890 539064
rect 479946 539008 479951 539064
rect 257889 539006 479951 539008
rect 257889 539003 257955 539006
rect 479885 539003 479951 539006
rect 119337 538930 119403 538933
rect 222285 538930 222351 538933
rect 119337 538928 222351 538930
rect 119337 538872 119342 538928
rect 119398 538872 222290 538928
rect 222346 538872 222351 538928
rect 119337 538870 222351 538872
rect 119337 538867 119403 538870
rect 222285 538867 222351 538870
rect 240225 538930 240291 538933
rect 483473 538930 483539 538933
rect 240225 538928 483539 538930
rect 240225 538872 240230 538928
rect 240286 538872 483478 538928
rect 483534 538872 483539 538928
rect 240225 538870 483539 538872
rect 240225 538867 240291 538870
rect 483473 538867 483539 538870
rect 61561 538794 61627 538797
rect 336917 538794 336983 538797
rect 61561 538792 336983 538794
rect 61561 538736 61566 538792
rect 61622 538736 336922 538792
rect 336978 538736 336983 538792
rect 61561 538734 336983 538736
rect 61561 538731 61627 538734
rect 336917 538731 336983 538734
rect 71589 538658 71655 538661
rect 140957 538658 141023 538661
rect 71589 538656 141023 538658
rect 71589 538600 71594 538656
rect 71650 538600 140962 538656
rect 141018 538600 141023 538656
rect 71589 538598 141023 538600
rect 71589 538595 71655 538598
rect 140957 538595 141023 538598
rect 152457 538658 152523 538661
rect 311433 538658 311499 538661
rect 152457 538656 311499 538658
rect 152457 538600 152462 538656
rect 152518 538600 311438 538656
rect 311494 538600 311499 538656
rect 152457 538598 311499 538600
rect 152457 538595 152523 538598
rect 311433 538595 311499 538598
rect 50337 538522 50403 538525
rect 86861 538522 86927 538525
rect 50337 538520 86927 538522
rect 50337 538464 50342 538520
rect 50398 538464 86866 538520
rect 86922 538464 86927 538520
rect 50337 538462 86927 538464
rect 50337 538459 50403 538462
rect 86861 538459 86927 538462
rect 227069 538522 227135 538525
rect 256693 538522 256759 538525
rect 227069 538520 256759 538522
rect 227069 538464 227074 538520
rect 227130 538464 256698 538520
rect 256754 538464 256759 538520
rect 227069 538462 256759 538464
rect 227069 538459 227135 538462
rect 256693 538459 256759 538462
rect 55949 538386 56015 538389
rect 118693 538386 118759 538389
rect 55949 538384 118759 538386
rect 55949 538328 55954 538384
rect 56010 538328 118698 538384
rect 118754 538328 118759 538384
rect 55949 538326 118759 538328
rect 55949 538323 56015 538326
rect 118693 538323 118759 538326
rect 56409 538250 56475 538253
rect 131113 538250 131179 538253
rect 56409 538248 131179 538250
rect 56409 538192 56414 538248
rect 56470 538192 131118 538248
rect 131174 538192 131179 538248
rect 56409 538190 131179 538192
rect 56409 538187 56475 538190
rect 131113 538187 131179 538190
rect 59721 538114 59787 538117
rect 275461 538114 275527 538117
rect 59721 538112 275527 538114
rect 59721 538056 59726 538112
rect 59782 538056 275466 538112
rect 275522 538056 275527 538112
rect 59721 538054 275527 538056
rect 59721 538051 59787 538054
rect 275461 538051 275527 538054
rect 292389 538114 292455 538117
rect 482134 538114 482140 538116
rect 292389 538112 482140 538114
rect 292389 538056 292394 538112
rect 292450 538056 482140 538112
rect 292389 538054 482140 538056
rect 292389 538051 292455 538054
rect 482134 538052 482140 538054
rect 482204 538052 482210 538116
rect 251357 537978 251423 537981
rect 484761 537978 484827 537981
rect 251357 537976 484827 537978
rect 251357 537920 251362 537976
rect 251418 537920 484766 537976
rect 484822 537920 484827 537976
rect 251357 537918 484827 537920
rect 251357 537915 251423 537918
rect 484761 537915 484827 537918
rect 123201 537842 123267 537845
rect 230105 537842 230171 537845
rect 123201 537840 230171 537842
rect 123201 537784 123206 537840
rect 123262 537784 230110 537840
rect 230166 537784 230171 537840
rect 123201 537782 230171 537784
rect 123201 537779 123267 537782
rect 230105 537779 230171 537782
rect 236177 537842 236243 537845
rect 483381 537842 483447 537845
rect 236177 537840 483447 537842
rect 236177 537784 236182 537840
rect 236238 537784 483386 537840
rect 483442 537784 483447 537840
rect 236177 537782 483447 537784
rect 236177 537779 236243 537782
rect 483381 537779 483447 537782
rect 580533 537842 580599 537845
rect 583520 537842 584960 537932
rect 580533 537840 584960 537842
rect 580533 537784 580538 537840
rect 580594 537784 584960 537840
rect 580533 537782 584960 537784
rect 580533 537779 580599 537782
rect 43437 537706 43503 537709
rect 60825 537706 60891 537709
rect 43437 537704 60891 537706
rect 43437 537648 43442 537704
rect 43498 537648 60830 537704
rect 60886 537648 60891 537704
rect 43437 537646 60891 537648
rect 43437 537643 43503 537646
rect 60825 537643 60891 537646
rect 172053 537706 172119 537709
rect 419349 537706 419415 537709
rect 172053 537704 419415 537706
rect 172053 537648 172058 537704
rect 172114 537648 419354 537704
rect 419410 537648 419415 537704
rect 583520 537692 584960 537782
rect 172053 537646 419415 537648
rect 172053 537643 172119 537646
rect 419349 537643 419415 537646
rect 61469 537570 61535 537573
rect 125317 537570 125383 537573
rect 61469 537568 125383 537570
rect 61469 537512 61474 537568
rect 61530 537512 125322 537568
rect 125378 537512 125383 537568
rect 61469 537510 125383 537512
rect 61469 537507 61535 537510
rect 125317 537507 125383 537510
rect 164969 537570 165035 537573
rect 438117 537570 438183 537573
rect 164969 537568 438183 537570
rect 164969 537512 164974 537568
rect 165030 537512 438122 537568
rect 438178 537512 438183 537568
rect 164969 537510 438183 537512
rect 164969 537507 165035 537510
rect 438117 537507 438183 537510
rect 60181 537434 60247 537437
rect 82813 537434 82879 537437
rect 60181 537432 82879 537434
rect 60181 537376 60186 537432
rect 60242 537376 82818 537432
rect 82874 537376 82879 537432
rect 60181 537374 82879 537376
rect 60181 537371 60247 537374
rect 82813 537371 82879 537374
rect 83733 537434 83799 537437
rect 159725 537434 159791 537437
rect 83733 537432 159791 537434
rect 83733 537376 83738 537432
rect 83794 537376 159730 537432
rect 159786 537376 159791 537432
rect 83733 537374 159791 537376
rect 83733 537371 83799 537374
rect 159725 537371 159791 537374
rect 165470 537372 165476 537436
rect 165540 537434 165546 537436
rect 171041 537434 171107 537437
rect 445937 537434 446003 537437
rect 165540 537432 171107 537434
rect 165540 537376 171046 537432
rect 171102 537376 171107 537432
rect 165540 537374 171107 537376
rect 165540 537372 165546 537374
rect 171041 537371 171107 537374
rect 176610 537432 446003 537434
rect 176610 537376 445942 537432
rect 445998 537376 446003 537432
rect 176610 537374 446003 537376
rect 49049 537298 49115 537301
rect 124121 537298 124187 537301
rect 49049 537296 124187 537298
rect 49049 537240 49054 537296
rect 49110 537240 124126 537296
rect 124182 537240 124187 537296
rect 49049 537238 124187 537240
rect 49049 537235 49115 537238
rect 124121 537235 124187 537238
rect 170489 537298 170555 537301
rect 176610 537298 176670 537374
rect 445937 537371 446003 537374
rect 170489 537296 176670 537298
rect 170489 537240 170494 537296
rect 170550 537240 176670 537296
rect 170489 537238 176670 537240
rect 280797 537298 280863 537301
rect 359917 537298 359983 537301
rect 280797 537296 359983 537298
rect 280797 537240 280802 537296
rect 280858 537240 359922 537296
rect 359978 537240 359983 537296
rect 280797 537238 359983 537240
rect 170489 537235 170555 537238
rect 280797 537235 280863 537238
rect 359917 537235 359983 537238
rect 53005 537162 53071 537165
rect 171777 537162 171843 537165
rect 53005 537160 171843 537162
rect 53005 537104 53010 537160
rect 53066 537104 171782 537160
rect 171838 537104 171843 537160
rect 53005 537102 171843 537104
rect 53005 537099 53071 537102
rect 171777 537099 171843 537102
rect 45185 537026 45251 537029
rect 252461 537026 252527 537029
rect 45185 537024 252527 537026
rect 45185 536968 45190 537024
rect 45246 536968 252466 537024
rect 252522 536968 252527 537024
rect 45185 536966 252527 536968
rect 45185 536963 45251 536966
rect 252461 536963 252527 536966
rect 32438 536828 32444 536892
rect 32508 536890 32514 536892
rect 291837 536890 291903 536893
rect 32508 536888 291903 536890
rect 32508 536832 291842 536888
rect 291898 536832 291903 536888
rect 32508 536830 291903 536832
rect 32508 536828 32514 536830
rect 291837 536827 291903 536830
rect 171777 536754 171843 536757
rect 173985 536754 174051 536757
rect 171777 536752 174051 536754
rect 171777 536696 171782 536752
rect 171838 536696 173990 536752
rect 174046 536696 174051 536752
rect 171777 536694 174051 536696
rect 171777 536691 171843 536694
rect 173985 536691 174051 536694
rect 179045 536754 179111 536757
rect 397361 536754 397427 536757
rect 179045 536752 397427 536754
rect 179045 536696 179050 536752
rect 179106 536696 397366 536752
rect 397422 536696 397427 536752
rect 179045 536694 397427 536696
rect 179045 536691 179111 536694
rect 397361 536691 397427 536694
rect 66529 536618 66595 536621
rect 133137 536618 133203 536621
rect 66529 536616 133203 536618
rect 66529 536560 66534 536616
rect 66590 536560 133142 536616
rect 133198 536560 133203 536616
rect 66529 536558 133203 536560
rect 66529 536555 66595 536558
rect 133137 536555 133203 536558
rect 174997 536618 175063 536621
rect 399017 536618 399083 536621
rect 174997 536616 399083 536618
rect 174997 536560 175002 536616
rect 175058 536560 399022 536616
rect 399078 536560 399083 536616
rect 174997 536558 399083 536560
rect 174997 536555 175063 536558
rect 399017 536555 399083 536558
rect 59077 536482 59143 536485
rect 291101 536482 291167 536485
rect 59077 536480 291167 536482
rect 59077 536424 59082 536480
rect 59138 536424 291106 536480
rect 291162 536424 291167 536480
rect 59077 536422 291167 536424
rect 59077 536419 59143 536422
rect 291101 536419 291167 536422
rect 293769 536482 293835 536485
rect 482001 536482 482067 536485
rect 293769 536480 482067 536482
rect 293769 536424 293774 536480
rect 293830 536424 482006 536480
rect 482062 536424 482067 536480
rect 293769 536422 482067 536424
rect 293769 536419 293835 536422
rect 482001 536419 482067 536422
rect 129273 536346 129339 536349
rect 239489 536346 239555 536349
rect 129273 536344 239555 536346
rect 129273 536288 129278 536344
rect 129334 536288 239494 536344
rect 239550 536288 239555 536344
rect 129273 536286 239555 536288
rect 129273 536283 129339 536286
rect 239489 536283 239555 536286
rect 253381 536346 253447 536349
rect 490465 536346 490531 536349
rect 253381 536344 490531 536346
rect 253381 536288 253386 536344
rect 253442 536288 490470 536344
rect 490526 536288 490531 536344
rect 253381 536286 490531 536288
rect 253381 536283 253447 536286
rect 490465 536283 490531 536286
rect 97809 536210 97875 536213
rect 191005 536210 191071 536213
rect 97809 536208 191071 536210
rect 97809 536152 97814 536208
rect 97870 536152 191010 536208
rect 191066 536152 191071 536208
rect 97809 536150 191071 536152
rect 97809 536147 97875 536150
rect 191005 536147 191071 536150
rect 192661 536210 192727 536213
rect 205633 536210 205699 536213
rect 192661 536208 205699 536210
rect 192661 536152 192666 536208
rect 192722 536152 205638 536208
rect 205694 536152 205699 536208
rect 192661 536150 205699 536152
rect 192661 536147 192727 536150
rect 205633 536147 205699 536150
rect 206829 536210 206895 536213
rect 218053 536210 218119 536213
rect 206829 536208 218119 536210
rect 206829 536152 206834 536208
rect 206890 536152 218058 536208
rect 218114 536152 218119 536208
rect 206829 536150 218119 536152
rect 206829 536147 206895 536150
rect 218053 536147 218119 536150
rect 218973 536210 219039 536213
rect 499757 536210 499823 536213
rect 218973 536208 499823 536210
rect 218973 536152 218978 536208
rect 219034 536152 499762 536208
rect 499818 536152 499823 536208
rect 218973 536150 499823 536152
rect 218973 536147 219039 536150
rect 499757 536147 499823 536150
rect 30046 536012 30052 536076
rect 30116 536074 30122 536076
rect 382222 536074 382228 536076
rect 30116 536014 382228 536074
rect 30116 536012 30122 536014
rect 382222 536012 382228 536014
rect 382292 536012 382298 536076
rect 49325 535938 49391 535941
rect 97901 535938 97967 535941
rect 49325 535936 97967 535938
rect 49325 535880 49330 535936
rect 49386 535880 97906 535936
rect 97962 535880 97967 535936
rect 49325 535878 97967 535880
rect 49325 535875 49391 535878
rect 97901 535875 97967 535878
rect 291837 535938 291903 535941
rect 331765 535938 331831 535941
rect 291837 535936 331831 535938
rect 291837 535880 291842 535936
rect 291898 535880 331770 535936
rect 331826 535880 331831 535936
rect 291837 535878 331831 535880
rect 291837 535875 291903 535878
rect 331765 535875 331831 535878
rect 50429 535802 50495 535805
rect 128353 535802 128419 535805
rect 50429 535800 128419 535802
rect 50429 535744 50434 535800
rect 50490 535744 128358 535800
rect 128414 535744 128419 535800
rect 50429 535742 128419 535744
rect 50429 535739 50495 535742
rect 128353 535739 128419 535742
rect 54477 535666 54543 535669
rect 178033 535666 178099 535669
rect 54477 535664 178099 535666
rect 54477 535608 54482 535664
rect 54538 535608 178038 535664
rect 178094 535608 178099 535664
rect 54477 535606 178099 535608
rect 54477 535603 54543 535606
rect 178033 535603 178099 535606
rect 56317 535530 56383 535533
rect 292573 535530 292639 535533
rect 56317 535528 292639 535530
rect 56317 535472 56322 535528
rect 56378 535472 292578 535528
rect 292634 535472 292639 535528
rect 56317 535470 292639 535472
rect 56317 535467 56383 535470
rect 292573 535467 292639 535470
rect 96889 535394 96955 535397
rect 164141 535394 164207 535397
rect 96889 535392 164207 535394
rect 96889 535336 96894 535392
rect 96950 535336 164146 535392
rect 164202 535336 164207 535392
rect 96889 535334 164207 535336
rect 96889 535331 96955 535334
rect 164141 535331 164207 535334
rect 193673 535394 193739 535397
rect 212441 535394 212507 535397
rect 193673 535392 212507 535394
rect 193673 535336 193678 535392
rect 193734 535336 212446 535392
rect 212502 535336 212507 535392
rect 193673 535334 212507 535336
rect 193673 535331 193739 535334
rect 212441 535331 212507 535334
rect 243261 535394 243327 535397
rect 483565 535394 483631 535397
rect 243261 535392 483631 535394
rect 243261 535336 243266 535392
rect 243322 535336 483570 535392
rect 483626 535336 483631 535392
rect 243261 535334 483631 535336
rect 243261 535331 243327 535334
rect 483565 535331 483631 535334
rect 32622 535196 32628 535260
rect 32692 535258 32698 535260
rect 276974 535258 276980 535260
rect 32692 535198 276980 535258
rect 32692 535196 32698 535198
rect 276974 535196 276980 535198
rect 277044 535196 277050 535260
rect 279509 535258 279575 535261
rect 336457 535258 336523 535261
rect 279509 535256 336523 535258
rect 279509 535200 279514 535256
rect 279570 535200 336462 535256
rect 336518 535200 336523 535256
rect 279509 535198 336523 535200
rect 279509 535195 279575 535198
rect 336457 535195 336523 535198
rect 35750 535060 35756 535124
rect 35820 535122 35826 535124
rect 285254 535122 285260 535124
rect 35820 535062 285260 535122
rect 35820 535060 35826 535062
rect 285254 535060 285260 535062
rect 285324 535060 285330 535124
rect 296437 535122 296503 535125
rect 496077 535122 496143 535125
rect 296437 535120 496143 535122
rect 296437 535064 296442 535120
rect 296498 535064 496082 535120
rect 496138 535064 496143 535120
rect 296437 535062 496143 535064
rect 296437 535059 296503 535062
rect 496077 535059 496143 535062
rect 55489 534986 55555 534989
rect 306741 534986 306807 534989
rect 55489 534984 306807 534986
rect 55489 534928 55494 534984
rect 55550 534928 306746 534984
rect 306802 534928 306807 534984
rect 55489 534926 306807 534928
rect 55489 534923 55555 534926
rect 306741 534923 306807 534926
rect 42374 534788 42380 534852
rect 42444 534850 42450 534852
rect 379646 534850 379652 534852
rect 42444 534790 379652 534850
rect 42444 534788 42450 534790
rect 379646 534788 379652 534790
rect 379716 534788 379722 534852
rect 30966 534652 30972 534716
rect 31036 534714 31042 534716
rect 383694 534714 383700 534716
rect 31036 534654 383700 534714
rect 31036 534652 31042 534654
rect 383694 534652 383700 534654
rect 383764 534652 383770 534716
rect 155493 534578 155559 534581
rect 333329 534578 333395 534581
rect 155493 534576 333395 534578
rect 155493 534520 155498 534576
rect 155554 534520 333334 534576
rect 333390 534520 333395 534576
rect 155493 534518 333395 534520
rect 155493 534515 155559 534518
rect 333329 534515 333395 534518
rect 163497 534442 163563 534445
rect 184749 534442 184815 534445
rect 163497 534440 184815 534442
rect 163497 534384 163502 534440
rect 163558 534384 184754 534440
rect 184810 534384 184815 534440
rect 163497 534382 184815 534384
rect 163497 534379 163563 534382
rect 184749 534379 184815 534382
rect 185577 534442 185643 534445
rect 194501 534442 194567 534445
rect 185577 534440 194567 534442
rect 185577 534384 185582 534440
rect 185638 534384 194506 534440
rect 194562 534384 194567 534440
rect 185577 534382 194567 534384
rect 185577 534379 185643 534382
rect 194501 534379 194567 534382
rect 211889 534442 211955 534445
rect 243537 534442 243603 534445
rect 211889 534440 243603 534442
rect 211889 534384 211894 534440
rect 211950 534384 243542 534440
rect 243598 534384 243603 534440
rect 211889 534382 243603 534384
rect 211889 534379 211955 534382
rect 243537 534379 243603 534382
rect 60273 534306 60339 534309
rect 97901 534306 97967 534309
rect 60273 534304 97967 534306
rect 60273 534248 60278 534304
rect 60334 534248 97906 534304
rect 97962 534248 97967 534304
rect 60273 534246 97967 534248
rect 60273 534243 60339 534246
rect 97901 534243 97967 534246
rect 31702 534108 31708 534172
rect 31772 534170 31778 534172
rect 33041 534170 33107 534173
rect 31772 534168 33107 534170
rect 31772 534112 33046 534168
rect 33102 534112 33107 534168
rect 31772 534110 33107 534112
rect 31772 534108 31778 534110
rect 33041 534107 33107 534110
rect 56041 534170 56107 534173
rect 155861 534170 155927 534173
rect 56041 534168 155927 534170
rect 56041 534112 56046 534168
rect 56102 534112 155866 534168
rect 155922 534112 155927 534168
rect 56041 534110 155927 534112
rect 56041 534107 56107 534110
rect 155861 534107 155927 534110
rect 379605 534170 379671 534173
rect 379830 534170 379836 534172
rect 379605 534168 379836 534170
rect 379605 534112 379610 534168
rect 379666 534112 379836 534168
rect 379605 534110 379836 534112
rect 379605 534107 379671 534110
rect 379830 534108 379836 534110
rect 379900 534108 379906 534172
rect 176285 534034 176351 534037
rect 395889 534034 395955 534037
rect 176285 534032 395955 534034
rect 176285 533976 176290 534032
rect 176346 533976 395894 534032
rect 395950 533976 395955 534032
rect 176285 533974 395955 533976
rect 176285 533971 176351 533974
rect 395889 533971 395955 533974
rect 59077 533898 59143 533901
rect 295793 533898 295859 533901
rect 59077 533896 295859 533898
rect 59077 533840 59082 533896
rect 59138 533840 295798 533896
rect 295854 533840 295859 533896
rect 59077 533838 295859 533840
rect 59077 533835 59143 533838
rect 295793 533835 295859 533838
rect 296529 533898 296595 533901
rect 481909 533898 481975 533901
rect 296529 533896 481975 533898
rect 296529 533840 296534 533896
rect 296590 533840 481914 533896
rect 481970 533840 481975 533896
rect 296529 533838 481975 533840
rect 296529 533835 296595 533838
rect 481909 533835 481975 533838
rect 48957 533762 49023 533765
rect 60733 533762 60799 533765
rect 48957 533760 60799 533762
rect 48957 533704 48962 533760
rect 49018 533704 60738 533760
rect 60794 533704 60799 533760
rect 48957 533702 60799 533704
rect 48957 533699 49023 533702
rect 60733 533699 60799 533702
rect 162209 533762 162275 533765
rect 181621 533762 181687 533765
rect 162209 533760 181687 533762
rect 162209 533704 162214 533760
rect 162270 533704 181626 533760
rect 181682 533704 181687 533760
rect 162209 533702 181687 533704
rect 162209 533699 162275 533702
rect 181621 533699 181687 533702
rect 184565 533762 184631 533765
rect 191741 533762 191807 533765
rect 184565 533760 191807 533762
rect 184565 533704 184570 533760
rect 184626 533704 191746 533760
rect 191802 533704 191807 533760
rect 184565 533702 191807 533704
rect 184565 533699 184631 533702
rect 191741 533699 191807 533702
rect 191925 533762 191991 533765
rect 244365 533762 244431 533765
rect 191925 533760 244431 533762
rect 191925 533704 191930 533760
rect 191986 533704 244370 533760
rect 244426 533704 244431 533760
rect 191925 533702 244431 533704
rect 191925 533699 191991 533702
rect 244365 533699 244431 533702
rect 245285 533762 245351 533765
rect 486417 533762 486483 533765
rect 245285 533760 486483 533762
rect 245285 533704 245290 533760
rect 245346 533704 486422 533760
rect 486478 533704 486483 533760
rect 245285 533702 486483 533704
rect 245285 533699 245351 533702
rect 486417 533699 486483 533702
rect 39389 533626 39455 533629
rect 59169 533626 59235 533629
rect 39389 533624 59235 533626
rect 39389 533568 39394 533624
rect 39450 533568 59174 533624
rect 59230 533568 59235 533624
rect 39389 533566 59235 533568
rect 39389 533563 39455 533566
rect 59169 533563 59235 533566
rect 70669 533626 70735 533629
rect 139301 533626 139367 533629
rect 70669 533624 139367 533626
rect 70669 533568 70674 533624
rect 70730 533568 139306 533624
rect 139362 533568 139367 533624
rect 70669 533566 139367 533568
rect 70669 533563 70735 533566
rect 139301 533563 139367 533566
rect 167821 533626 167887 533629
rect 427169 533626 427235 533629
rect 167821 533624 427235 533626
rect 167821 533568 167826 533624
rect 167882 533568 427174 533624
rect 427230 533568 427235 533624
rect 167821 533566 427235 533568
rect 167821 533563 167887 533566
rect 427169 533563 427235 533566
rect 42517 533490 42583 533493
rect 324773 533490 324839 533493
rect 42517 533488 324839 533490
rect 42517 533432 42522 533488
rect 42578 533432 324778 533488
rect 324834 533432 324839 533488
rect 42517 533430 324839 533432
rect 42517 533427 42583 533430
rect 324773 533427 324839 533430
rect 29126 533292 29132 533356
rect 29196 533354 29202 533356
rect 30281 533354 30347 533357
rect 379462 533354 379468 533356
rect 29196 533352 30347 533354
rect 29196 533296 30286 533352
rect 30342 533296 30347 533352
rect 29196 533294 30347 533296
rect 29196 533292 29202 533294
rect 30281 533291 30347 533294
rect 35850 533294 379468 533354
rect 29862 533156 29868 533220
rect 29932 533218 29938 533220
rect 35850 533218 35910 533294
rect 379462 533292 379468 533294
rect 379532 533292 379538 533356
rect 29932 533158 35910 533218
rect 60733 533218 60799 533221
rect 255129 533218 255195 533221
rect 60733 533216 255195 533218
rect 60733 533160 60738 533216
rect 60794 533160 255134 533216
rect 255190 533160 255195 533216
rect 60733 533158 255195 533160
rect 29932 533156 29938 533158
rect 60733 533155 60799 533158
rect 255129 533155 255195 533158
rect 283414 533156 283420 533220
rect 283484 533218 283490 533220
rect 495382 533218 495388 533220
rect 283484 533158 495388 533218
rect 283484 533156 283490 533158
rect 495382 533156 495388 533158
rect 495452 533156 495458 533220
rect 34145 533082 34211 533085
rect 70393 533082 70459 533085
rect 34145 533080 70459 533082
rect 34145 533024 34150 533080
rect 34206 533024 70398 533080
rect 70454 533024 70459 533080
rect 34145 533022 70459 533024
rect 34145 533019 34211 533022
rect 70393 533019 70459 533022
rect 55857 532946 55923 532949
rect 166993 532946 167059 532949
rect 55857 532944 167059 532946
rect 55857 532888 55862 532944
rect 55918 532888 166998 532944
rect 167054 532888 167059 532944
rect 55857 532886 167059 532888
rect 55857 532883 55923 532886
rect 166993 532883 167059 532886
rect 54385 532810 54451 532813
rect 175825 532810 175891 532813
rect 54385 532808 175891 532810
rect 54385 532752 54390 532808
rect 54446 532752 175830 532808
rect 175886 532752 175891 532808
rect 54385 532750 175891 532752
rect 54385 532747 54451 532750
rect 175825 532747 175891 532750
rect 178953 532674 179019 532677
rect 394325 532674 394391 532677
rect 178953 532672 394391 532674
rect 178953 532616 178958 532672
rect 179014 532616 394330 532672
rect 394386 532616 394391 532672
rect 178953 532614 394391 532616
rect 178953 532611 179019 532614
rect 394325 532611 394391 532614
rect 58985 532538 59051 532541
rect 286409 532538 286475 532541
rect 58985 532536 286475 532538
rect 58985 532480 58990 532536
rect 59046 532480 286414 532536
rect 286470 532480 286475 532536
rect 58985 532478 286475 532480
rect 58985 532475 59051 532478
rect 286409 532475 286475 532478
rect 132309 532402 132375 532405
rect 218697 532402 218763 532405
rect 132309 532400 218763 532402
rect 132309 532344 132314 532400
rect 132370 532344 218702 532400
rect 218758 532344 218763 532400
rect 132309 532342 218763 532344
rect 132309 532339 132375 532342
rect 218697 532339 218763 532342
rect 266854 532340 266860 532404
rect 266924 532402 266930 532404
rect 502926 532402 502932 532404
rect 266924 532342 502932 532402
rect 266924 532340 266930 532342
rect 502926 532340 502932 532342
rect 502996 532340 503002 532404
rect 50245 532266 50311 532269
rect 96521 532266 96587 532269
rect 50245 532264 96587 532266
rect 50245 532208 50250 532264
rect 50306 532208 96526 532264
rect 96582 532208 96587 532264
rect 50245 532206 96587 532208
rect 50245 532203 50311 532206
rect 96521 532203 96587 532206
rect 117129 532266 117195 532269
rect 220721 532266 220787 532269
rect 117129 532264 220787 532266
rect 117129 532208 117134 532264
rect 117190 532208 220726 532264
rect 220782 532208 220787 532264
rect 117129 532206 220787 532208
rect 117129 532203 117195 532206
rect 220721 532203 220787 532206
rect 248321 532266 248387 532269
rect 484945 532266 485011 532269
rect 248321 532264 485011 532266
rect 248321 532208 248326 532264
rect 248382 532208 484950 532264
rect 485006 532208 485011 532264
rect 248321 532206 485011 532208
rect 248321 532203 248387 532206
rect 484945 532203 485011 532206
rect 68553 532130 68619 532133
rect 136265 532130 136331 532133
rect 68553 532128 136331 532130
rect 68553 532072 68558 532128
rect 68614 532072 136270 532128
rect 136326 532072 136331 532128
rect 68553 532070 136331 532072
rect 68553 532067 68619 532070
rect 136265 532067 136331 532070
rect 148317 532130 148383 532133
rect 180057 532130 180123 532133
rect 148317 532128 180123 532130
rect 148317 532072 148322 532128
rect 148378 532072 180062 532128
rect 180118 532072 180123 532128
rect 148317 532070 180123 532072
rect 148317 532067 148383 532070
rect 180057 532067 180123 532070
rect 212901 532130 212967 532133
rect 481081 532130 481147 532133
rect 212901 532128 481147 532130
rect 212901 532072 212906 532128
rect 212962 532072 481086 532128
rect 481142 532072 481147 532128
rect 212901 532070 481147 532072
rect 212901 532067 212967 532070
rect 481081 532067 481147 532070
rect 484301 532130 484367 532133
rect 507945 532130 508011 532133
rect 484301 532128 508011 532130
rect 484301 532072 484306 532128
rect 484362 532072 507950 532128
rect 508006 532072 508011 532128
rect 484301 532070 508011 532072
rect 484301 532067 484367 532070
rect 507945 532067 508011 532070
rect 95877 531994 95943 531997
rect 189441 531994 189507 531997
rect 95877 531992 189507 531994
rect 95877 531936 95882 531992
rect 95938 531936 189446 531992
rect 189502 531936 189507 531992
rect 95877 531934 189507 531936
rect 95877 531931 95943 531934
rect 189441 531931 189507 531934
rect 198733 531994 198799 531997
rect 498377 531994 498443 531997
rect 198733 531992 498443 531994
rect 198733 531936 198738 531992
rect 198794 531936 498382 531992
rect 498438 531936 498443 531992
rect 198733 531934 498443 531936
rect 198733 531931 198799 531934
rect 498377 531931 498443 531934
rect 59813 531858 59879 531861
rect 267641 531858 267707 531861
rect 59813 531856 267707 531858
rect 59813 531800 59818 531856
rect 59874 531800 267646 531856
rect 267702 531800 267707 531856
rect 59813 531798 267707 531800
rect 59813 531795 59879 531798
rect 267641 531795 267707 531798
rect 286174 531796 286180 531860
rect 286244 531858 286250 531860
rect 498142 531858 498148 531860
rect 286244 531798 498148 531858
rect 286244 531796 286250 531798
rect 498142 531796 498148 531798
rect 498212 531796 498218 531860
rect 40769 531722 40835 531725
rect 117221 531722 117287 531725
rect 40769 531720 117287 531722
rect 40769 531664 40774 531720
rect 40830 531664 117226 531720
rect 117282 531664 117287 531720
rect 40769 531662 117287 531664
rect 40769 531659 40835 531662
rect 117221 531659 117287 531662
rect 197721 531722 197787 531725
rect 213821 531722 213887 531725
rect 197721 531720 213887 531722
rect 197721 531664 197726 531720
rect 197782 531664 213826 531720
rect 213882 531664 213887 531720
rect 197721 531662 213887 531664
rect 197721 531659 197787 531662
rect 213821 531659 213887 531662
rect 39573 531586 39639 531589
rect 131113 531586 131179 531589
rect 39573 531584 131179 531586
rect 39573 531528 39578 531584
rect 39634 531528 131118 531584
rect 131174 531528 131179 531584
rect 39573 531526 131179 531528
rect 39573 531523 39639 531526
rect 131113 531523 131179 531526
rect 37038 531388 37044 531452
rect 37108 531450 37114 531452
rect 178033 531450 178099 531453
rect 37108 531448 178099 531450
rect 37108 531392 178038 531448
rect 178094 531392 178099 531448
rect 37108 531390 178099 531392
rect 37108 531388 37114 531390
rect 178033 531387 178099 531390
rect 211061 531450 211127 531453
rect 211061 531448 211354 531450
rect 211061 531392 211066 531448
rect 211122 531392 211354 531448
rect 211061 531390 211354 531392
rect 211061 531387 211127 531390
rect 39481 531314 39547 531317
rect 211061 531314 211127 531317
rect 39481 531312 211127 531314
rect 39481 531256 39486 531312
rect 39542 531256 211066 531312
rect 211122 531256 211127 531312
rect 39481 531254 211127 531256
rect 211294 531314 211354 531390
rect 251081 531314 251147 531317
rect 211294 531312 251147 531314
rect 211294 531256 251086 531312
rect 251142 531256 251147 531312
rect 211294 531254 251147 531256
rect 39481 531251 39547 531254
rect 211061 531251 211127 531254
rect 251081 531251 251147 531254
rect 282126 531252 282132 531316
rect 282196 531314 282202 531316
rect 295333 531314 295399 531317
rect 282196 531312 295399 531314
rect 282196 531256 295338 531312
rect 295394 531256 295399 531312
rect 282196 531254 295399 531256
rect 282196 531252 282202 531254
rect 295333 531251 295399 531254
rect 67633 531178 67699 531181
rect 134701 531178 134767 531181
rect 67633 531176 134767 531178
rect 67633 531120 67638 531176
rect 67694 531120 134706 531176
rect 134762 531120 134767 531176
rect 67633 531118 134767 531120
rect 67633 531115 67699 531118
rect 134701 531115 134767 531118
rect 173157 531178 173223 531181
rect 449065 531178 449131 531181
rect 173157 531176 449131 531178
rect 173157 531120 173162 531176
rect 173218 531120 449070 531176
rect 449126 531120 449131 531176
rect 173157 531118 449131 531120
rect 173157 531115 173223 531118
rect 449065 531115 449131 531118
rect 40953 531042 41019 531045
rect 319713 531042 319779 531045
rect 40953 531040 319779 531042
rect 40953 530984 40958 531040
rect 41014 530984 319718 531040
rect 319774 530984 319779 531040
rect 40953 530982 319779 530984
rect 40953 530979 41019 530982
rect 319713 530979 319779 530982
rect 112069 530906 112135 530909
rect 212901 530906 212967 530909
rect 112069 530904 212967 530906
rect 112069 530848 112074 530904
rect 112130 530848 212906 530904
rect 212962 530848 212967 530904
rect 112069 530846 212967 530848
rect 112069 530843 112135 530846
rect 212901 530843 212967 530846
rect 220997 530906 221063 530909
rect 499941 530906 500007 530909
rect 220997 530904 500007 530906
rect 220997 530848 221002 530904
rect 221058 530848 499946 530904
rect 500002 530848 500007 530904
rect 220997 530846 500007 530848
rect 220997 530843 221063 530846
rect 499941 530843 500007 530846
rect 59537 530770 59603 530773
rect 376753 530770 376819 530773
rect 59537 530768 376819 530770
rect 59537 530712 59542 530768
rect 59598 530712 376758 530768
rect 376814 530712 376819 530768
rect 59537 530710 376819 530712
rect 59537 530707 59603 530710
rect 376753 530707 376819 530710
rect 34053 530634 34119 530637
rect 383837 530634 383903 530637
rect 34053 530632 383903 530634
rect 34053 530576 34058 530632
rect 34114 530576 383842 530632
rect 383898 530576 383903 530632
rect 34053 530574 383903 530576
rect 34053 530571 34119 530574
rect 383837 530571 383903 530574
rect 58893 530498 58959 530501
rect 280061 530498 280127 530501
rect 58893 530496 280127 530498
rect 58893 530440 58898 530496
rect 58954 530440 280066 530496
rect 280122 530440 280127 530496
rect 58893 530438 280127 530440
rect 58893 530435 58959 530438
rect 280061 530435 280127 530438
rect 288566 530436 288572 530500
rect 288636 530498 288642 530500
rect 289721 530498 289787 530501
rect 288636 530496 289787 530498
rect 288636 530440 289726 530496
rect 289782 530440 289787 530496
rect 288636 530438 289787 530440
rect 288636 530436 288642 530438
rect 289721 530435 289787 530438
rect 296621 530498 296687 530501
rect 482093 530498 482159 530501
rect 296621 530496 482159 530498
rect 296621 530440 296626 530496
rect 296682 530440 482098 530496
rect 482154 530440 482159 530496
rect 296621 530438 482159 530440
rect 296621 530435 296687 530438
rect 482093 530435 482159 530438
rect 38285 530362 38351 530365
rect 59169 530362 59235 530365
rect 38285 530360 59235 530362
rect 38285 530304 38290 530360
rect 38346 530304 59174 530360
rect 59230 530304 59235 530360
rect 38285 530302 59235 530304
rect 38285 530299 38351 530302
rect 59169 530299 59235 530302
rect 250345 530362 250411 530365
rect 483657 530362 483723 530365
rect 250345 530360 483723 530362
rect 250345 530304 250350 530360
rect 250406 530304 483662 530360
rect 483718 530304 483723 530360
rect 250345 530302 483723 530304
rect 250345 530299 250411 530302
rect 483657 530299 483723 530302
rect 36721 530226 36787 530229
rect 67541 530226 67607 530229
rect 36721 530224 67607 530226
rect 36721 530168 36726 530224
rect 36782 530168 67546 530224
rect 67602 530168 67607 530224
rect 36721 530166 67607 530168
rect 36721 530163 36787 530166
rect 67541 530163 67607 530166
rect 46381 530090 46447 530093
rect 111793 530090 111859 530093
rect 46381 530088 111859 530090
rect 46381 530032 46386 530088
rect 46442 530032 111798 530088
rect 111854 530032 111859 530088
rect 46381 530030 111859 530032
rect 46381 530027 46447 530030
rect 111793 530027 111859 530030
rect 52913 529954 52979 529957
rect 59905 529954 59971 529957
rect 52913 529952 59971 529954
rect 52913 529896 52918 529952
rect 52974 529896 59910 529952
rect 59966 529896 59971 529952
rect 52913 529894 59971 529896
rect 52913 529891 52979 529894
rect 59905 529891 59971 529894
rect 55673 529820 55739 529821
rect 55622 529818 55628 529820
rect 55582 529758 55628 529818
rect 55692 529816 55739 529820
rect 55734 529760 55739 529816
rect 55622 529756 55628 529758
rect 55692 529756 55739 529760
rect 55673 529755 55739 529756
rect 59905 529818 59971 529821
rect 292665 529818 292731 529821
rect 59905 529816 292731 529818
rect 59905 529760 59910 529816
rect 59966 529760 292670 529816
rect 292726 529760 292731 529816
rect 59905 529758 292731 529760
rect 59905 529755 59971 529758
rect 292665 529755 292731 529758
rect 127249 529682 127315 529685
rect 236361 529682 236427 529685
rect 127249 529680 236427 529682
rect 127249 529624 127254 529680
rect 127310 529624 236366 529680
rect 236422 529624 236427 529680
rect 127249 529622 236427 529624
rect 127249 529619 127315 529622
rect 236361 529619 236427 529622
rect 242249 529682 242315 529685
rect 486509 529682 486575 529685
rect 242249 529680 486575 529682
rect 242249 529624 242254 529680
rect 242310 529624 486514 529680
rect 486570 529624 486575 529680
rect 242249 529622 486575 529624
rect 242249 529619 242315 529622
rect 486509 529619 486575 529622
rect 51717 529546 51783 529549
rect 334893 529546 334959 529549
rect 51717 529544 334959 529546
rect 51717 529488 51722 529544
rect 51778 529488 334898 529544
rect 334954 529488 334959 529544
rect 51717 529486 334959 529488
rect 51717 529483 51783 529486
rect 334893 529483 334959 529486
rect 57830 529348 57836 529412
rect 57900 529410 57906 529412
rect 166257 529410 166323 529413
rect 57900 529408 166323 529410
rect 57900 529352 166262 529408
rect 166318 529352 166323 529408
rect 57900 529350 166323 529352
rect 57900 529348 57906 529350
rect 166257 529347 166323 529350
rect 177062 529348 177068 529412
rect 177132 529410 177138 529412
rect 177481 529410 177547 529413
rect 177132 529408 177547 529410
rect 177132 529352 177486 529408
rect 177542 529352 177547 529408
rect 177132 529350 177547 529352
rect 177132 529348 177138 529350
rect 177481 529347 177547 529350
rect 288382 529348 288388 529412
rect 288452 529410 288458 529412
rect 289721 529410 289787 529413
rect 288452 529408 289787 529410
rect 288452 529352 289726 529408
rect 289782 529352 289787 529408
rect 288452 529350 289787 529352
rect 288452 529348 288458 529350
rect 289721 529347 289787 529350
rect 59077 529274 59143 529277
rect 376845 529274 376911 529277
rect 59077 529272 376911 529274
rect 59077 529216 59082 529272
rect 59138 529216 376850 529272
rect 376906 529216 376911 529272
rect 59077 529214 376911 529216
rect 59077 529211 59143 529214
rect 376845 529211 376911 529214
rect 57421 529138 57487 529141
rect 59445 529138 59511 529141
rect 377622 529138 377628 529140
rect 57421 529136 59511 529138
rect 57421 529080 57426 529136
rect 57482 529080 59450 529136
rect 59506 529080 59511 529136
rect 57421 529078 59511 529080
rect 57421 529075 57487 529078
rect 59445 529075 59511 529078
rect 64830 529078 377628 529138
rect 55990 528940 55996 529004
rect 56060 529002 56066 529004
rect 64830 529002 64890 529078
rect 377622 529076 377628 529078
rect 377692 529076 377698 529140
rect 56060 528942 64890 529002
rect 134517 529002 134583 529005
rect 325509 529002 325575 529005
rect 134517 529000 325575 529002
rect 134517 528944 134522 529000
rect 134578 528944 325514 529000
rect 325570 528944 325575 529000
rect 134517 528942 325575 528944
rect 56060 528940 56066 528942
rect 134517 528939 134583 528942
rect 325509 528939 325575 528942
rect 57789 528866 57855 528869
rect 127617 528866 127683 528869
rect 57789 528864 127683 528866
rect 57789 528808 57794 528864
rect 57850 528808 127622 528864
rect 127678 528808 127683 528864
rect 57789 528806 127683 528808
rect 57789 528803 57855 528806
rect 127617 528803 127683 528806
rect 51533 528730 51599 528733
rect 59169 528730 59235 528733
rect 135161 528730 135227 528733
rect 51533 528728 59235 528730
rect 51533 528672 51538 528728
rect 51594 528672 59174 528728
rect 59230 528672 59235 528728
rect 51533 528670 59235 528672
rect 51533 528667 51599 528670
rect 59169 528667 59235 528670
rect 64830 528728 135227 528730
rect 64830 528672 135166 528728
rect 135222 528672 135227 528728
rect 64830 528670 135227 528672
rect 56869 528594 56935 528597
rect 64830 528594 64890 528670
rect 135161 528667 135227 528670
rect 166257 528730 166323 528733
rect 460013 528730 460079 528733
rect 166257 528728 460079 528730
rect 166257 528672 166262 528728
rect 166318 528672 460018 528728
rect 460074 528672 460079 528728
rect 166257 528670 460079 528672
rect 166257 528667 166323 528670
rect 460013 528667 460079 528670
rect 56869 528592 64890 528594
rect 56869 528536 56874 528592
rect 56930 528536 64890 528592
rect 56869 528534 64890 528536
rect 56869 528531 56935 528534
rect 155309 528458 155375 528461
rect 334893 528458 334959 528461
rect 155309 528456 334959 528458
rect 155309 528400 155314 528456
rect 155370 528400 334898 528456
rect 334954 528400 334959 528456
rect 155309 528398 334959 528400
rect 155309 528395 155375 528398
rect 334893 528395 334959 528398
rect 174721 528322 174787 528325
rect 411529 528322 411595 528325
rect 174721 528320 411595 528322
rect 174721 528264 174726 528320
rect 174782 528264 411534 528320
rect 411590 528264 411595 528320
rect 174721 528262 411595 528264
rect 174721 528259 174787 528262
rect 411529 528259 411595 528262
rect 170397 528186 170463 528189
rect 425605 528186 425671 528189
rect 170397 528184 425671 528186
rect 170397 528128 170402 528184
rect 170458 528128 425610 528184
rect 425666 528128 425671 528184
rect 170397 528126 425671 528128
rect 170397 528123 170463 528126
rect 425605 528123 425671 528126
rect 169201 528050 169267 528053
rect 441245 528050 441311 528053
rect 169201 528048 441311 528050
rect -960 527914 480 528004
rect 169201 527992 169206 528048
rect 169262 527992 441250 528048
rect 441306 527992 441311 528048
rect 169201 527990 441311 527992
rect 169201 527987 169267 527990
rect 441245 527987 441311 527990
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 164877 527914 164943 527917
rect 169753 527914 169819 527917
rect 164877 527912 169819 527914
rect 164877 527856 164882 527912
rect 164938 527856 169758 527912
rect 169814 527856 169819 527912
rect 164877 527854 169819 527856
rect 164877 527851 164943 527854
rect 169753 527851 169819 527854
rect 219985 527914 220051 527917
rect 498561 527914 498627 527917
rect 219985 527912 498627 527914
rect 219985 527856 219990 527912
rect 220046 527856 498566 527912
rect 498622 527856 498627 527912
rect 219985 527854 498627 527856
rect 219985 527851 220051 527854
rect 498561 527851 498627 527854
rect 175774 527716 175780 527780
rect 175844 527778 175850 527780
rect 458449 527778 458515 527781
rect 175844 527776 458515 527778
rect 175844 527720 458454 527776
rect 458510 527720 458515 527776
rect 175844 527718 458515 527720
rect 175844 527716 175850 527718
rect 458449 527715 458515 527718
rect 57513 527642 57579 527645
rect 175181 527642 175247 527645
rect 57513 527640 175247 527642
rect 57513 527584 57518 527640
rect 57574 527584 175186 527640
rect 175242 527584 175247 527640
rect 57513 527582 175247 527584
rect 57513 527579 57579 527582
rect 175181 527579 175247 527582
rect 285622 527580 285628 527644
rect 285692 527642 285698 527644
rect 286317 527642 286383 527645
rect 326981 527642 327047 527645
rect 285692 527640 286383 527642
rect 285692 527584 286322 527640
rect 286378 527584 286383 527640
rect 285692 527582 286383 527584
rect 285692 527580 285698 527582
rect 286317 527579 286383 527582
rect 287010 527640 327047 527642
rect 287010 527584 326986 527640
rect 327042 527584 327047 527640
rect 287010 527582 327047 527584
rect 57881 527506 57947 527509
rect 175825 527506 175891 527509
rect 57881 527504 175891 527506
rect 57881 527448 57886 527504
rect 57942 527448 175830 527504
rect 175886 527448 175891 527504
rect 57881 527446 175891 527448
rect 57881 527443 57947 527446
rect 175825 527443 175891 527446
rect 279417 527506 279483 527509
rect 287010 527506 287070 527582
rect 326981 527579 327047 527582
rect 279417 527504 287070 527506
rect 279417 527448 279422 527504
rect 279478 527448 287070 527504
rect 279417 527446 287070 527448
rect 279417 527443 279483 527446
rect 32857 527370 32923 527373
rect 220629 527370 220695 527373
rect 32857 527368 220695 527370
rect 32857 527312 32862 527368
rect 32918 527312 220634 527368
rect 220690 527312 220695 527368
rect 32857 527310 220695 527312
rect 32857 527307 32923 527310
rect 220629 527307 220695 527310
rect 36486 527172 36492 527236
rect 36556 527234 36562 527236
rect 279969 527234 280035 527237
rect 36556 527232 280035 527234
rect 36556 527176 279974 527232
rect 280030 527176 280035 527232
rect 36556 527174 280035 527176
rect 36556 527172 36562 527174
rect 279969 527171 280035 527174
rect 103973 527098 104039 527101
rect 200389 527098 200455 527101
rect 103973 527096 200455 527098
rect 103973 527040 103978 527096
rect 104034 527040 200394 527096
rect 200450 527040 200455 527096
rect 103973 527038 200455 527040
rect 103973 527035 104039 527038
rect 200389 527035 200455 527038
rect 286869 527098 286935 527101
rect 289721 527098 289787 527101
rect 286869 527096 289787 527098
rect 286869 527040 286874 527096
rect 286930 527040 289726 527096
rect 289782 527040 289787 527096
rect 286869 527038 289787 527040
rect 286869 527035 286935 527038
rect 289721 527035 289787 527038
rect 105997 526962 106063 526965
rect 203517 526962 203583 526965
rect 105997 526960 203583 526962
rect 105997 526904 106002 526960
rect 106058 526904 203522 526960
rect 203578 526904 203583 526960
rect 105997 526902 203583 526904
rect 105997 526899 106063 526902
rect 203517 526899 203583 526902
rect 246297 526962 246363 526965
rect 486601 526962 486667 526965
rect 246297 526960 486667 526962
rect 246297 526904 246302 526960
rect 246358 526904 486606 526960
rect 486662 526904 486667 526960
rect 246297 526902 486667 526904
rect 246297 526899 246363 526902
rect 486601 526899 486667 526902
rect 107009 526826 107075 526829
rect 205081 526826 205147 526829
rect 107009 526824 205147 526826
rect 107009 526768 107014 526824
rect 107070 526768 205086 526824
rect 205142 526768 205147 526824
rect 107009 526766 205147 526768
rect 107009 526763 107075 526766
rect 205081 526763 205147 526766
rect 235165 526826 235231 526829
rect 484853 526826 484919 526829
rect 235165 526824 484919 526826
rect 235165 526768 235170 526824
rect 235226 526768 484858 526824
rect 484914 526768 484919 526824
rect 235165 526766 484919 526768
rect 235165 526763 235231 526766
rect 484853 526763 484919 526766
rect 108021 526690 108087 526693
rect 206645 526690 206711 526693
rect 108021 526688 206711 526690
rect 108021 526632 108026 526688
rect 108082 526632 206650 526688
rect 206706 526632 206711 526688
rect 108021 526630 206711 526632
rect 108021 526627 108087 526630
rect 206645 526627 206711 526630
rect 222009 526690 222075 526693
rect 483238 526690 483244 526692
rect 222009 526688 483244 526690
rect 222009 526632 222014 526688
rect 222070 526632 483244 526688
rect 222009 526630 483244 526632
rect 222009 526627 222075 526630
rect 483238 526628 483244 526630
rect 483308 526628 483314 526692
rect 109309 526554 109375 526557
rect 208209 526554 208275 526557
rect 109309 526552 208275 526554
rect 109309 526496 109314 526552
rect 109370 526496 208214 526552
rect 208270 526496 208275 526552
rect 109309 526494 208275 526496
rect 109309 526491 109375 526494
rect 208209 526491 208275 526494
rect 214925 526554 214991 526557
rect 491569 526554 491635 526557
rect 214925 526552 491635 526554
rect 214925 526496 214930 526552
rect 214986 526496 491574 526552
rect 491630 526496 491635 526552
rect 214925 526494 491635 526496
rect 214925 526491 214991 526494
rect 491569 526491 491635 526494
rect 46289 526418 46355 526421
rect 107561 526418 107627 526421
rect 46289 526416 107627 526418
rect 46289 526360 46294 526416
rect 46350 526360 107566 526416
rect 107622 526360 107627 526416
rect 46289 526358 107627 526360
rect 46289 526355 46355 526358
rect 107561 526355 107627 526358
rect 110045 526418 110111 526421
rect 209681 526418 209747 526421
rect 110045 526416 209747 526418
rect 110045 526360 110050 526416
rect 110106 526360 209686 526416
rect 209742 526360 209747 526416
rect 110045 526358 209747 526360
rect 110045 526355 110111 526358
rect 209681 526355 209747 526358
rect 217961 526418 218027 526421
rect 495617 526418 495683 526421
rect 217961 526416 495683 526418
rect 217961 526360 217966 526416
rect 218022 526360 495622 526416
rect 495678 526360 495683 526416
rect 217961 526358 495683 526360
rect 217961 526355 218027 526358
rect 495617 526355 495683 526358
rect 105077 526282 105143 526285
rect 201953 526282 202019 526285
rect 105077 526280 202019 526282
rect 105077 526224 105082 526280
rect 105138 526224 201958 526280
rect 202014 526224 202019 526280
rect 105077 526222 202019 526224
rect 105077 526219 105143 526222
rect 201953 526219 202019 526222
rect 299790 526220 299796 526284
rect 299860 526282 299866 526284
rect 503662 526282 503668 526284
rect 299860 526222 503668 526282
rect 299860 526220 299866 526222
rect 503662 526220 503668 526222
rect 503732 526220 503738 526284
rect 43805 526146 43871 526149
rect 109033 526146 109099 526149
rect 43805 526144 109099 526146
rect 43805 526088 43810 526144
rect 43866 526088 109038 526144
rect 109094 526088 109099 526144
rect 43805 526086 109099 526088
rect 43805 526083 43871 526086
rect 109033 526083 109099 526086
rect 171542 526084 171548 526148
rect 171612 526146 171618 526148
rect 172421 526146 172487 526149
rect 171612 526144 172487 526146
rect 171612 526088 172426 526144
rect 172482 526088 172487 526144
rect 171612 526086 172487 526088
rect 171612 526084 171618 526086
rect 172421 526083 172487 526086
rect 201769 526146 201835 526149
rect 300761 526146 300827 526149
rect 201769 526144 300827 526146
rect 201769 526088 201774 526144
rect 201830 526088 300766 526144
rect 300822 526088 300827 526144
rect 201769 526086 300827 526088
rect 201769 526083 201835 526086
rect 300761 526083 300827 526086
rect 40585 526010 40651 526013
rect 108297 526010 108363 526013
rect 40585 526008 108363 526010
rect 40585 525952 40590 526008
rect 40646 525952 108302 526008
rect 108358 525952 108363 526008
rect 40585 525950 108363 525952
rect 40585 525947 40651 525950
rect 108297 525947 108363 525950
rect 288934 525948 288940 526012
rect 289004 526010 289010 526012
rect 493174 526010 493180 526012
rect 289004 525950 493180 526010
rect 289004 525948 289010 525950
rect 493174 525948 493180 525950
rect 493244 525948 493250 526012
rect 37222 525812 37228 525876
rect 37292 525874 37298 525876
rect 109125 525874 109191 525877
rect 37292 525872 109191 525874
rect 37292 525816 109130 525872
rect 109186 525816 109191 525872
rect 37292 525814 109191 525816
rect 37292 525812 37298 525814
rect 109125 525811 109191 525814
rect 175038 525676 175044 525740
rect 175108 525738 175114 525740
rect 175181 525738 175247 525741
rect 175108 525736 175247 525738
rect 175108 525680 175186 525736
rect 175242 525680 175247 525736
rect 175108 525678 175247 525680
rect 175108 525676 175114 525678
rect 175181 525675 175247 525678
rect 179822 525676 179828 525740
rect 179892 525738 179898 525740
rect 180241 525738 180307 525741
rect 179892 525736 180307 525738
rect 179892 525680 180246 525736
rect 180302 525680 180307 525736
rect 179892 525678 180307 525680
rect 179892 525676 179898 525678
rect 180241 525675 180307 525678
rect 295926 525676 295932 525740
rect 295996 525738 296002 525740
rect 497038 525738 497044 525740
rect 295996 525678 497044 525738
rect 295996 525676 296002 525678
rect 497038 525676 497044 525678
rect 497108 525676 497114 525740
rect 101949 525602 102015 525605
rect 197261 525602 197327 525605
rect 101949 525600 197327 525602
rect 101949 525544 101954 525600
rect 102010 525544 197266 525600
rect 197322 525544 197327 525600
rect 101949 525542 197327 525544
rect 101949 525539 102015 525542
rect 197261 525539 197327 525542
rect 294454 525540 294460 525604
rect 294524 525602 294530 525604
rect 507894 525602 507900 525604
rect 294524 525542 507900 525602
rect 294524 525540 294530 525542
rect 507894 525540 507900 525542
rect 507964 525540 507970 525604
rect 176101 525466 176167 525469
rect 402145 525466 402211 525469
rect 176101 525464 402211 525466
rect 176101 525408 176106 525464
rect 176162 525408 402150 525464
rect 402206 525408 402211 525464
rect 176101 525406 402211 525408
rect 176101 525403 176167 525406
rect 402145 525403 402211 525406
rect 43713 525330 43779 525333
rect 102133 525330 102199 525333
rect 43713 525328 102199 525330
rect 43713 525272 43718 525328
rect 43774 525272 102138 525328
rect 102194 525272 102199 525328
rect 43713 525270 102199 525272
rect 43713 525267 43779 525270
rect 102133 525267 102199 525270
rect 102961 525330 103027 525333
rect 198825 525330 198891 525333
rect 102961 525328 198891 525330
rect 102961 525272 102966 525328
rect 103022 525272 198830 525328
rect 198886 525272 198891 525328
rect 102961 525270 198891 525272
rect 102961 525267 103027 525270
rect 198825 525267 198891 525270
rect 244273 525330 244339 525333
rect 485037 525330 485103 525333
rect 244273 525328 485103 525330
rect 244273 525272 244278 525328
rect 244334 525272 485042 525328
rect 485098 525272 485103 525328
rect 244273 525270 485103 525272
rect 244273 525267 244339 525270
rect 485037 525267 485103 525270
rect 42149 525194 42215 525197
rect 100753 525194 100819 525197
rect 42149 525192 100819 525194
rect 42149 525136 42154 525192
rect 42210 525136 100758 525192
rect 100814 525136 100819 525192
rect 42149 525134 100819 525136
rect 42149 525131 42215 525134
rect 100753 525131 100819 525134
rect 119153 525194 119219 525197
rect 223849 525194 223915 525197
rect 119153 525192 223915 525194
rect 119153 525136 119158 525192
rect 119214 525136 223854 525192
rect 223910 525136 223915 525192
rect 119153 525134 223915 525136
rect 119153 525131 119219 525134
rect 223849 525131 223915 525134
rect 231117 525194 231183 525197
rect 489177 525194 489243 525197
rect 231117 525192 489243 525194
rect 231117 525136 231122 525192
rect 231178 525136 489182 525192
rect 489238 525136 489243 525192
rect 231117 525134 489243 525136
rect 231117 525131 231183 525134
rect 489177 525131 489243 525134
rect 51625 525058 51691 525061
rect 120073 525058 120139 525061
rect 51625 525056 120139 525058
rect 51625 525000 51630 525056
rect 51686 525000 120078 525056
rect 120134 525000 120139 525056
rect 51625 524998 120139 525000
rect 51625 524995 51691 524998
rect 120073 524995 120139 524998
rect 121177 525058 121243 525061
rect 226977 525058 227043 525061
rect 121177 525056 227043 525058
rect 121177 525000 121182 525056
rect 121238 525000 226982 525056
rect 227038 525000 227043 525056
rect 121177 524998 227043 525000
rect 121177 524995 121243 524998
rect 226977 524995 227043 524998
rect 234153 525058 234219 525061
rect 501229 525058 501295 525061
rect 234153 525056 501295 525058
rect 234153 525000 234158 525056
rect 234214 525000 501234 525056
rect 501290 525000 501295 525056
rect 234153 524998 501295 525000
rect 234153 524995 234219 524998
rect 501229 524995 501295 524998
rect 43621 524922 43687 524925
rect 118693 524922 118759 524925
rect 43621 524920 118759 524922
rect 43621 524864 43626 524920
rect 43682 524864 118698 524920
rect 118754 524864 118759 524920
rect 43621 524862 118759 524864
rect 43621 524859 43687 524862
rect 118693 524859 118759 524862
rect 133321 524922 133387 524925
rect 211061 524922 211127 524925
rect 133321 524920 211127 524922
rect 133321 524864 133326 524920
rect 133382 524864 211066 524920
rect 211122 524864 211127 524920
rect 133321 524862 211127 524864
rect 133321 524859 133387 524862
rect 211061 524859 211127 524862
rect 299238 524860 299244 524924
rect 299308 524922 299314 524924
rect 499982 524922 499988 524924
rect 299308 524862 499988 524922
rect 299308 524860 299314 524862
rect 499982 524860 499988 524862
rect 500052 524860 500058 524924
rect 40861 524786 40927 524789
rect 133781 524786 133847 524789
rect 40861 524784 133847 524786
rect 40861 524728 40866 524784
rect 40922 524728 133786 524784
rect 133842 524728 133847 524784
rect 40861 524726 133847 524728
rect 40861 524723 40927 524726
rect 133781 524723 133847 524726
rect 44633 524650 44699 524653
rect 175917 524650 175983 524653
rect 44633 524648 175983 524650
rect 44633 524592 44638 524648
rect 44694 524592 175922 524648
rect 175978 524592 175983 524648
rect 44633 524590 175983 524592
rect 44633 524587 44699 524590
rect 175917 524587 175983 524590
rect 32949 524514 33015 524517
rect 299381 524514 299447 524517
rect 32949 524512 299447 524514
rect 32949 524456 32954 524512
rect 33010 524456 299386 524512
rect 299442 524456 299447 524512
rect 32949 524454 299447 524456
rect 32949 524451 33015 524454
rect 299381 524451 299447 524454
rect 547086 524452 547092 524516
rect 547156 524514 547162 524516
rect 583520 524514 584960 524604
rect 547156 524454 584960 524514
rect 547156 524452 547162 524454
rect 137553 524378 137619 524381
rect 324313 524378 324379 524381
rect 137553 524376 324379 524378
rect 137553 524320 137558 524376
rect 137614 524320 324318 524376
rect 324374 524320 324379 524376
rect 137553 524318 324379 524320
rect 137553 524315 137619 524318
rect 324313 524315 324379 524318
rect 471605 524378 471671 524381
rect 473353 524378 473419 524381
rect 471605 524376 473419 524378
rect 471605 524320 471610 524376
rect 471666 524320 473358 524376
rect 473414 524320 473419 524376
rect 583520 524364 584960 524454
rect 471605 524318 473419 524320
rect 471605 524315 471671 524318
rect 473353 524315 473419 524318
rect 56961 524242 57027 524245
rect 63493 524242 63559 524245
rect 56961 524240 63559 524242
rect 56961 524184 56966 524240
rect 57022 524184 63498 524240
rect 63554 524184 63559 524240
rect 56961 524182 63559 524184
rect 56961 524179 57027 524182
rect 63493 524179 63559 524182
rect 170765 524242 170831 524245
rect 377121 524242 377187 524245
rect 170765 524240 377187 524242
rect 170765 524184 170770 524240
rect 170826 524184 377126 524240
rect 377182 524184 377187 524240
rect 170765 524182 377187 524184
rect 170765 524179 170831 524182
rect 377121 524179 377187 524182
rect 35198 524044 35204 524108
rect 35268 524106 35274 524108
rect 66161 524106 66227 524109
rect 35268 524104 66227 524106
rect 35268 524048 66166 524104
rect 66222 524048 66227 524104
rect 35268 524046 66227 524048
rect 35268 524044 35274 524046
rect 66161 524043 66227 524046
rect 69565 524106 69631 524109
rect 137737 524106 137803 524109
rect 69565 524104 137803 524106
rect 69565 524048 69570 524104
rect 69626 524048 137742 524104
rect 137798 524048 137803 524104
rect 69565 524046 137803 524048
rect 69565 524043 69631 524046
rect 137737 524043 137803 524046
rect 178769 524106 178835 524109
rect 392761 524106 392827 524109
rect 178769 524104 392827 524106
rect 178769 524048 178774 524104
rect 178830 524048 392766 524104
rect 392822 524048 392827 524104
rect 178769 524046 392827 524048
rect 178769 524043 178835 524046
rect 392761 524043 392827 524046
rect 59169 523970 59235 523973
rect 45510 523968 59235 523970
rect 45510 523912 59174 523968
rect 59230 523912 59235 523968
rect 45510 523910 59235 523912
rect 42241 523834 42307 523837
rect 45510 523834 45570 523910
rect 59169 523907 59235 523910
rect 64505 523970 64571 523973
rect 130009 523970 130075 523973
rect 64505 523968 130075 523970
rect 64505 523912 64510 523968
rect 64566 523912 130014 523968
rect 130070 523912 130075 523968
rect 64505 523910 130075 523912
rect 64505 523907 64571 523910
rect 130009 523907 130075 523910
rect 130285 523970 130351 523973
rect 241053 523970 241119 523973
rect 130285 523968 241119 523970
rect 130285 523912 130290 523968
rect 130346 523912 241058 523968
rect 241114 523912 241119 523968
rect 130285 523910 241119 523912
rect 130285 523907 130351 523910
rect 241053 523907 241119 523910
rect 257981 523970 258047 523973
rect 485221 523970 485287 523973
rect 257981 523968 485287 523970
rect 257981 523912 257986 523968
rect 258042 523912 485226 523968
rect 485282 523912 485287 523968
rect 257981 523910 485287 523912
rect 257981 523907 258047 523910
rect 485221 523907 485287 523910
rect 42241 523832 45570 523834
rect 42241 523776 42246 523832
rect 42302 523776 45570 523832
rect 42241 523774 45570 523776
rect 57973 523834 58039 523837
rect 58566 523834 58572 523836
rect 57973 523832 58572 523834
rect 57973 523776 57978 523832
rect 58034 523776 58572 523832
rect 57973 523774 58572 523776
rect 42241 523771 42307 523774
rect 57973 523771 58039 523774
rect 58566 523772 58572 523774
rect 58636 523772 58642 523836
rect 65517 523834 65583 523837
rect 131573 523834 131639 523837
rect 65517 523832 131639 523834
rect 65517 523776 65522 523832
rect 65578 523776 131578 523832
rect 131634 523776 131639 523832
rect 65517 523774 131639 523776
rect 65517 523771 65583 523774
rect 131573 523771 131639 523774
rect 137369 523834 137435 523837
rect 367001 523834 367067 523837
rect 137369 523832 367067 523834
rect 137369 523776 137374 523832
rect 137430 523776 367006 523832
rect 367062 523776 367067 523832
rect 137369 523774 367067 523776
rect 137369 523771 137435 523774
rect 367001 523771 367067 523774
rect 39614 523636 39620 523700
rect 39684 523698 39690 523700
rect 280838 523698 280844 523700
rect 39684 523638 280844 523698
rect 39684 523636 39690 523638
rect 280838 523636 280844 523638
rect 280908 523636 280914 523700
rect 293861 523698 293927 523701
rect 482185 523698 482251 523701
rect 293861 523696 482251 523698
rect 293861 523640 293866 523696
rect 293922 523640 482190 523696
rect 482246 523640 482251 523696
rect 293861 523638 482251 523640
rect 293861 523635 293927 523638
rect 482185 523635 482251 523638
rect 42057 523562 42123 523565
rect 69657 523562 69723 523565
rect 42057 523560 69723 523562
rect 42057 523504 42062 523560
rect 42118 523504 69662 523560
rect 69718 523504 69723 523560
rect 42057 523502 69723 523504
rect 42057 523499 42123 523502
rect 69657 523499 69723 523502
rect 275185 523562 275251 523565
rect 292573 523562 292639 523565
rect 275185 523560 292639 523562
rect 275185 523504 275190 523560
rect 275246 523504 292578 523560
rect 292634 523504 292639 523560
rect 275185 523502 292639 523504
rect 275185 523499 275251 523502
rect 292573 523499 292639 523502
rect 299289 523562 299355 523565
rect 482553 523562 482619 523565
rect 299289 523560 482619 523562
rect 299289 523504 299294 523560
rect 299350 523504 482558 523560
rect 482614 523504 482619 523560
rect 299289 523502 482619 523504
rect 299289 523499 299355 523502
rect 482553 523499 482619 523502
rect 36670 523364 36676 523428
rect 36740 523426 36746 523428
rect 169753 523426 169819 523429
rect 36740 523424 169819 523426
rect 36740 523368 169758 523424
rect 169814 523368 169819 523424
rect 36740 523366 169819 523368
rect 36740 523364 36746 523366
rect 169753 523363 169819 523366
rect 292481 523426 292547 523429
rect 299381 523426 299447 523429
rect 292481 523424 299447 523426
rect 292481 523368 292486 523424
rect 292542 523368 299386 523424
rect 299442 523368 299447 523424
rect 292481 523366 299447 523368
rect 292481 523363 292547 523366
rect 299381 523363 299447 523366
rect 38101 523290 38167 523293
rect 178033 523290 178099 523293
rect 38101 523288 178099 523290
rect 38101 523232 38106 523288
rect 38162 523232 178038 523288
rect 178094 523232 178099 523288
rect 38101 523230 178099 523232
rect 38101 523227 38167 523230
rect 178033 523227 178099 523230
rect 58382 523092 58388 523156
rect 58452 523154 58458 523156
rect 274633 523154 274699 523157
rect 58452 523152 274699 523154
rect 58452 523096 274638 523152
rect 274694 523096 274699 523152
rect 58452 523094 274699 523096
rect 58452 523092 58458 523094
rect 274633 523091 274699 523094
rect 481633 523154 481699 523157
rect 482318 523154 482324 523156
rect 481633 523152 482324 523154
rect 481633 523096 481638 523152
rect 481694 523096 482324 523152
rect 481633 523094 482324 523096
rect 481633 523091 481699 523094
rect 482318 523092 482324 523094
rect 482388 523092 482394 523156
rect 55765 523020 55831 523021
rect 59537 523020 59603 523021
rect 55765 523018 55812 523020
rect 55720 523016 55812 523018
rect 55720 522960 55770 523016
rect 55720 522958 55812 522960
rect 55765 522956 55812 522958
rect 55876 522956 55882 523020
rect 59486 523018 59492 523020
rect 59446 522958 59492 523018
rect 59556 523016 59603 523020
rect 59598 522960 59603 523016
rect 59486 522956 59492 522958
rect 59556 522956 59603 522960
rect 55765 522955 55831 522956
rect 59537 522955 59603 522956
rect 62481 523018 62547 523021
rect 126881 523018 126947 523021
rect 62481 523016 126947 523018
rect 62481 522960 62486 523016
rect 62542 522960 126886 523016
rect 126942 522960 126947 523016
rect 62481 522958 126947 522960
rect 62481 522955 62547 522958
rect 126881 522955 126947 522958
rect 174537 523018 174603 523021
rect 176929 523018 176995 523021
rect 174537 523016 176995 523018
rect 174537 522960 174542 523016
rect 174598 522960 176934 523016
rect 176990 522960 176995 523016
rect 174537 522958 176995 522960
rect 174537 522955 174603 522958
rect 176929 522955 176995 522958
rect 177573 523018 177639 523021
rect 471881 523018 471947 523021
rect 177573 523016 471947 523018
rect 177573 522960 177578 523016
rect 177634 522960 471886 523016
rect 471942 522960 471947 523016
rect 177573 522958 471947 522960
rect 177573 522955 177639 522958
rect 471881 522955 471947 522958
rect 63677 522882 63743 522885
rect 128445 522882 128511 522885
rect 63677 522880 128511 522882
rect 63677 522824 63682 522880
rect 63738 522824 128450 522880
rect 128506 522824 128511 522880
rect 63677 522822 128511 522824
rect 63677 522819 63743 522822
rect 128445 522819 128511 522822
rect 257102 522820 257108 522884
rect 257172 522882 257178 522884
rect 480294 522882 480300 522884
rect 257172 522822 480300 522882
rect 257172 522820 257178 522822
rect 480294 522820 480300 522822
rect 480364 522820 480370 522884
rect 40493 522746 40559 522749
rect 63493 522746 63559 522749
rect 40493 522744 63559 522746
rect 40493 522688 40498 522744
rect 40554 522688 63498 522744
rect 63554 522688 63559 522744
rect 40493 522686 63559 522688
rect 40493 522683 40559 522686
rect 63493 522683 63559 522686
rect 80697 522746 80763 522749
rect 155033 522746 155099 522749
rect 80697 522744 155099 522746
rect 80697 522688 80702 522744
rect 80758 522688 155038 522744
rect 155094 522688 155099 522744
rect 80697 522686 155099 522688
rect 80697 522683 80763 522686
rect 155033 522683 155099 522686
rect 176009 522746 176075 522749
rect 405273 522746 405339 522749
rect 176009 522744 405339 522746
rect 176009 522688 176014 522744
rect 176070 522688 405278 522744
rect 405334 522688 405339 522744
rect 176009 522686 405339 522688
rect 176009 522683 176075 522686
rect 405273 522683 405339 522686
rect 464613 522746 464679 522749
rect 501321 522746 501387 522749
rect 464613 522744 501387 522746
rect 464613 522688 464618 522744
rect 464674 522688 501326 522744
rect 501382 522688 501387 522744
rect 464613 522686 501387 522688
rect 464613 522683 464679 522686
rect 501321 522683 501387 522686
rect 43662 522548 43668 522612
rect 43732 522610 43738 522612
rect 56501 522610 56567 522613
rect 43732 522608 56567 522610
rect 43732 522552 56506 522608
rect 56562 522552 56567 522608
rect 43732 522550 56567 522552
rect 43732 522548 43738 522550
rect 56501 522547 56567 522550
rect 59854 522548 59860 522612
rect 59924 522610 59930 522612
rect 297357 522610 297423 522613
rect 59924 522608 297423 522610
rect 59924 522552 297362 522608
rect 297418 522552 297423 522608
rect 59924 522550 297423 522552
rect 59924 522548 59930 522550
rect 297357 522547 297423 522550
rect 464337 522610 464403 522613
rect 502701 522610 502767 522613
rect 464337 522608 502767 522610
rect 464337 522552 464342 522608
rect 464398 522552 502706 522608
rect 502762 522552 502767 522608
rect 464337 522550 502767 522552
rect 464337 522547 464403 522550
rect 502701 522547 502767 522550
rect 55990 522412 55996 522476
rect 56060 522474 56066 522476
rect 296846 522474 296852 522476
rect 56060 522414 296852 522474
rect 56060 522412 56066 522414
rect 296846 522412 296852 522414
rect 296916 522412 296922 522476
rect 298686 522412 298692 522476
rect 298756 522474 298762 522476
rect 495566 522474 495572 522476
rect 298756 522414 495572 522474
rect 298756 522412 298762 522414
rect 495566 522412 495572 522414
rect 495636 522412 495642 522476
rect 34094 522276 34100 522340
rect 34164 522338 34170 522340
rect 280654 522338 280660 522340
rect 34164 522278 280660 522338
rect 34164 522276 34170 522278
rect 280654 522276 280660 522278
rect 280724 522276 280730 522340
rect 295149 522338 295215 522341
rect 496813 522338 496879 522341
rect 295149 522336 496879 522338
rect 295149 522280 295154 522336
rect 295210 522280 496818 522336
rect 496874 522280 496879 522336
rect 295149 522278 496879 522280
rect 295149 522275 295215 522278
rect 496813 522275 496879 522278
rect 35382 522140 35388 522204
rect 35452 522202 35458 522204
rect 62113 522202 62179 522205
rect 35452 522200 62179 522202
rect 35452 522144 62118 522200
rect 62174 522144 62179 522200
rect 35452 522142 62179 522144
rect 35452 522140 35458 522142
rect 62113 522139 62179 522142
rect 114093 522202 114159 522205
rect 175917 522202 175983 522205
rect 114093 522200 175983 522202
rect 114093 522144 114098 522200
rect 114154 522144 175922 522200
rect 175978 522144 175983 522200
rect 114093 522142 175983 522144
rect 114093 522139 114159 522142
rect 175917 522139 175983 522142
rect 177665 522202 177731 522205
rect 293953 522202 294019 522205
rect 177665 522200 294019 522202
rect 177665 522144 177670 522200
rect 177726 522144 293958 522200
rect 294014 522144 294019 522200
rect 177665 522142 294019 522144
rect 177665 522139 177731 522142
rect 293953 522139 294019 522142
rect 295241 522202 295307 522205
rect 482369 522202 482435 522205
rect 295241 522200 482435 522202
rect 295241 522144 295246 522200
rect 295302 522144 482374 522200
rect 482430 522144 482435 522200
rect 295241 522142 482435 522144
rect 295241 522139 295307 522142
rect 482369 522139 482435 522142
rect 31385 522066 31451 522069
rect 59905 522066 59971 522069
rect 31385 522064 59971 522066
rect 31385 522008 31390 522064
rect 31446 522008 59910 522064
rect 59966 522008 59971 522064
rect 31385 522006 59971 522008
rect 31385 522003 31451 522006
rect 59905 522003 59971 522006
rect 471513 522066 471579 522069
rect 498745 522066 498811 522069
rect 471513 522064 498811 522066
rect 471513 522008 471518 522064
rect 471574 522008 498750 522064
rect 498806 522008 498811 522064
rect 471513 522006 498811 522008
rect 471513 522003 471579 522006
rect 498745 522003 498811 522006
rect 46105 521930 46171 521933
rect 80053 521930 80119 521933
rect 46105 521928 80119 521930
rect 46105 521872 46110 521928
rect 46166 521872 80058 521928
rect 80114 521872 80119 521928
rect 46105 521870 80119 521872
rect 46105 521867 46171 521870
rect 80053 521867 80119 521870
rect 39246 521732 39252 521796
rect 39316 521794 39322 521796
rect 114461 521794 114527 521797
rect 39316 521792 114527 521794
rect 39316 521736 114466 521792
rect 114522 521736 114527 521792
rect 39316 521734 114527 521736
rect 39316 521732 39322 521734
rect 114461 521731 114527 521734
rect 58934 521596 58940 521660
rect 59004 521658 59010 521660
rect 59077 521658 59143 521661
rect 59004 521656 59143 521658
rect 59004 521600 59082 521656
rect 59138 521600 59143 521656
rect 59004 521598 59143 521600
rect 59004 521596 59010 521598
rect 59077 521595 59143 521598
rect 111241 521658 111307 521661
rect 136725 521658 136791 521661
rect 111241 521656 136791 521658
rect 111241 521600 111246 521656
rect 111302 521600 136730 521656
rect 136786 521600 136791 521656
rect 111241 521598 136791 521600
rect 111241 521595 111307 521598
rect 136725 521595 136791 521598
rect 179689 521658 179755 521661
rect 258441 521658 258507 521661
rect 179689 521656 258507 521658
rect 179689 521600 179694 521656
rect 179750 521600 258446 521656
rect 258502 521600 258507 521656
rect 179689 521598 258507 521600
rect 179689 521595 179755 521598
rect 258441 521595 258507 521598
rect 258717 521658 258783 521661
rect 265985 521658 266051 521661
rect 283189 521658 283255 521661
rect 258717 521656 266051 521658
rect 258717 521600 258722 521656
rect 258778 521600 265990 521656
rect 266046 521600 266051 521656
rect 258717 521598 266051 521600
rect 258717 521595 258783 521598
rect 265985 521595 266051 521598
rect 267690 521656 283255 521658
rect 267690 521600 283194 521656
rect 283250 521600 283255 521656
rect 267690 521598 283255 521600
rect 100293 521522 100359 521525
rect 134793 521522 134859 521525
rect 100293 521520 134859 521522
rect 100293 521464 100298 521520
rect 100354 521464 134798 521520
rect 134854 521464 134859 521520
rect 100293 521462 134859 521464
rect 100293 521459 100359 521462
rect 134793 521459 134859 521462
rect 134977 521522 135043 521525
rect 186221 521522 186287 521525
rect 134977 521520 186287 521522
rect 134977 521464 134982 521520
rect 135038 521464 186226 521520
rect 186282 521464 186287 521520
rect 134977 521462 186287 521464
rect 134977 521459 135043 521462
rect 186221 521459 186287 521462
rect 211061 521522 211127 521525
rect 240777 521522 240843 521525
rect 242525 521522 242591 521525
rect 211061 521520 240426 521522
rect 211061 521464 211066 521520
rect 211122 521464 240426 521520
rect 211061 521462 240426 521464
rect 211061 521459 211127 521462
rect 115105 521386 115171 521389
rect 217501 521386 217567 521389
rect 115105 521384 217567 521386
rect 115105 521328 115110 521384
rect 115166 521328 217506 521384
rect 217562 521328 217567 521384
rect 115105 521326 217567 521328
rect 115105 521323 115171 521326
rect 217501 521323 217567 521326
rect 218697 521386 218763 521389
rect 238753 521386 238819 521389
rect 218697 521384 238819 521386
rect 218697 521328 218702 521384
rect 218758 521328 238758 521384
rect 238814 521328 238819 521384
rect 218697 521326 238819 521328
rect 218697 521323 218763 521326
rect 238753 521323 238819 521326
rect 116117 521250 116183 521253
rect 219065 521250 219131 521253
rect 116117 521248 219131 521250
rect 116117 521192 116122 521248
rect 116178 521192 219070 521248
rect 219126 521192 219131 521248
rect 116117 521190 219131 521192
rect 116117 521187 116183 521190
rect 219065 521187 219131 521190
rect 231209 521250 231275 521253
rect 233141 521250 233207 521253
rect 231209 521248 233207 521250
rect 231209 521192 231214 521248
rect 231270 521192 233146 521248
rect 233202 521192 233207 521248
rect 231209 521190 233207 521192
rect 231209 521187 231275 521190
rect 233141 521187 233207 521190
rect 233877 521250 233943 521253
rect 234705 521250 234771 521253
rect 233877 521248 234771 521250
rect 233877 521192 233882 521248
rect 233938 521192 234710 521248
rect 234766 521192 234771 521248
rect 233877 521190 234771 521192
rect 240366 521250 240426 521462
rect 240777 521520 242591 521522
rect 240777 521464 240782 521520
rect 240838 521464 242530 521520
rect 242586 521464 242591 521520
rect 240777 521462 242591 521464
rect 240777 521459 240843 521462
rect 242525 521459 242591 521462
rect 246389 521522 246455 521525
rect 264421 521522 264487 521525
rect 246389 521520 264487 521522
rect 246389 521464 246394 521520
rect 246450 521464 264426 521520
rect 264482 521464 264487 521520
rect 246389 521462 264487 521464
rect 246389 521459 246455 521462
rect 264421 521459 264487 521462
rect 264605 521522 264671 521525
rect 267690 521522 267750 521598
rect 283189 521595 283255 521598
rect 294597 521658 294663 521661
rect 314469 521658 314535 521661
rect 294597 521656 314535 521658
rect 294597 521600 294602 521656
rect 294658 521600 314474 521656
rect 314530 521600 314535 521656
rect 294597 521598 314535 521600
rect 294597 521595 294663 521598
rect 314469 521595 314535 521598
rect 473261 521658 473327 521661
rect 497641 521658 497707 521661
rect 473261 521656 497707 521658
rect 473261 521600 473266 521656
rect 473322 521600 497646 521656
rect 497702 521600 497707 521656
rect 473261 521598 497707 521600
rect 473261 521595 473327 521598
rect 497641 521595 497707 521598
rect 264605 521520 267750 521522
rect 264605 521464 264610 521520
rect 264666 521464 267750 521520
rect 264605 521462 267750 521464
rect 278037 521522 278103 521525
rect 317597 521522 317663 521525
rect 278037 521520 317663 521522
rect 278037 521464 278042 521520
rect 278098 521464 317602 521520
rect 317658 521464 317663 521520
rect 278037 521462 317663 521464
rect 264605 521459 264671 521462
rect 278037 521459 278103 521462
rect 317597 521459 317663 521462
rect 472617 521522 472683 521525
rect 504357 521522 504423 521525
rect 472617 521520 504423 521522
rect 472617 521464 472622 521520
rect 472678 521464 504362 521520
rect 504418 521464 504423 521520
rect 472617 521462 504423 521464
rect 472617 521459 472683 521462
rect 504357 521459 504423 521462
rect 256141 521386 256207 521389
rect 319161 521386 319227 521389
rect 256141 521384 319227 521386
rect 256141 521328 256146 521384
rect 256202 521328 319166 521384
rect 319222 521328 319227 521384
rect 256141 521326 319227 521328
rect 256141 521323 256207 521326
rect 319161 521323 319227 521326
rect 372245 521386 372311 521389
rect 378593 521386 378659 521389
rect 372245 521384 378659 521386
rect 372245 521328 372250 521384
rect 372306 521328 378598 521384
rect 378654 521328 378659 521384
rect 372245 521326 378659 521328
rect 372245 521323 372311 521326
rect 378593 521323 378659 521326
rect 464521 521386 464587 521389
rect 495985 521386 496051 521389
rect 464521 521384 496051 521386
rect 464521 521328 464526 521384
rect 464582 521328 495990 521384
rect 496046 521328 496051 521384
rect 464521 521326 496051 521328
rect 464521 521323 464587 521326
rect 495985 521323 496051 521326
rect 245653 521250 245719 521253
rect 240366 521248 245719 521250
rect 240366 521192 245658 521248
rect 245714 521192 245719 521248
rect 240366 521190 245719 521192
rect 233877 521187 233943 521190
rect 234705 521187 234771 521190
rect 245653 521187 245719 521190
rect 255957 521250 256023 521253
rect 322289 521250 322355 521253
rect 255957 521248 322355 521250
rect 255957 521192 255962 521248
rect 256018 521192 322294 521248
rect 322350 521192 322355 521248
rect 255957 521190 322355 521192
rect 255957 521187 256023 521190
rect 322289 521187 322355 521190
rect 367001 521250 367067 521253
rect 391105 521250 391171 521253
rect 367001 521248 391171 521250
rect 367001 521192 367006 521248
rect 367062 521192 391110 521248
rect 391166 521192 391171 521248
rect 367001 521190 391171 521192
rect 367001 521187 367067 521190
rect 391105 521187 391171 521190
rect 461853 521250 461919 521253
rect 501413 521250 501479 521253
rect 461853 521248 501479 521250
rect 461853 521192 461858 521248
rect 461914 521192 501418 521248
rect 501474 521192 501479 521248
rect 461853 521190 501479 521192
rect 461853 521187 461919 521190
rect 501413 521187 501479 521190
rect 59302 521052 59308 521116
rect 59372 521114 59378 521116
rect 279366 521114 279372 521116
rect 59372 521054 279372 521114
rect 59372 521052 59378 521054
rect 279366 521052 279372 521054
rect 279436 521052 279442 521116
rect 287697 521114 287763 521117
rect 316033 521114 316099 521117
rect 287697 521112 316099 521114
rect 287697 521056 287702 521112
rect 287758 521056 316038 521112
rect 316094 521056 316099 521112
rect 287697 521054 316099 521056
rect 287697 521051 287763 521054
rect 316033 521051 316099 521054
rect 324313 521114 324379 521117
rect 384849 521114 384915 521117
rect 324313 521112 384915 521114
rect 324313 521056 324318 521112
rect 324374 521056 384854 521112
rect 384910 521056 384915 521112
rect 324313 521054 384915 521056
rect 324313 521051 324379 521054
rect 384849 521051 384915 521054
rect 461669 521114 461735 521117
rect 505553 521114 505619 521117
rect 461669 521112 505619 521114
rect 461669 521056 461674 521112
rect 461730 521056 505558 521112
rect 505614 521056 505619 521112
rect 461669 521054 505619 521056
rect 461669 521051 461735 521054
rect 505553 521051 505619 521054
rect 36854 520916 36860 520980
rect 36924 520978 36930 520980
rect 287830 520978 287836 520980
rect 36924 520918 287836 520978
rect 36924 520916 36930 520918
rect 287830 520916 287836 520918
rect 287900 520916 287906 520980
rect 299841 520978 299907 520981
rect 482461 520978 482527 520981
rect 299841 520976 482527 520978
rect 299841 520920 299846 520976
rect 299902 520920 482466 520976
rect 482522 520920 482527 520976
rect 299841 520918 482527 520920
rect 299841 520915 299907 520918
rect 482461 520915 482527 520918
rect 46013 520842 46079 520845
rect 99373 520842 99439 520845
rect 46013 520840 99439 520842
rect 46013 520784 46018 520840
rect 46074 520784 99378 520840
rect 99434 520784 99439 520840
rect 46013 520782 99439 520784
rect 46013 520779 46079 520782
rect 99373 520779 99439 520782
rect 114369 520842 114435 520845
rect 136633 520842 136699 520845
rect 114369 520840 136699 520842
rect 114369 520784 114374 520840
rect 114430 520784 136638 520840
rect 136694 520784 136699 520840
rect 114369 520782 136699 520784
rect 114369 520779 114435 520782
rect 136633 520779 136699 520782
rect 175917 520842 175983 520845
rect 215937 520842 216003 520845
rect 175917 520840 216003 520842
rect 175917 520784 175922 520840
rect 175978 520784 215942 520840
rect 215998 520784 216003 520840
rect 175917 520782 216003 520784
rect 175917 520779 175983 520782
rect 215937 520779 216003 520782
rect 238753 520842 238819 520845
rect 244089 520842 244155 520845
rect 238753 520840 244155 520842
rect 238753 520784 238758 520840
rect 238814 520784 244094 520840
rect 244150 520784 244155 520840
rect 238753 520782 244155 520784
rect 238753 520779 238819 520782
rect 244089 520779 244155 520782
rect 253197 520842 253263 520845
rect 269205 520842 269271 520845
rect 253197 520840 269271 520842
rect 253197 520784 253202 520840
rect 253258 520784 269210 520840
rect 269266 520784 269271 520840
rect 253197 520782 269271 520784
rect 253197 520779 253263 520782
rect 269205 520779 269271 520782
rect 275553 520842 275619 520845
rect 289445 520842 289511 520845
rect 275553 520840 289511 520842
rect 275553 520784 275558 520840
rect 275614 520784 289450 520840
rect 289506 520784 289511 520840
rect 275553 520782 289511 520784
rect 275553 520779 275619 520782
rect 289445 520779 289511 520782
rect 473353 520842 473419 520845
rect 482921 520842 482987 520845
rect 473353 520840 482987 520842
rect 473353 520784 473358 520840
rect 473414 520784 482926 520840
rect 482982 520784 482987 520840
rect 473353 520782 482987 520784
rect 473353 520779 473419 520782
rect 482921 520779 482987 520782
rect 50470 520644 50476 520708
rect 50540 520706 50546 520708
rect 110413 520706 110479 520709
rect 50540 520704 110479 520706
rect 50540 520648 110418 520704
rect 110474 520648 110479 520704
rect 50540 520646 110479 520648
rect 50540 520644 50546 520646
rect 110413 520643 110479 520646
rect 269757 520706 269823 520709
rect 278497 520706 278563 520709
rect 269757 520704 278563 520706
rect 269757 520648 269762 520704
rect 269818 520648 278502 520704
rect 278558 520648 278563 520704
rect 269757 520646 278563 520648
rect 269757 520643 269823 520646
rect 278497 520643 278563 520646
rect 47577 520570 47643 520573
rect 114461 520570 114527 520573
rect 47577 520568 114527 520570
rect 47577 520512 47582 520568
rect 47638 520512 114466 520568
rect 114522 520512 114527 520568
rect 47577 520510 114527 520512
rect 47577 520507 47643 520510
rect 114461 520507 114527 520510
rect 43897 520434 43963 520437
rect 117221 520434 117287 520437
rect 43897 520432 117287 520434
rect 43897 520376 43902 520432
rect 43958 520376 117226 520432
rect 117282 520376 117287 520432
rect 43897 520374 117287 520376
rect 43897 520371 43963 520374
rect 117221 520371 117287 520374
rect 42558 520236 42564 520300
rect 42628 520298 42634 520300
rect 115749 520298 115815 520301
rect 42628 520296 115815 520298
rect 42628 520240 115754 520296
rect 115810 520240 115815 520296
rect 42628 520238 115815 520240
rect 42628 520236 42634 520238
rect 115749 520235 115815 520238
rect 290917 520162 290983 520165
rect 492029 520162 492095 520165
rect 290917 520160 492095 520162
rect 290917 520104 290922 520160
rect 290978 520104 492034 520160
rect 492090 520104 492095 520160
rect 290917 520102 492095 520104
rect 290917 520099 290983 520102
rect 492029 520099 492095 520102
rect 495382 520100 495388 520164
rect 495452 520162 495458 520164
rect 495801 520162 495867 520165
rect 495452 520160 495867 520162
rect 495452 520104 495806 520160
rect 495862 520104 495867 520160
rect 495452 520102 495867 520104
rect 495452 520100 495458 520102
rect 495801 520099 495867 520102
rect 44909 520026 44975 520029
rect 57697 520026 57763 520029
rect 44909 520024 57763 520026
rect 44909 519968 44914 520024
rect 44970 519968 57702 520024
rect 57758 519968 57763 520024
rect 44909 519966 57763 519968
rect 44909 519963 44975 519966
rect 57697 519963 57763 519966
rect 283598 519964 283604 520028
rect 283668 520026 283674 520028
rect 490046 520026 490052 520028
rect 283668 519966 490052 520026
rect 283668 519964 283674 519966
rect 490046 519964 490052 519966
rect 490116 519964 490122 520028
rect 35566 519828 35572 519892
rect 35636 519890 35642 519892
rect 291929 519890 291995 519893
rect 35636 519888 291995 519890
rect 35636 519832 291934 519888
rect 291990 519832 291995 519888
rect 35636 519830 291995 519832
rect 35636 519828 35642 519830
rect 291929 519827 291995 519830
rect 45093 519754 45159 519757
rect 164141 519754 164207 519757
rect 45093 519752 164207 519754
rect 45093 519696 45098 519752
rect 45154 519696 164146 519752
rect 164202 519696 164207 519752
rect 45093 519694 164207 519696
rect 45093 519691 45159 519694
rect 164141 519691 164207 519694
rect 164325 519754 164391 519757
rect 375465 519754 375531 519757
rect 164325 519752 375531 519754
rect 164325 519696 164330 519752
rect 164386 519696 375470 519752
rect 375526 519696 375531 519752
rect 164325 519694 375531 519696
rect 164325 519691 164391 519694
rect 375465 519691 375531 519694
rect 462957 519754 463023 519757
rect 501505 519754 501571 519757
rect 462957 519752 501571 519754
rect 462957 519696 462962 519752
rect 463018 519696 501510 519752
rect 501566 519696 501571 519752
rect 462957 519694 501571 519696
rect 462957 519691 463023 519694
rect 501505 519691 501571 519694
rect 37406 519556 37412 519620
rect 37476 519618 37482 519620
rect 37476 519558 45570 519618
rect 37476 519556 37482 519558
rect 40677 519482 40743 519485
rect 44173 519482 44239 519485
rect 40677 519480 44239 519482
rect 40677 519424 40682 519480
rect 40738 519424 44178 519480
rect 44234 519424 44239 519480
rect 40677 519422 44239 519424
rect 45510 519482 45570 519558
rect 54886 519556 54892 519620
rect 54956 519618 54962 519620
rect 55121 519618 55187 519621
rect 54956 519616 55187 519618
rect 54956 519560 55126 519616
rect 55182 519560 55187 519616
rect 54956 519558 55187 519560
rect 54956 519556 54962 519558
rect 55121 519555 55187 519558
rect 57646 519556 57652 519620
rect 57716 519618 57722 519620
rect 255814 519618 255820 519620
rect 57716 519558 255820 519618
rect 57716 519556 57722 519558
rect 255814 519556 255820 519558
rect 255884 519556 255890 519620
rect 265750 519556 265756 519620
rect 265820 519618 265826 519620
rect 490230 519618 490236 519620
rect 265820 519558 490236 519618
rect 265820 519556 265826 519558
rect 490230 519556 490236 519558
rect 490300 519556 490306 519620
rect 285070 519482 285076 519484
rect 45510 519422 285076 519482
rect 40677 519419 40743 519422
rect 44173 519419 44239 519422
rect 285070 519420 285076 519422
rect 285140 519420 285146 519484
rect 290958 519420 290964 519484
rect 291028 519482 291034 519484
rect 291028 519422 495266 519482
rect 291028 519420 291034 519422
rect 42333 519346 42399 519349
rect 50153 519346 50219 519349
rect 42333 519344 50219 519346
rect 42333 519288 42338 519344
rect 42394 519288 50158 519344
rect 50214 519288 50219 519344
rect 42333 519286 50219 519288
rect 42333 519283 42399 519286
rect 50153 519283 50219 519286
rect 50286 519284 50292 519348
rect 50356 519346 50362 519348
rect 270401 519346 270467 519349
rect 50356 519344 270467 519346
rect 50356 519288 270406 519344
rect 270462 519288 270467 519344
rect 50356 519286 270467 519288
rect 50356 519284 50362 519286
rect 270401 519283 270467 519286
rect 291694 519284 291700 519348
rect 291764 519346 291770 519348
rect 491334 519346 491340 519348
rect 291764 519286 491340 519346
rect 291764 519284 291770 519286
rect 491334 519284 491340 519286
rect 491404 519284 491410 519348
rect 46422 519148 46428 519212
rect 46492 519210 46498 519212
rect 282913 519210 282979 519213
rect 46492 519208 282979 519210
rect 46492 519152 282918 519208
rect 282974 519152 282979 519208
rect 46492 519150 282979 519152
rect 46492 519148 46498 519150
rect 282913 519147 282979 519150
rect 284886 519148 284892 519212
rect 284956 519210 284962 519212
rect 494646 519210 494652 519212
rect 284956 519150 494652 519210
rect 284956 519148 284962 519150
rect 494646 519148 494652 519150
rect 494716 519148 494722 519212
rect 43478 519012 43484 519076
rect 43548 519074 43554 519076
rect 291009 519074 291075 519077
rect 43548 519072 291075 519074
rect 43548 519016 291014 519072
rect 291070 519016 291075 519072
rect 43548 519014 291075 519016
rect 43548 519012 43554 519014
rect 291009 519011 291075 519014
rect 483013 519074 483079 519077
rect 483422 519074 483428 519076
rect 483013 519072 483428 519074
rect 483013 519016 483018 519072
rect 483074 519016 483428 519072
rect 483013 519014 483428 519016
rect 483013 519011 483079 519014
rect 483422 519012 483428 519014
rect 483492 519012 483498 519076
rect 43345 518938 43411 518941
rect 45921 518938 45987 518941
rect 43345 518936 45987 518938
rect 43345 518880 43350 518936
rect 43406 518880 45926 518936
rect 45982 518880 45987 518936
rect 43345 518878 45987 518880
rect 43345 518875 43411 518878
rect 45921 518875 45987 518878
rect 54518 518876 54524 518940
rect 54588 518938 54594 518940
rect 55121 518938 55187 518941
rect 54588 518936 55187 518938
rect 54588 518880 55126 518936
rect 55182 518880 55187 518936
rect 54588 518878 55187 518880
rect 54588 518876 54594 518878
rect 55121 518875 55187 518878
rect 269614 518876 269620 518940
rect 269684 518938 269690 518940
rect 291837 518938 291903 518941
rect 495206 518940 495266 519422
rect 269684 518936 291903 518938
rect 269684 518880 291842 518936
rect 291898 518880 291903 518936
rect 269684 518878 291903 518880
rect 269684 518876 269690 518878
rect 291837 518875 291903 518878
rect 495198 518876 495204 518940
rect 495268 518876 495274 518940
rect 58525 518802 58591 518805
rect 269021 518802 269087 518805
rect 58525 518800 269087 518802
rect 58525 518744 58530 518800
rect 58586 518744 269026 518800
rect 269082 518744 269087 518800
rect 58525 518742 269087 518744
rect 58525 518739 58591 518742
rect 269021 518739 269087 518742
rect 476062 518740 476068 518804
rect 476132 518802 476138 518804
rect 477401 518802 477467 518805
rect 476132 518800 477467 518802
rect 476132 518744 477406 518800
rect 477462 518744 477467 518800
rect 476132 518742 477467 518744
rect 476132 518740 476138 518742
rect 477401 518739 477467 518742
rect 478086 518740 478092 518804
rect 478156 518802 478162 518804
rect 478781 518802 478847 518805
rect 478156 518800 478847 518802
rect 478156 518744 478786 518800
rect 478842 518744 478847 518800
rect 478156 518742 478847 518744
rect 478156 518740 478162 518742
rect 478781 518739 478847 518742
rect 58566 518604 58572 518668
rect 58636 518666 58642 518668
rect 271086 518666 271092 518668
rect 58636 518606 271092 518666
rect 58636 518604 58642 518606
rect 271086 518604 271092 518606
rect 271156 518604 271162 518668
rect 298870 518604 298876 518668
rect 298940 518666 298946 518668
rect 497222 518666 497228 518668
rect 298940 518606 497228 518666
rect 298940 518604 298946 518606
rect 497222 518604 497228 518606
rect 497292 518604 497298 518668
rect 268326 518468 268332 518532
rect 268396 518530 268402 518532
rect 503846 518530 503852 518532
rect 268396 518470 503852 518530
rect 268396 518468 268402 518470
rect 503846 518468 503852 518470
rect 503916 518468 503922 518532
rect 50654 518332 50660 518396
rect 50724 518394 50730 518396
rect 379830 518394 379836 518396
rect 50724 518334 379836 518394
rect 50724 518332 50730 518334
rect 379830 518332 379836 518334
rect 379900 518332 379906 518396
rect 461577 518394 461643 518397
rect 476113 518394 476179 518397
rect 461577 518392 476179 518394
rect 461577 518336 461582 518392
rect 461638 518336 476118 518392
rect 476174 518336 476179 518392
rect 461577 518334 476179 518336
rect 461577 518331 461643 518334
rect 476113 518331 476179 518334
rect 476798 518332 476804 518396
rect 476868 518394 476874 518396
rect 476868 518334 480270 518394
rect 476868 518332 476874 518334
rect 44582 518196 44588 518260
rect 44652 518258 44658 518260
rect 381302 518258 381308 518260
rect 44652 518198 381308 518258
rect 44652 518196 44658 518198
rect 381302 518196 381308 518198
rect 381372 518196 381378 518260
rect 476941 518258 477007 518261
rect 478505 518258 478571 518261
rect 476941 518256 478571 518258
rect 476941 518200 476946 518256
rect 477002 518200 478510 518256
rect 478566 518200 478571 518256
rect 476941 518198 478571 518200
rect 480210 518258 480270 518334
rect 491518 518258 491524 518260
rect 480210 518198 491524 518258
rect 476941 518195 477007 518198
rect 478505 518195 478571 518198
rect 491518 518196 491524 518198
rect 491588 518196 491594 518260
rect 44817 518122 44883 518125
rect 382273 518122 382339 518125
rect 44817 518120 382339 518122
rect 44817 518064 44822 518120
rect 44878 518064 382278 518120
rect 382334 518064 382339 518120
rect 44817 518062 382339 518064
rect 44817 518059 44883 518062
rect 382273 518059 382339 518062
rect 474406 518060 474412 518124
rect 474476 518122 474482 518124
rect 477309 518122 477375 518125
rect 474476 518120 477375 518122
rect 474476 518064 477314 518120
rect 477370 518064 477375 518120
rect 474476 518062 477375 518064
rect 474476 518060 474482 518062
rect 477309 518059 477375 518062
rect 478270 518060 478276 518124
rect 478340 518122 478346 518124
rect 478781 518122 478847 518125
rect 493358 518122 493364 518124
rect 478340 518120 478847 518122
rect 478340 518064 478786 518120
rect 478842 518064 478847 518120
rect 478340 518062 478847 518064
rect 478340 518060 478346 518062
rect 478781 518059 478847 518062
rect 479014 518062 493364 518122
rect 54518 517924 54524 517988
rect 54588 517986 54594 517988
rect 58985 517986 59051 517989
rect 61561 517986 61627 517989
rect 54588 517984 59051 517986
rect 54588 517928 58990 517984
rect 59046 517928 59051 517984
rect 54588 517926 59051 517928
rect 54588 517924 54594 517926
rect 58985 517923 59051 517926
rect 60598 517984 61627 517986
rect 60598 517928 61566 517984
rect 61622 517928 61627 517984
rect 60598 517926 61627 517928
rect 47485 517850 47551 517853
rect 58893 517850 58959 517853
rect 47485 517848 58959 517850
rect 47485 517792 47490 517848
rect 47546 517792 58898 517848
rect 58954 517792 58959 517848
rect 47485 517790 58959 517792
rect 47485 517787 47551 517790
rect 58893 517787 58959 517790
rect 60598 517684 60658 517926
rect 61561 517923 61627 517926
rect 476614 517924 476620 517988
rect 476684 517986 476690 517988
rect 479014 517986 479074 518062
rect 493358 518060 493364 518062
rect 493428 518060 493434 518124
rect 476684 517926 479074 517986
rect 476684 517924 476690 517926
rect 478505 517850 478571 517853
rect 478505 517848 479442 517850
rect 478505 517792 478510 517848
rect 478566 517792 479442 517848
rect 478505 517790 479442 517792
rect 478505 517787 478571 517790
rect 479382 517684 479442 517790
rect 58065 517578 58131 517581
rect 58750 517578 58756 517580
rect 58065 517576 58756 517578
rect 58065 517520 58070 517576
rect 58126 517520 58756 517576
rect 58065 517518 58756 517520
rect 58065 517515 58131 517518
rect 58750 517516 58756 517518
rect 58820 517516 58826 517580
rect 480069 517578 480135 517581
rect 483013 517578 483079 517581
rect 480069 517576 483079 517578
rect 480069 517520 480074 517576
rect 480130 517520 483018 517576
rect 483074 517520 483079 517576
rect 480069 517518 483079 517520
rect 480069 517515 480135 517518
rect 483013 517515 483079 517518
rect 481766 517306 481772 517308
rect 479934 517246 481772 517306
rect 57421 517170 57487 517173
rect 57421 517168 60076 517170
rect 57421 517112 57426 517168
rect 57482 517112 60076 517168
rect 479934 517140 479994 517246
rect 481766 517244 481772 517246
rect 481836 517244 481842 517308
rect 57421 517110 60076 517112
rect 57421 517107 57487 517110
rect 480161 516898 480227 516901
rect 481766 516898 481772 516900
rect 480161 516896 481772 516898
rect 480161 516840 480166 516896
rect 480222 516840 481772 516896
rect 480161 516838 481772 516840
rect 480161 516835 480227 516838
rect 481766 516836 481772 516838
rect 481836 516836 481842 516900
rect 482318 516762 482324 516764
rect 479934 516702 482324 516762
rect 57789 516626 57855 516629
rect 57789 516624 60076 516626
rect 57789 516568 57794 516624
rect 57850 516568 60076 516624
rect 479934 516596 479994 516702
rect 482318 516700 482324 516702
rect 482388 516700 482394 516764
rect 57789 516566 60076 516568
rect 57789 516563 57855 516566
rect 57329 516082 57395 516085
rect 57329 516080 60076 516082
rect 57329 516024 57334 516080
rect 57390 516024 60076 516080
rect 57329 516022 60076 516024
rect 57329 516019 57395 516022
rect 479934 515946 479994 516052
rect 482134 515946 482140 515948
rect 479934 515886 482140 515946
rect 482134 515884 482140 515886
rect 482204 515884 482210 515948
rect 482185 515810 482251 515813
rect 479934 515808 482251 515810
rect 479934 515752 482190 515808
rect 482246 515752 482251 515808
rect 479934 515750 482251 515752
rect 56869 515538 56935 515541
rect 56869 515536 60076 515538
rect 56869 515480 56874 515536
rect 56930 515480 60076 515536
rect 479934 515508 479994 515750
rect 482185 515747 482251 515750
rect 56869 515478 60076 515480
rect 56869 515475 56935 515478
rect 482001 515266 482067 515269
rect 479934 515264 482067 515266
rect 479934 515208 482006 515264
rect 482062 515208 482067 515264
rect 479934 515206 482067 515208
rect -960 514858 480 514948
rect 57830 514932 57836 514996
rect 57900 514994 57906 514996
rect 57900 514934 60076 514994
rect 479934 514964 479994 515206
rect 482001 515203 482067 515206
rect 57900 514932 57906 514934
rect 2998 514858 3004 514860
rect -960 514798 3004 514858
rect -960 514708 480 514798
rect 2998 514796 3004 514798
rect 3068 514796 3074 514860
rect 482185 514858 482251 514861
rect 482921 514858 482987 514861
rect 482185 514856 482987 514858
rect 482185 514800 482190 514856
rect 482246 514800 482926 514856
rect 482982 514800 482987 514856
rect 482185 514798 482987 514800
rect 482185 514795 482251 514798
rect 482921 514795 482987 514798
rect 481817 514722 481883 514725
rect 479934 514720 481883 514722
rect 479934 514664 481822 514720
rect 481878 514664 481883 514720
rect 479934 514662 481883 514664
rect 56961 514450 57027 514453
rect 56961 514448 60076 514450
rect 56961 514392 56966 514448
rect 57022 514392 60076 514448
rect 479934 514420 479994 514662
rect 481817 514659 481883 514662
rect 56961 514390 60076 514392
rect 56961 514387 57027 514390
rect 482369 514178 482435 514181
rect 479934 514176 482435 514178
rect 479934 514120 482374 514176
rect 482430 514120 482435 514176
rect 479934 514118 482435 514120
rect 57513 513906 57579 513909
rect 57513 513904 60076 513906
rect 57513 513848 57518 513904
rect 57574 513848 60076 513904
rect 479934 513876 479994 514118
rect 482369 514115 482435 514118
rect 57513 513846 60076 513848
rect 57513 513843 57579 513846
rect 57145 513362 57211 513365
rect 481725 513362 481791 513365
rect 57145 513360 60076 513362
rect 57145 513304 57150 513360
rect 57206 513304 60076 513360
rect 480210 513360 481791 513362
rect 57145 513302 60076 513304
rect 57145 513299 57211 513302
rect 479934 513226 479994 513332
rect 480210 513304 481730 513360
rect 481786 513304 481791 513360
rect 480210 513302 481791 513304
rect 480210 513226 480270 513302
rect 481725 513299 481791 513302
rect 479934 513166 480270 513226
rect 482553 513090 482619 513093
rect 479934 513088 482619 513090
rect 479934 513032 482558 513088
rect 482614 513032 482619 513088
rect 479934 513030 482619 513032
rect 57605 512818 57671 512821
rect 57605 512816 60076 512818
rect 57605 512760 57610 512816
rect 57666 512760 60076 512816
rect 479934 512788 479994 513030
rect 482553 513027 482619 513030
rect 57605 512758 60076 512760
rect 57605 512755 57671 512758
rect 481950 512410 481956 512412
rect 479934 512350 481956 512410
rect 57881 512274 57947 512277
rect 57881 512272 60076 512274
rect 57881 512216 57886 512272
rect 57942 512216 60076 512272
rect 479934 512244 479994 512350
rect 481950 512348 481956 512350
rect 482020 512348 482026 512412
rect 57881 512214 60076 512216
rect 57881 512211 57947 512214
rect 482369 512002 482435 512005
rect 483054 512002 483060 512004
rect 482369 512000 483060 512002
rect 482369 511944 482374 512000
rect 482430 511944 483060 512000
rect 482369 511942 483060 511944
rect 482369 511939 482435 511942
rect 483054 511940 483060 511942
rect 483124 511940 483130 512004
rect 503069 512002 503135 512005
rect 504081 512002 504147 512005
rect 503069 512000 504147 512002
rect 503069 511944 503074 512000
rect 503130 511944 504086 512000
rect 504142 511944 504147 512000
rect 503069 511942 504147 511944
rect 503069 511939 503135 511942
rect 504081 511939 504147 511942
rect 481633 511866 481699 511869
rect 479934 511864 481699 511866
rect 479934 511808 481638 511864
rect 481694 511808 481699 511864
rect 479934 511806 481699 511808
rect 58893 511730 58959 511733
rect 58893 511728 60076 511730
rect 58893 511672 58898 511728
rect 58954 511672 60076 511728
rect 479934 511700 479994 511806
rect 481633 511803 481699 511806
rect 58893 511670 60076 511672
rect 58893 511667 58959 511670
rect 481909 511594 481975 511597
rect 480210 511592 481975 511594
rect 480210 511536 481914 511592
rect 481970 511536 481975 511592
rect 480210 511534 481975 511536
rect 480210 511458 480270 511534
rect 481909 511531 481975 511534
rect 479934 511398 480270 511458
rect 36813 511186 36879 511189
rect 36813 511184 60076 511186
rect 36813 511128 36818 511184
rect 36874 511128 60076 511184
rect 479934 511156 479994 511398
rect 504081 511322 504147 511325
rect 583520 511322 584960 511412
rect 504081 511320 584960 511322
rect 504081 511264 504086 511320
rect 504142 511264 584960 511320
rect 504081 511262 584960 511264
rect 504081 511259 504147 511262
rect 583520 511172 584960 511262
rect 36813 511126 60076 511128
rect 36813 511123 36879 511126
rect 482277 510914 482343 510917
rect 479934 510912 482343 510914
rect 479934 510856 482282 510912
rect 482338 510856 482343 510912
rect 479934 510854 482343 510856
rect 44766 510580 44772 510644
rect 44836 510642 44842 510644
rect 44836 510582 60076 510642
rect 479934 510612 479994 510854
rect 482277 510851 482343 510854
rect 44836 510580 44842 510582
rect 43294 510444 43300 510508
rect 43364 510506 43370 510508
rect 43437 510506 43503 510509
rect 482277 510506 482343 510509
rect 483013 510506 483079 510509
rect 43364 510504 43503 510506
rect 43364 510448 43442 510504
rect 43498 510448 43503 510504
rect 43364 510446 43503 510448
rect 43364 510444 43370 510446
rect 43437 510443 43503 510446
rect 480210 510446 481466 510506
rect 480210 510370 480270 510446
rect 479934 510310 480270 510370
rect 481406 510370 481466 510446
rect 482277 510504 483079 510506
rect 482277 510448 482282 510504
rect 482338 510448 483018 510504
rect 483074 510448 483079 510504
rect 482277 510446 483079 510448
rect 482277 510443 482343 510446
rect 483013 510443 483079 510446
rect 482461 510370 482527 510373
rect 481406 510368 482527 510370
rect 481406 510312 482466 510368
rect 482522 510312 482527 510368
rect 481406 510310 482527 510312
rect 39798 510036 39804 510100
rect 39868 510098 39874 510100
rect 39868 510038 60076 510098
rect 479934 510068 479994 510310
rect 482461 510307 482527 510310
rect 39868 510036 39874 510038
rect 57789 509962 57855 509965
rect 59537 509962 59603 509965
rect 57789 509960 59603 509962
rect 57789 509904 57794 509960
rect 57850 509904 59542 509960
rect 59598 509904 59603 509960
rect 57789 509902 59603 509904
rect 57789 509899 57855 509902
rect 59537 509899 59603 509902
rect 44030 509492 44036 509556
rect 44100 509554 44106 509556
rect 491937 509554 492003 509557
rect 44100 509494 60076 509554
rect 480210 509552 492003 509554
rect 44100 509492 44106 509494
rect 479934 509418 479994 509524
rect 480210 509496 491942 509552
rect 491998 509496 492003 509552
rect 480210 509494 492003 509496
rect 480210 509418 480270 509494
rect 491937 509491 492003 509494
rect 479934 509358 480270 509418
rect 57881 509146 57947 509149
rect 58985 509146 59051 509149
rect 57881 509144 59051 509146
rect 57881 509088 57886 509144
rect 57942 509088 58990 509144
rect 59046 509088 59051 509144
rect 57881 509086 59051 509088
rect 57881 509083 57947 509086
rect 58985 509083 59051 509086
rect 42609 509010 42675 509013
rect 495566 509010 495572 509012
rect 42609 509008 60076 509010
rect 42609 508952 42614 509008
rect 42670 508952 60076 509008
rect 42609 508950 60076 508952
rect 42609 508947 42675 508950
rect 479934 508874 479994 508980
rect 480210 508950 495572 509010
rect 480210 508874 480270 508950
rect 495566 508948 495572 508950
rect 495636 508948 495642 509012
rect 479934 508814 480270 508874
rect 482645 508602 482711 508605
rect 490414 508602 490420 508604
rect 482645 508600 490420 508602
rect 482645 508544 482650 508600
rect 482706 508544 490420 508600
rect 482645 508542 490420 508544
rect 482645 508539 482711 508542
rect 490414 508540 490420 508542
rect 490484 508540 490490 508604
rect 41270 508404 41276 508468
rect 41340 508466 41346 508468
rect 496813 508466 496879 508469
rect 41340 508406 60076 508466
rect 480210 508464 496879 508466
rect 41340 508404 41346 508406
rect 479934 508330 479994 508436
rect 480210 508408 496818 508464
rect 496874 508408 496879 508464
rect 480210 508406 496879 508408
rect 480210 508330 480270 508406
rect 496813 508403 496879 508406
rect 479934 508270 480270 508330
rect 479934 507998 480270 508058
rect 50286 507860 50292 507924
rect 50356 507922 50362 507924
rect 50356 507862 60076 507922
rect 479934 507892 479994 507998
rect 480210 507922 480270 507998
rect 494462 507922 494468 507924
rect 480210 507862 494468 507922
rect 50356 507860 50362 507862
rect 494462 507860 494468 507862
rect 494532 507860 494538 507924
rect 47485 507378 47551 507381
rect 500166 507378 500172 507380
rect 47485 507376 60076 507378
rect 47485 507320 47490 507376
rect 47546 507320 60076 507376
rect 47485 507318 60076 507320
rect 47485 507315 47551 507318
rect 479934 507242 479994 507348
rect 480210 507318 500172 507378
rect 480210 507242 480270 507318
rect 500166 507316 500172 507318
rect 500236 507316 500242 507380
rect 479934 507182 480270 507242
rect 481633 507106 481699 507109
rect 479934 507104 481699 507106
rect 479934 507048 481638 507104
rect 481694 507048 481699 507104
rect 479934 507046 481699 507048
rect 54518 506772 54524 506836
rect 54588 506834 54594 506836
rect 54588 506774 60076 506834
rect 479934 506804 479994 507046
rect 481633 507043 481699 507046
rect 54588 506772 54594 506774
rect 57513 506426 57579 506429
rect 58525 506426 58591 506429
rect 57513 506424 58591 506426
rect 57513 506368 57518 506424
rect 57574 506368 58530 506424
rect 58586 506368 58591 506424
rect 57513 506366 58591 506368
rect 57513 506363 57579 506366
rect 58525 506363 58591 506366
rect 479934 506366 480270 506426
rect 46013 506290 46079 506293
rect 46013 506288 60076 506290
rect 46013 506232 46018 506288
rect 46074 506232 60076 506288
rect 479934 506260 479994 506366
rect 480210 506290 480270 506366
rect 482921 506290 482987 506293
rect 480210 506288 482987 506290
rect 46013 506230 60076 506232
rect 480210 506232 482926 506288
rect 482982 506232 482987 506288
rect 480210 506230 482987 506232
rect 46013 506227 46079 506230
rect 482921 506227 482987 506230
rect 482829 506154 482895 506157
rect 480210 506152 482895 506154
rect 480210 506096 482834 506152
rect 482890 506096 482895 506152
rect 480210 506094 482895 506096
rect 480210 506018 480270 506094
rect 482829 506091 482895 506094
rect 479934 505958 480270 506018
rect 43662 505684 43668 505748
rect 43732 505746 43738 505748
rect 43732 505686 60076 505746
rect 479934 505716 479994 505958
rect 43732 505684 43738 505686
rect 479934 505278 480270 505338
rect 43989 505204 44055 505205
rect 43989 505202 44036 505204
rect 43944 505200 44036 505202
rect 43944 505144 43994 505200
rect 43944 505142 44036 505144
rect 43989 505140 44036 505142
rect 44100 505140 44106 505204
rect 55622 505140 55628 505204
rect 55692 505202 55698 505204
rect 55692 505142 60076 505202
rect 479934 505172 479994 505278
rect 480210 505202 480270 505278
rect 501270 505202 501276 505204
rect 480210 505142 501276 505202
rect 55692 505140 55698 505142
rect 501270 505140 501276 505142
rect 501340 505140 501346 505204
rect 43989 505139 44055 505140
rect 50470 505004 50476 505068
rect 50540 505066 50546 505068
rect 57462 505066 57468 505068
rect 50540 505006 57468 505066
rect 50540 505004 50546 505006
rect 57462 505004 57468 505006
rect 57532 505004 57538 505068
rect 59486 504596 59492 504660
rect 59556 504658 59562 504660
rect 502926 504658 502932 504660
rect 59556 504598 60076 504658
rect 59556 504596 59562 504598
rect 57329 504522 57395 504525
rect 58985 504522 59051 504525
rect 57329 504520 59051 504522
rect 57329 504464 57334 504520
rect 57390 504464 58990 504520
rect 59046 504464 59051 504520
rect 57329 504462 59051 504464
rect 479934 504522 479994 504628
rect 480210 504598 502932 504658
rect 480210 504522 480270 504598
rect 502926 504596 502932 504598
rect 502996 504596 503002 504660
rect 479934 504462 480270 504522
rect 57329 504459 57395 504462
rect 58985 504459 59051 504462
rect 44633 504386 44699 504389
rect 57605 504386 57671 504389
rect 44633 504384 57671 504386
rect 44633 504328 44638 504384
rect 44694 504328 57610 504384
rect 57666 504328 57671 504384
rect 44633 504326 57671 504328
rect 44633 504323 44699 504326
rect 57605 504323 57671 504326
rect 35198 504052 35204 504116
rect 35268 504114 35274 504116
rect 498510 504114 498516 504116
rect 35268 504054 60076 504114
rect 35268 504052 35274 504054
rect 479934 503978 479994 504084
rect 480210 504054 498516 504114
rect 480210 503978 480270 504054
rect 498510 504052 498516 504054
rect 498580 504052 498586 504116
rect 479934 503918 480270 503978
rect 32857 503570 32923 503573
rect 32857 503568 60076 503570
rect 32857 503512 32862 503568
rect 32918 503512 60076 503568
rect 32857 503510 60076 503512
rect 32857 503507 32923 503510
rect 479934 503434 479994 503540
rect 485221 503434 485287 503437
rect 479934 503432 485287 503434
rect 479934 503376 485226 503432
rect 485282 503376 485287 503432
rect 479934 503374 485287 503376
rect 485221 503371 485287 503374
rect 57881 503026 57947 503029
rect 505461 503026 505527 503029
rect 57881 503024 60076 503026
rect 57881 502968 57886 503024
rect 57942 502968 60076 503024
rect 480210 503024 505527 503026
rect 57881 502966 60076 502968
rect 57881 502963 57947 502966
rect 479934 502890 479994 502996
rect 480210 502968 505466 503024
rect 505522 502968 505527 503024
rect 480210 502966 505527 502968
rect 480210 502890 480270 502966
rect 505461 502963 505527 502966
rect 479934 502830 480270 502890
rect 479934 502558 480270 502618
rect 58750 502420 58756 502484
rect 58820 502482 58826 502484
rect 59169 502482 59235 502485
rect 58820 502422 59048 502482
rect 58820 502420 58826 502422
rect 58988 502350 59048 502422
rect 59169 502480 60076 502482
rect 59169 502424 59174 502480
rect 59230 502424 60076 502480
rect 479934 502452 479994 502558
rect 480210 502482 480270 502558
rect 502742 502482 502748 502484
rect 59169 502422 60076 502424
rect 480210 502422 502748 502482
rect 59169 502419 59235 502422
rect 502742 502420 502748 502422
rect 502812 502420 502818 502484
rect 59118 502350 59124 502352
rect 58988 502290 59124 502350
rect 59118 502288 59124 502290
rect 59188 502288 59194 502352
rect 31385 501938 31451 501941
rect 506606 501938 506612 501940
rect 31385 501936 60076 501938
rect -960 501802 480 501892
rect 31385 501880 31390 501936
rect 31446 501880 60076 501936
rect 31385 501878 60076 501880
rect 31385 501875 31451 501878
rect 4654 501802 4660 501804
rect -960 501742 4660 501802
rect -960 501652 480 501742
rect 4654 501740 4660 501742
rect 4724 501740 4730 501804
rect 479934 501802 479994 501908
rect 480210 501878 506612 501938
rect 480210 501802 480270 501878
rect 506606 501876 506612 501878
rect 506676 501876 506682 501940
rect 479934 501742 480270 501802
rect 479885 501666 479951 501669
rect 479885 501664 479994 501666
rect 479885 501608 479890 501664
rect 479946 501608 479994 501664
rect 479885 501603 479994 501608
rect 36486 501332 36492 501396
rect 36556 501394 36562 501396
rect 36556 501334 60076 501394
rect 479934 501364 479994 501603
rect 36556 501332 36562 501334
rect 35382 500788 35388 500852
rect 35452 500850 35458 500852
rect 35452 500790 60076 500850
rect 35452 500788 35458 500790
rect 479934 500714 479994 500820
rect 480294 500714 480300 500716
rect 479934 500654 480300 500714
rect 480294 500652 480300 500654
rect 480364 500652 480370 500716
rect 482921 500578 482987 500581
rect 479934 500576 482987 500578
rect 479934 500520 482926 500576
rect 482982 500520 482987 500576
rect 479934 500518 482987 500520
rect 57513 500306 57579 500309
rect 57513 500304 60076 500306
rect 57513 500248 57518 500304
rect 57574 500248 60076 500304
rect 479934 500276 479994 500518
rect 482921 500515 482987 500518
rect 57513 500246 60076 500248
rect 57513 500243 57579 500246
rect 482829 500034 482895 500037
rect 479934 500032 482895 500034
rect 479934 499976 482834 500032
rect 482890 499976 482895 500032
rect 479934 499974 482895 499976
rect 42057 499762 42123 499765
rect 42057 499760 60076 499762
rect 42057 499704 42062 499760
rect 42118 499704 60076 499760
rect 479934 499732 479994 499974
rect 482829 499971 482895 499974
rect 42057 499702 60076 499704
rect 42057 499699 42123 499702
rect 57605 499354 57671 499357
rect 57605 499352 60106 499354
rect 57605 499296 57610 499352
rect 57666 499296 60106 499352
rect 57605 499294 60106 499296
rect 57605 499291 57671 499294
rect 47577 499218 47643 499221
rect 57513 499218 57579 499221
rect 47577 499216 57579 499218
rect 47577 499160 47582 499216
rect 47638 499160 57518 499216
rect 57574 499160 57579 499216
rect 60046 499188 60106 499294
rect 496077 499218 496143 499221
rect 480210 499216 496143 499218
rect 47577 499158 57579 499160
rect 47577 499155 47643 499158
rect 57513 499155 57579 499158
rect 46422 499020 46428 499084
rect 46492 499082 46498 499084
rect 57462 499082 57468 499084
rect 46492 499022 57468 499082
rect 46492 499020 46498 499022
rect 57462 499020 57468 499022
rect 57532 499020 57538 499084
rect 479934 499082 479994 499188
rect 480210 499160 496082 499216
rect 496138 499160 496143 499216
rect 480210 499158 496143 499160
rect 480210 499082 480270 499158
rect 496077 499155 496143 499158
rect 479934 499022 480270 499082
rect 40493 498946 40559 498949
rect 57605 498946 57671 498949
rect 40493 498944 57671 498946
rect 40493 498888 40498 498944
rect 40554 498888 57610 498944
rect 57666 498888 57671 498944
rect 40493 498886 57671 498888
rect 40493 498883 40559 498886
rect 57605 498883 57671 498886
rect 40585 498810 40651 498813
rect 57697 498810 57763 498813
rect 40585 498808 57763 498810
rect 40585 498752 40590 498808
rect 40646 498752 57702 498808
rect 57758 498752 57763 498808
rect 40585 498750 57763 498752
rect 40585 498747 40651 498750
rect 57697 498747 57763 498750
rect 57278 498612 57284 498676
rect 57348 498674 57354 498676
rect 501086 498674 501092 498676
rect 57348 498614 60076 498674
rect 57348 498612 57354 498614
rect 479934 498538 479994 498644
rect 480210 498614 501092 498674
rect 480210 498538 480270 498614
rect 501086 498612 501092 498614
rect 501156 498612 501162 498676
rect 479934 498478 480270 498538
rect 46238 498204 46244 498268
rect 46308 498266 46314 498268
rect 46473 498266 46539 498269
rect 46308 498264 46539 498266
rect 46308 498208 46478 498264
rect 46534 498208 46539 498264
rect 46308 498206 46539 498208
rect 46308 498204 46314 498206
rect 46473 498203 46539 498206
rect 34053 498130 34119 498133
rect 497222 498130 497228 498132
rect 34053 498128 60076 498130
rect 34053 498072 34058 498128
rect 34114 498072 60076 498128
rect 34053 498070 60076 498072
rect 34053 498067 34119 498070
rect 479934 497994 479994 498100
rect 480210 498070 497228 498130
rect 480210 497994 480270 498070
rect 497222 498068 497228 498070
rect 497292 498068 497298 498132
rect 479934 497934 480270 497994
rect 46105 497858 46171 497861
rect 57421 497858 57487 497861
rect 46105 497856 57487 497858
rect 46105 497800 46110 497856
rect 46166 497800 57426 497856
rect 57482 497800 57487 497856
rect 583520 497844 584960 498084
rect 46105 497798 57487 497800
rect 46105 497795 46171 497798
rect 57421 497795 57487 497798
rect 44817 497722 44883 497725
rect 57329 497722 57395 497725
rect 44817 497720 57395 497722
rect 44817 497664 44822 497720
rect 44878 497664 57334 497720
rect 57390 497664 57395 497720
rect 44817 497662 57395 497664
rect 44817 497659 44883 497662
rect 57329 497659 57395 497662
rect 57605 497586 57671 497589
rect 490230 497586 490236 497588
rect 57605 497584 60076 497586
rect 57605 497528 57610 497584
rect 57666 497528 60076 497584
rect 57605 497526 60076 497528
rect 57605 497523 57671 497526
rect 43529 497450 43595 497453
rect 57605 497450 57671 497453
rect 43529 497448 57671 497450
rect 43529 497392 43534 497448
rect 43590 497392 57610 497448
rect 57666 497392 57671 497448
rect 43529 497390 57671 497392
rect 479934 497450 479994 497556
rect 480210 497526 490236 497586
rect 480210 497450 480270 497526
rect 490230 497524 490236 497526
rect 490300 497524 490306 497588
rect 479934 497390 480270 497450
rect 43529 497387 43595 497390
rect 57605 497387 57671 497390
rect 57513 497042 57579 497045
rect 491518 497042 491524 497044
rect 57513 497040 60076 497042
rect 57513 496984 57518 497040
rect 57574 496984 60076 497040
rect 57513 496982 60076 496984
rect 57513 496979 57579 496982
rect 479934 496906 479994 497012
rect 480210 496982 491524 497042
rect 480210 496906 480270 496982
rect 491518 496980 491524 496982
rect 491588 496980 491594 497044
rect 479934 496846 480270 496906
rect 50654 496708 50660 496772
rect 50724 496770 50730 496772
rect 57278 496770 57284 496772
rect 50724 496710 57284 496770
rect 50724 496708 50730 496710
rect 57278 496708 57284 496710
rect 57348 496708 57354 496772
rect 38193 496498 38259 496501
rect 503846 496498 503852 496500
rect 38193 496496 60076 496498
rect 38193 496440 38198 496496
rect 38254 496440 60076 496496
rect 38193 496438 60076 496440
rect 38193 496435 38259 496438
rect 45001 496362 45067 496365
rect 57053 496362 57119 496365
rect 45001 496360 57119 496362
rect 45001 496304 45006 496360
rect 45062 496304 57058 496360
rect 57114 496304 57119 496360
rect 45001 496302 57119 496304
rect 479934 496362 479994 496468
rect 480210 496438 503852 496498
rect 480210 496362 480270 496438
rect 503846 496436 503852 496438
rect 503916 496436 503922 496500
rect 479934 496302 480270 496362
rect 45001 496299 45067 496302
rect 57053 496299 57119 496302
rect 57462 495892 57468 495956
rect 57532 495954 57538 495956
rect 493358 495954 493364 495956
rect 57532 495894 60076 495954
rect 57532 495892 57538 495894
rect 479934 495818 479994 495924
rect 480210 495894 493364 495954
rect 480210 495818 480270 495894
rect 493358 495892 493364 495894
rect 493428 495892 493434 495956
rect 479934 495758 480270 495818
rect 57145 495546 57211 495549
rect 58893 495546 58959 495549
rect 57145 495544 58959 495546
rect 57145 495488 57150 495544
rect 57206 495488 58898 495544
rect 58954 495488 58959 495544
rect 57145 495486 58959 495488
rect 57145 495483 57211 495486
rect 58893 495483 58959 495486
rect 482461 495546 482527 495549
rect 487654 495546 487660 495548
rect 482461 495544 487660 495546
rect 482461 495488 482466 495544
rect 482522 495488 487660 495544
rect 482461 495486 487660 495488
rect 482461 495483 482527 495486
rect 487654 495484 487660 495486
rect 487724 495484 487730 495548
rect 57697 495410 57763 495413
rect 494646 495410 494652 495412
rect 57697 495408 60076 495410
rect 57697 495352 57702 495408
rect 57758 495352 60076 495408
rect 57697 495350 60076 495352
rect 57697 495347 57763 495350
rect 479934 495274 479994 495380
rect 480210 495350 494652 495410
rect 480210 495274 480270 495350
rect 494646 495348 494652 495350
rect 494716 495348 494722 495412
rect 479934 495214 480270 495274
rect 33726 494804 33732 494868
rect 33796 494866 33802 494868
rect 506933 494866 506999 494869
rect 33796 494806 60076 494866
rect 480210 494864 506999 494866
rect 33796 494804 33802 494806
rect 479934 494730 479994 494836
rect 480210 494808 506938 494864
rect 506994 494808 506999 494864
rect 480210 494806 506999 494808
rect 480210 494730 480270 494806
rect 506933 494803 506999 494806
rect 479934 494670 480270 494730
rect 482829 494730 482895 494733
rect 485129 494730 485195 494733
rect 482829 494728 485195 494730
rect 482829 494672 482834 494728
rect 482890 494672 485134 494728
rect 485190 494672 485195 494728
rect 482829 494670 485195 494672
rect 482829 494667 482895 494670
rect 485129 494667 485195 494670
rect 57605 494322 57671 494325
rect 497038 494322 497044 494324
rect 57605 494320 60076 494322
rect 57605 494264 57610 494320
rect 57666 494264 60076 494320
rect 57605 494262 60076 494264
rect 57605 494259 57671 494262
rect 53281 494186 53347 494189
rect 57513 494186 57579 494189
rect 53281 494184 57579 494186
rect 53281 494128 53286 494184
rect 53342 494128 57518 494184
rect 57574 494128 57579 494184
rect 53281 494126 57579 494128
rect 479934 494186 479994 494292
rect 480210 494262 497044 494322
rect 480210 494186 480270 494262
rect 497038 494260 497044 494262
rect 497108 494260 497114 494324
rect 479934 494126 480270 494186
rect 53281 494123 53347 494126
rect 57513 494123 57579 494126
rect 32949 493778 33015 493781
rect 498694 493778 498700 493780
rect 32949 493776 60076 493778
rect 32949 493720 32954 493776
rect 33010 493720 60076 493776
rect 32949 493718 60076 493720
rect 32949 493715 33015 493718
rect 479934 493642 479994 493748
rect 480210 493718 498700 493778
rect 480210 493642 480270 493718
rect 498694 493716 498700 493718
rect 498764 493716 498770 493780
rect 479934 493582 480270 493642
rect 57421 493234 57487 493237
rect 500902 493234 500908 493236
rect 57421 493232 60076 493234
rect 57421 493176 57426 493232
rect 57482 493176 60076 493232
rect 57421 493174 60076 493176
rect 57421 493171 57487 493174
rect 479934 493098 479994 493204
rect 480210 493174 500908 493234
rect 480210 493098 480270 493174
rect 500902 493172 500908 493174
rect 500972 493172 500978 493236
rect 479934 493038 480270 493098
rect 57697 492962 57763 492965
rect 59629 492962 59695 492965
rect 57697 492960 59695 492962
rect 57697 492904 57702 492960
rect 57758 492904 59634 492960
rect 59690 492904 59695 492960
rect 57697 492902 59695 492904
rect 57697 492899 57763 492902
rect 59629 492899 59695 492902
rect 38101 492826 38167 492829
rect 38101 492824 60106 492826
rect 38101 492768 38106 492824
rect 38162 492768 60106 492824
rect 38101 492766 60106 492768
rect 38101 492763 38167 492766
rect 52126 492628 52132 492692
rect 52196 492690 52202 492692
rect 57145 492690 57211 492693
rect 52196 492688 57211 492690
rect 52196 492632 57150 492688
rect 57206 492632 57211 492688
rect 52196 492630 57211 492632
rect 52196 492628 52202 492630
rect 57145 492627 57211 492630
rect 58985 492690 59051 492693
rect 59445 492690 59511 492693
rect 58985 492688 59511 492690
rect 58985 492632 58990 492688
rect 59046 492632 59450 492688
rect 59506 492632 59511 492688
rect 60046 492660 60106 492766
rect 479934 492766 480270 492826
rect 479934 492660 479994 492766
rect 480210 492690 480270 492766
rect 490046 492690 490052 492692
rect 58985 492630 59511 492632
rect 480210 492630 490052 492690
rect 58985 492627 59051 492630
rect 59445 492627 59511 492630
rect 490046 492628 490052 492630
rect 490116 492628 490122 492692
rect 36670 492084 36676 492148
rect 36740 492146 36746 492148
rect 502558 492146 502564 492148
rect 36740 492086 60076 492146
rect 36740 492084 36746 492086
rect 479934 492010 479994 492116
rect 480210 492086 502564 492146
rect 480210 492010 480270 492086
rect 502558 492084 502564 492086
rect 502628 492084 502634 492148
rect 479934 491950 480270 492010
rect 482737 492010 482803 492013
rect 495709 492010 495775 492013
rect 482737 492008 495775 492010
rect 482737 491952 482742 492008
rect 482798 491952 495714 492008
rect 495770 491952 495775 492008
rect 482737 491950 495775 491952
rect 482737 491947 482803 491950
rect 495709 491947 495775 491950
rect 482921 491874 482987 491877
rect 497365 491874 497431 491877
rect 482921 491872 497431 491874
rect 482921 491816 482926 491872
rect 482982 491816 497370 491872
rect 497426 491816 497431 491872
rect 482921 491814 497431 491816
rect 482921 491811 482987 491814
rect 497365 491811 497431 491814
rect 57329 491602 57395 491605
rect 492029 491602 492095 491605
rect 57329 491600 60076 491602
rect 57329 491544 57334 491600
rect 57390 491544 60076 491600
rect 480210 491600 492095 491602
rect 57329 491542 60076 491544
rect 57329 491539 57395 491542
rect 479934 491466 479994 491572
rect 480210 491544 492034 491600
rect 492090 491544 492095 491600
rect 480210 491542 492095 491544
rect 480210 491466 480270 491542
rect 492029 491539 492095 491542
rect 479934 491406 480270 491466
rect 57513 491330 57579 491333
rect 57973 491330 58039 491333
rect 57513 491328 58039 491330
rect 57513 491272 57518 491328
rect 57574 491272 57978 491328
rect 58034 491272 58039 491328
rect 57513 491270 58039 491272
rect 57513 491267 57579 491270
rect 57973 491267 58039 491270
rect 42149 491194 42215 491197
rect 42558 491194 42564 491196
rect 42149 491192 42564 491194
rect 42149 491136 42154 491192
rect 42210 491136 42564 491192
rect 42149 491134 42564 491136
rect 42149 491131 42215 491134
rect 42558 491132 42564 491134
rect 42628 491132 42634 491196
rect 43478 490996 43484 491060
rect 43548 491058 43554 491060
rect 502374 491058 502380 491060
rect 43548 490998 60076 491058
rect 43548 490996 43554 490998
rect 479934 490922 479994 491028
rect 480210 490998 502380 491058
rect 480210 490922 480270 490998
rect 502374 490996 502380 490998
rect 502444 490996 502450 491060
rect 479934 490862 480270 490922
rect 42742 490452 42748 490516
rect 42812 490514 42818 490516
rect 494605 490514 494671 490517
rect 42812 490454 60076 490514
rect 480210 490512 494671 490514
rect 42812 490452 42818 490454
rect 479934 490378 479994 490484
rect 480210 490456 494610 490512
rect 494666 490456 494671 490512
rect 480210 490454 494671 490456
rect 480210 490378 480270 490454
rect 494605 490451 494671 490454
rect 479934 490318 480270 490378
rect 41086 490044 41092 490108
rect 41156 490106 41162 490108
rect 41156 490046 45570 490106
rect 41156 490044 41162 490046
rect 45510 489970 45570 490046
rect 495382 489970 495388 489972
rect 45510 489910 60076 489970
rect 479934 489930 479994 489940
rect 480118 489930 495388 489970
rect 479934 489910 495388 489930
rect 479934 489870 480178 489910
rect 495382 489908 495388 489910
rect 495452 489908 495458 489972
rect 57605 489834 57671 489837
rect 58065 489834 58131 489837
rect 57605 489832 58131 489834
rect 57605 489776 57610 489832
rect 57666 489776 58070 489832
rect 58126 489776 58131 489832
rect 57605 489774 58131 489776
rect 57605 489771 57671 489774
rect 58065 489771 58131 489774
rect 59169 489834 59235 489837
rect 59445 489834 59511 489837
rect 59169 489832 59511 489834
rect 59169 489776 59174 489832
rect 59230 489776 59450 489832
rect 59506 489776 59511 489832
rect 59169 489774 59511 489776
rect 59169 489771 59235 489774
rect 59445 489771 59511 489774
rect 479934 489502 480270 489562
rect 39246 489364 39252 489428
rect 39316 489426 39322 489428
rect 39316 489366 60076 489426
rect 479934 489396 479994 489502
rect 480210 489426 480270 489502
rect 498326 489426 498332 489428
rect 480210 489366 498332 489426
rect 39316 489364 39322 489366
rect 498326 489364 498332 489366
rect 498396 489364 498402 489428
rect 479934 488958 480270 489018
rect -960 488596 480 488836
rect 57278 488820 57284 488884
rect 57348 488882 57354 488884
rect 57348 488822 60076 488882
rect 479934 488852 479994 488958
rect 480210 488882 480270 488958
rect 491334 488882 491340 488884
rect 480210 488822 491340 488882
rect 57348 488820 57354 488822
rect 491334 488820 491340 488822
rect 491404 488820 491410 488884
rect 479934 488414 480270 488474
rect 44582 488276 44588 488340
rect 44652 488338 44658 488340
rect 44652 488278 60076 488338
rect 479934 488308 479994 488414
rect 480210 488338 480270 488414
rect 499798 488338 499804 488340
rect 480210 488278 499804 488338
rect 44652 488276 44658 488278
rect 499798 488276 499804 488278
rect 499868 488276 499874 488340
rect 479934 487870 480270 487930
rect 55438 487732 55444 487796
rect 55508 487794 55514 487796
rect 55508 487734 60076 487794
rect 479934 487764 479994 487870
rect 480210 487794 480270 487870
rect 514150 487794 514156 487796
rect 480210 487734 514156 487794
rect 55508 487732 55514 487734
rect 514150 487732 514156 487734
rect 514220 487732 514226 487796
rect 487470 487386 487476 487388
rect 479934 487326 487476 487386
rect 31569 487250 31635 487253
rect 31569 487248 60076 487250
rect 31569 487192 31574 487248
rect 31630 487192 60076 487248
rect 479934 487220 479994 487326
rect 487470 487324 487476 487326
rect 487540 487324 487546 487388
rect 31569 487190 60076 487192
rect 31569 487187 31635 487190
rect 479934 486782 480270 486842
rect 31477 486706 31543 486709
rect 31477 486704 60076 486706
rect 31477 486648 31482 486704
rect 31538 486648 60076 486704
rect 479934 486676 479994 486782
rect 480210 486706 480270 486782
rect 511390 486706 511396 486708
rect 31477 486646 60076 486648
rect 480210 486646 511396 486706
rect 31477 486643 31543 486646
rect 511390 486644 511396 486646
rect 511460 486644 511466 486708
rect 479934 486238 480270 486298
rect 33910 486100 33916 486164
rect 33980 486162 33986 486164
rect 33980 486102 60076 486162
rect 479934 486132 479994 486238
rect 480210 486162 480270 486238
rect 512126 486162 512132 486164
rect 480210 486102 512132 486162
rect 33980 486100 33986 486102
rect 512126 486100 512132 486102
rect 512196 486100 512202 486164
rect 511206 485828 511212 485892
rect 511276 485890 511282 485892
rect 511901 485890 511967 485893
rect 511276 485888 511967 485890
rect 511276 485832 511906 485888
rect 511962 485832 511967 485888
rect 511276 485830 511967 485832
rect 511276 485828 511282 485830
rect 511901 485827 511967 485830
rect 479934 485694 480270 485754
rect 39430 485556 39436 485620
rect 39500 485618 39506 485620
rect 39500 485558 60076 485618
rect 479934 485588 479994 485694
rect 480210 485618 480270 485694
rect 510654 485618 510660 485620
rect 480210 485558 510660 485618
rect 39500 485556 39506 485558
rect 510654 485556 510660 485558
rect 510724 485556 510730 485620
rect 479934 485150 480270 485210
rect 30966 485012 30972 485076
rect 31036 485074 31042 485076
rect 31036 485014 60076 485074
rect 479934 485044 479994 485150
rect 480210 485074 480270 485150
rect 507894 485074 507900 485076
rect 480210 485014 507900 485074
rect 31036 485012 31042 485014
rect 507894 485012 507900 485014
rect 507964 485012 507970 485076
rect 479934 484606 480270 484666
rect 29862 484468 29868 484532
rect 29932 484530 29938 484532
rect 29932 484470 60076 484530
rect 479934 484500 479994 484606
rect 480210 484530 480270 484606
rect 580206 484604 580212 484668
rect 580276 484666 580282 484668
rect 583520 484666 584960 484756
rect 580276 484606 584960 484666
rect 580276 484604 580282 484606
rect 503662 484530 503668 484532
rect 480210 484470 503668 484530
rect 29932 484468 29938 484470
rect 503662 484468 503668 484470
rect 503732 484468 503738 484532
rect 583520 484516 584960 484606
rect 479934 484062 480270 484122
rect 30046 483924 30052 483988
rect 30116 483986 30122 483988
rect 30116 483926 60076 483986
rect 479934 483956 479994 484062
rect 480210 483986 480270 484062
rect 499982 483986 499988 483988
rect 480210 483926 499988 483986
rect 30116 483924 30122 483926
rect 499982 483924 499988 483926
rect 500052 483924 500058 483988
rect 479934 483518 480270 483578
rect 32438 483380 32444 483444
rect 32508 483442 32514 483444
rect 32508 483382 60076 483442
rect 479934 483412 479994 483518
rect 480210 483442 480270 483518
rect 505134 483442 505140 483444
rect 480210 483382 505140 483442
rect 32508 483380 32514 483382
rect 505134 483380 505140 483382
rect 505204 483380 505210 483444
rect 42374 482972 42380 483036
rect 42444 483034 42450 483036
rect 42444 482974 42626 483034
rect 42444 482972 42450 482974
rect 42241 482898 42307 482901
rect 42374 482898 42380 482900
rect 42241 482896 42380 482898
rect 42241 482840 42246 482896
rect 42302 482840 42380 482896
rect 42241 482838 42380 482840
rect 42241 482835 42307 482838
rect 42374 482836 42380 482838
rect 42444 482836 42450 482900
rect 42566 482898 42626 482974
rect 493174 482898 493180 482900
rect 42566 482838 60076 482898
rect 479934 482762 479994 482868
rect 480210 482838 493180 482898
rect 480210 482762 480270 482838
rect 493174 482836 493180 482838
rect 493244 482836 493250 482900
rect 479934 482702 480270 482762
rect 479934 482430 480270 482490
rect 36905 482354 36971 482357
rect 36905 482352 60076 482354
rect 36905 482296 36910 482352
rect 36966 482296 60076 482352
rect 479934 482324 479994 482430
rect 480210 482354 480270 482430
rect 501505 482354 501571 482357
rect 480210 482352 501571 482354
rect 36905 482294 60076 482296
rect 480210 482296 501510 482352
rect 501566 482296 501571 482352
rect 480210 482294 501571 482296
rect 36905 482291 36971 482294
rect 501505 482291 501571 482294
rect 479934 481886 480270 481946
rect 50797 481810 50863 481813
rect 50797 481808 60076 481810
rect 50797 481752 50802 481808
rect 50858 481752 60076 481808
rect 479934 481780 479994 481886
rect 480210 481810 480270 481886
rect 504357 481810 504423 481813
rect 480210 481808 504423 481810
rect 50797 481750 60076 481752
rect 480210 481752 504362 481808
rect 504418 481752 504423 481808
rect 480210 481750 504423 481752
rect 50797 481747 50863 481750
rect 504357 481747 504423 481750
rect 479934 481342 480270 481402
rect 35709 481266 35775 481269
rect 35709 481264 60076 481266
rect 35709 481208 35714 481264
rect 35770 481208 60076 481264
rect 479934 481236 479994 481342
rect 480210 481266 480270 481342
rect 505553 481266 505619 481269
rect 480210 481264 505619 481266
rect 35709 481206 60076 481208
rect 480210 481208 505558 481264
rect 505614 481208 505619 481264
rect 480210 481206 505619 481208
rect 35709 481203 35775 481206
rect 505553 481203 505619 481206
rect 479934 480798 480270 480858
rect 36997 480722 37063 480725
rect 36997 480720 60076 480722
rect 36997 480664 37002 480720
rect 37058 480664 60076 480720
rect 479934 480692 479994 480798
rect 480210 480722 480270 480798
rect 501413 480722 501479 480725
rect 480210 480720 501479 480722
rect 36997 480662 60076 480664
rect 480210 480664 501418 480720
rect 501474 480664 501479 480720
rect 480210 480662 501479 480664
rect 36997 480659 37063 480662
rect 501413 480659 501479 480662
rect 57145 480178 57211 480181
rect 57145 480176 60076 480178
rect 57145 480120 57150 480176
rect 57206 480120 60076 480176
rect 57145 480118 60076 480120
rect 57145 480115 57211 480118
rect 479934 480042 479994 480148
rect 485957 480042 486023 480045
rect 479934 480040 486023 480042
rect 479934 479984 485962 480040
rect 486018 479984 486023 480040
rect 479934 479982 486023 479984
rect 485957 479979 486023 479982
rect 479977 479906 480043 479909
rect 479934 479904 480043 479906
rect 479934 479848 479982 479904
rect 480038 479848 480043 479904
rect 479934 479843 480043 479848
rect 35617 479634 35683 479637
rect 35617 479632 60076 479634
rect 35617 479576 35622 479632
rect 35678 479576 60076 479632
rect 479934 479604 479994 479843
rect 35617 479574 60076 479576
rect 35617 479571 35683 479574
rect 482093 479362 482159 479365
rect 479934 479360 482159 479362
rect 479934 479304 482098 479360
rect 482154 479304 482159 479360
rect 479934 479302 482159 479304
rect 40677 479090 40743 479093
rect 40677 479088 60076 479090
rect 40677 479032 40682 479088
rect 40738 479032 60076 479088
rect 479934 479060 479994 479302
rect 482093 479299 482159 479302
rect 40677 479030 60076 479032
rect 40677 479027 40743 479030
rect 39389 478546 39455 478549
rect 495985 478546 496051 478549
rect 39389 478544 60076 478546
rect 39389 478488 39394 478544
rect 39450 478488 60076 478544
rect 480210 478544 496051 478546
rect 39389 478486 60076 478488
rect 39389 478483 39455 478486
rect 479934 478410 479994 478516
rect 480210 478488 495990 478544
rect 496046 478488 496051 478544
rect 480210 478486 496051 478488
rect 480210 478410 480270 478486
rect 495985 478483 496051 478486
rect 479934 478350 480270 478410
rect 482093 478274 482159 478277
rect 479934 478272 482159 478274
rect 479934 478216 482098 478272
rect 482154 478216 482159 478272
rect 479934 478214 482159 478216
rect 53465 478002 53531 478005
rect 53465 478000 60076 478002
rect 53465 477944 53470 478000
rect 53526 477944 60076 478000
rect 479934 477972 479994 478214
rect 482093 478211 482159 478214
rect 53465 477942 60076 477944
rect 53465 477939 53531 477942
rect 38285 477458 38351 477461
rect 498745 477458 498811 477461
rect 38285 477456 60076 477458
rect 38285 477400 38290 477456
rect 38346 477400 60076 477456
rect 480210 477456 498811 477458
rect 38285 477398 60076 477400
rect 38285 477395 38351 477398
rect 479934 477322 479994 477428
rect 480210 477400 498750 477456
rect 498806 477400 498811 477456
rect 480210 477398 498811 477400
rect 480210 477322 480270 477398
rect 498745 477395 498811 477398
rect 479934 477262 480270 477322
rect 54702 476852 54708 476916
rect 54772 476914 54778 476916
rect 54772 476854 60076 476914
rect 54772 476852 54778 476854
rect 479934 476778 479994 476884
rect 488993 476778 489059 476781
rect 479934 476776 489059 476778
rect 479934 476720 488998 476776
rect 489054 476720 489059 476776
rect 479934 476718 489059 476720
rect 488993 476715 489059 476718
rect 43345 476370 43411 476373
rect 501321 476370 501387 476373
rect 43345 476368 60076 476370
rect 43345 476312 43350 476368
rect 43406 476312 60076 476368
rect 480210 476368 501387 476370
rect 43345 476310 60076 476312
rect 43345 476307 43411 476310
rect 479934 476234 479994 476340
rect 480210 476312 501326 476368
rect 501382 476312 501387 476368
rect 480210 476310 501387 476312
rect 480210 476234 480270 476310
rect 501321 476307 501387 476310
rect 479934 476174 480270 476234
rect 479517 476098 479583 476101
rect 479517 476096 479626 476098
rect 479517 476040 479522 476096
rect 479578 476040 479626 476096
rect 479517 476035 479626 476040
rect 38561 475826 38627 475829
rect 38561 475824 60076 475826
rect -960 475690 480 475780
rect 38561 475768 38566 475824
rect 38622 475768 60076 475824
rect 479566 475796 479626 476035
rect 38561 475766 60076 475768
rect 38561 475763 38627 475766
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 57513 475282 57579 475285
rect 57513 475280 60076 475282
rect 57513 475224 57518 475280
rect 57574 475224 60076 475280
rect 57513 475222 60076 475224
rect 57513 475219 57579 475222
rect 479934 475146 479994 475252
rect 487521 475146 487587 475149
rect 479934 475144 487587 475146
rect 479934 475088 487526 475144
rect 487582 475088 487587 475144
rect 479934 475086 487587 475088
rect 487521 475083 487587 475086
rect 38377 474738 38443 474741
rect 482093 474738 482159 474741
rect 38377 474736 60076 474738
rect 38377 474680 38382 474736
rect 38438 474680 60076 474736
rect 480210 474736 482159 474738
rect 38377 474678 60076 474680
rect 38377 474675 38443 474678
rect 479934 474602 479994 474708
rect 480210 474680 482098 474736
rect 482154 474680 482159 474736
rect 480210 474678 482159 474680
rect 480210 474602 480270 474678
rect 482093 474675 482159 474678
rect 479934 474542 480270 474602
rect 480345 474466 480411 474469
rect 479934 474464 480411 474466
rect 479934 474408 480350 474464
rect 480406 474408 480411 474464
rect 479934 474406 480411 474408
rect 53649 474194 53715 474197
rect 53649 474192 60076 474194
rect 53649 474136 53654 474192
rect 53710 474136 60076 474192
rect 479934 474164 479994 474406
rect 480345 474403 480411 474406
rect 53649 474134 60076 474136
rect 53649 474131 53715 474134
rect 480437 474058 480503 474061
rect 480210 474056 480503 474058
rect 480210 474000 480442 474056
rect 480498 474000 480503 474056
rect 480210 473998 480503 474000
rect 480210 473922 480270 473998
rect 480437 473995 480503 473998
rect 479934 473862 480270 473922
rect 52085 473650 52151 473653
rect 52085 473648 60076 473650
rect 52085 473592 52090 473648
rect 52146 473592 60076 473648
rect 479934 473620 479994 473862
rect 52085 473590 60076 473592
rect 52085 473587 52151 473590
rect 53741 473106 53807 473109
rect 53741 473104 60076 473106
rect 53741 473048 53746 473104
rect 53802 473048 60076 473104
rect 53741 473046 60076 473048
rect 53741 473043 53807 473046
rect 479934 472970 479994 473076
rect 488901 472970 488967 472973
rect 479934 472968 488967 472970
rect 479934 472912 488906 472968
rect 488962 472912 488967 472968
rect 479934 472910 488967 472912
rect 488901 472907 488967 472910
rect 52177 472562 52243 472565
rect 502701 472562 502767 472565
rect 52177 472560 60076 472562
rect 52177 472504 52182 472560
rect 52238 472504 60076 472560
rect 480210 472560 502767 472562
rect 52177 472502 60076 472504
rect 52177 472499 52243 472502
rect 479934 472426 479994 472532
rect 480210 472504 502706 472560
rect 502762 472504 502767 472560
rect 480210 472502 502767 472504
rect 480210 472426 480270 472502
rect 502701 472499 502767 472502
rect 479934 472366 480270 472426
rect 482093 472290 482159 472293
rect 479934 472288 482159 472290
rect 479934 472232 482098 472288
rect 482154 472232 482159 472288
rect 479934 472230 482159 472232
rect 39849 472018 39915 472021
rect 39849 472016 60076 472018
rect 39849 471960 39854 472016
rect 39910 471960 60076 472016
rect 479934 471988 479994 472230
rect 482093 472227 482159 472230
rect 39849 471958 60076 471960
rect 39849 471955 39915 471958
rect 482001 471746 482067 471749
rect 479934 471744 482067 471746
rect 479934 471688 482006 471744
rect 482062 471688 482067 471744
rect 479934 471686 482067 471688
rect 51993 471474 52059 471477
rect 51993 471472 60076 471474
rect 51993 471416 51998 471472
rect 52054 471416 60076 471472
rect 479934 471444 479994 471686
rect 482001 471683 482067 471686
rect 51993 471414 60076 471416
rect 51993 471411 52059 471414
rect 544326 471412 544332 471476
rect 544396 471474 544402 471476
rect 583520 471474 584960 471564
rect 544396 471414 584960 471474
rect 544396 471412 544402 471414
rect 583520 471324 584960 471414
rect 482093 471202 482159 471205
rect 479934 471200 482159 471202
rect 479934 471144 482098 471200
rect 482154 471144 482159 471200
rect 479934 471142 482159 471144
rect 53557 470930 53623 470933
rect 53557 470928 60076 470930
rect 53557 470872 53562 470928
rect 53618 470872 60076 470928
rect 479934 470900 479994 471142
rect 482093 471139 482159 471142
rect 53557 470870 60076 470872
rect 53557 470867 53623 470870
rect 42333 470386 42399 470389
rect 482001 470386 482067 470389
rect 42333 470384 60076 470386
rect 42333 470328 42338 470384
rect 42394 470328 60076 470384
rect 480210 470384 482067 470386
rect 42333 470326 60076 470328
rect 42333 470323 42399 470326
rect 479934 470250 479994 470356
rect 480210 470328 482006 470384
rect 482062 470328 482067 470384
rect 480210 470326 482067 470328
rect 480210 470250 480270 470326
rect 482001 470323 482067 470326
rect 479934 470190 480270 470250
rect 44909 469842 44975 469845
rect 44909 469840 60076 469842
rect 44909 469784 44914 469840
rect 44970 469784 60076 469840
rect 44909 469782 60076 469784
rect 44909 469779 44975 469782
rect 479934 469706 479994 469812
rect 488717 469706 488783 469709
rect 479934 469704 488783 469706
rect 479934 469648 488722 469704
rect 488778 469648 488783 469704
rect 479934 469646 488783 469648
rect 488717 469643 488783 469646
rect 482093 469570 482159 469573
rect 479934 469568 482159 469570
rect 479934 469512 482098 469568
rect 482154 469512 482159 469568
rect 479934 469510 482159 469512
rect 54293 469298 54359 469301
rect 54293 469296 60076 469298
rect 54293 469240 54298 469296
rect 54354 469240 60076 469296
rect 479934 469268 479994 469510
rect 482093 469507 482159 469510
rect 54293 469238 60076 469240
rect 54293 469235 54359 469238
rect 482093 469026 482159 469029
rect 479934 469024 482159 469026
rect 479934 468968 482098 469024
rect 482154 468968 482159 469024
rect 479934 468966 482159 468968
rect 57421 468754 57487 468757
rect 57421 468752 60076 468754
rect 57421 468696 57426 468752
rect 57482 468696 60076 468752
rect 479934 468724 479994 468966
rect 482093 468963 482159 468966
rect 57421 468694 60076 468696
rect 57421 468691 57487 468694
rect 482001 468618 482067 468621
rect 480210 468616 482067 468618
rect 480210 468560 482006 468616
rect 482062 468560 482067 468616
rect 480210 468558 482067 468560
rect 480210 468482 480270 468558
rect 482001 468555 482067 468558
rect 479934 468422 480270 468482
rect 55029 468210 55095 468213
rect 55029 468208 60076 468210
rect 55029 468152 55034 468208
rect 55090 468152 60076 468208
rect 479934 468180 479994 468422
rect 55029 468150 60076 468152
rect 55029 468147 55095 468150
rect 482001 467802 482067 467805
rect 479934 467800 482067 467802
rect 479934 467744 482006 467800
rect 482062 467744 482067 467800
rect 479934 467742 482067 467744
rect 55765 467666 55831 467669
rect 55765 467664 60076 467666
rect 55765 467608 55770 467664
rect 55826 467608 60076 467664
rect 479934 467636 479994 467742
rect 482001 467739 482067 467742
rect 55765 467606 60076 467608
rect 55765 467603 55831 467606
rect 479333 467394 479399 467397
rect 479333 467392 479442 467394
rect 479333 467336 479338 467392
rect 479394 467336 479442 467392
rect 479333 467331 479442 467336
rect 41321 467122 41387 467125
rect 41321 467120 60076 467122
rect 41321 467064 41326 467120
rect 41382 467064 60076 467120
rect 479382 467092 479442 467331
rect 41321 467062 60076 467064
rect 41321 467059 41387 467062
rect 482093 466850 482159 466853
rect 479934 466848 482159 466850
rect 479934 466792 482098 466848
rect 482154 466792 482159 466848
rect 479934 466790 482159 466792
rect 59077 466578 59143 466581
rect 59077 466576 60076 466578
rect 59077 466520 59082 466576
rect 59138 466520 60076 466576
rect 479934 466548 479994 466790
rect 482093 466787 482159 466790
rect 59077 466518 60076 466520
rect 59077 466515 59143 466518
rect 43621 466034 43687 466037
rect 43621 466032 60076 466034
rect 43621 465976 43626 466032
rect 43682 465976 60076 466032
rect 43621 465974 60076 465976
rect 43621 465971 43687 465974
rect 479934 465898 479994 466004
rect 486182 465898 486188 465900
rect 479934 465838 486188 465898
rect 486182 465836 486188 465838
rect 486252 465836 486258 465900
rect 480253 465762 480319 465765
rect 479934 465760 480319 465762
rect 479934 465704 480258 465760
rect 480314 465704 480319 465760
rect 479934 465702 480319 465704
rect 42701 465490 42767 465493
rect 42701 465488 60076 465490
rect 42701 465432 42706 465488
rect 42762 465432 60076 465488
rect 479934 465460 479994 465702
rect 480253 465699 480319 465702
rect 42701 465430 60076 465432
rect 42701 465427 42767 465430
rect 36629 464946 36695 464949
rect 482093 464946 482159 464949
rect 36629 464944 60076 464946
rect 36629 464888 36634 464944
rect 36690 464888 60076 464944
rect 480210 464944 482159 464946
rect 36629 464886 60076 464888
rect 36629 464883 36695 464886
rect 479934 464810 479994 464916
rect 480210 464888 482098 464944
rect 482154 464888 482159 464944
rect 480210 464886 482159 464888
rect 480210 464810 480270 464886
rect 482093 464883 482159 464886
rect 479934 464750 480270 464810
rect 482001 464674 482067 464677
rect 479934 464672 482067 464674
rect 479934 464616 482006 464672
rect 482062 464616 482067 464672
rect 479934 464614 482067 464616
rect 35433 464402 35499 464405
rect 35433 464400 60076 464402
rect 35433 464344 35438 464400
rect 35494 464344 60076 464400
rect 479934 464372 479994 464614
rect 482001 464611 482067 464614
rect 35433 464342 60076 464344
rect 35433 464339 35499 464342
rect 482093 464130 482159 464133
rect 479934 464128 482159 464130
rect 479934 464072 482098 464128
rect 482154 464072 482159 464128
rect 479934 464070 482159 464072
rect 57605 463858 57671 463861
rect 57605 463856 60076 463858
rect 57605 463800 57610 463856
rect 57666 463800 60076 463856
rect 479934 463828 479994 464070
rect 482093 464067 482159 464070
rect 57605 463798 60076 463800
rect 57605 463795 57671 463798
rect 482093 463450 482159 463453
rect 479934 463448 482159 463450
rect 479934 463392 482098 463448
rect 482154 463392 482159 463448
rect 479934 463390 482159 463392
rect 37089 463314 37155 463317
rect 37089 463312 60076 463314
rect 37089 463256 37094 463312
rect 37150 463256 60076 463312
rect 479934 463284 479994 463390
rect 482093 463387 482159 463390
rect 37089 463254 60076 463256
rect 37089 463251 37155 463254
rect 482093 463042 482159 463045
rect 479934 463040 482159 463042
rect 479934 462984 482098 463040
rect 482154 462984 482159 463040
rect 479934 462982 482159 462984
rect 50981 462770 51047 462773
rect 50981 462768 60076 462770
rect -960 462634 480 462724
rect 50981 462712 50986 462768
rect 51042 462712 60076 462768
rect 479934 462740 479994 462982
rect 482093 462979 482159 462982
rect 50981 462710 60076 462712
rect 50981 462707 51047 462710
rect 3366 462634 3372 462636
rect -960 462574 3372 462634
rect -960 462484 480 462574
rect 3366 462572 3372 462574
rect 3436 462572 3442 462636
rect 35341 462226 35407 462229
rect 35341 462224 60076 462226
rect 35341 462168 35346 462224
rect 35402 462168 60076 462224
rect 35341 462166 60076 462168
rect 35341 462163 35407 462166
rect 479934 462090 479994 462196
rect 482093 462090 482159 462093
rect 479934 462088 482159 462090
rect 479934 462032 482098 462088
rect 482154 462032 482159 462088
rect 479934 462030 482159 462032
rect 482093 462027 482159 462030
rect 482001 461954 482067 461957
rect 479934 461952 482067 461954
rect 479934 461896 482006 461952
rect 482062 461896 482067 461952
rect 479934 461894 482067 461896
rect 50889 461682 50955 461685
rect 50889 461680 60076 461682
rect 50889 461624 50894 461680
rect 50950 461624 60076 461680
rect 479934 461652 479994 461894
rect 482001 461891 482067 461894
rect 50889 461622 60076 461624
rect 50889 461619 50955 461622
rect 481909 461410 481975 461413
rect 479934 461408 481975 461410
rect 479934 461352 481914 461408
rect 481970 461352 481975 461408
rect 479934 461350 481975 461352
rect 52269 461138 52335 461141
rect 52269 461136 60076 461138
rect 52269 461080 52274 461136
rect 52330 461080 60076 461136
rect 479934 461108 479994 461350
rect 481909 461347 481975 461350
rect 52269 461078 60076 461080
rect 52269 461075 52335 461078
rect 482093 460730 482159 460733
rect 479934 460728 482159 460730
rect 479934 460672 482098 460728
rect 482154 460672 482159 460728
rect 479934 460670 482159 460672
rect 52361 460594 52427 460597
rect 52361 460592 60076 460594
rect 52361 460536 52366 460592
rect 52422 460536 60076 460592
rect 479934 460564 479994 460670
rect 482093 460667 482159 460670
rect 52361 460534 60076 460536
rect 52361 460531 52427 460534
rect 487102 460186 487108 460188
rect 479934 460126 487108 460186
rect 45093 460050 45159 460053
rect 45093 460048 60076 460050
rect 45093 459992 45098 460048
rect 45154 459992 60076 460048
rect 479934 460020 479994 460126
rect 487102 460124 487108 460126
rect 487172 460124 487178 460188
rect 45093 459990 60076 459992
rect 45093 459987 45159 459990
rect 43713 459506 43779 459509
rect 43713 459504 60076 459506
rect 43713 459448 43718 459504
rect 43774 459448 60076 459504
rect 43713 459446 60076 459448
rect 43713 459443 43779 459446
rect 479934 459370 479994 459476
rect 482093 459370 482159 459373
rect 479934 459368 482159 459370
rect 479934 459312 482098 459368
rect 482154 459312 482159 459368
rect 479934 459310 482159 459312
rect 482093 459307 482159 459310
rect 489494 459098 489500 459100
rect 479934 459038 489500 459098
rect 46749 458962 46815 458965
rect 46749 458960 60076 458962
rect 46749 458904 46754 458960
rect 46810 458904 60076 458960
rect 479934 458932 479994 459038
rect 489494 459036 489500 459038
rect 489564 459036 489570 459100
rect 46749 458902 60076 458904
rect 46749 458899 46815 458902
rect 482001 458690 482067 458693
rect 479934 458688 482067 458690
rect 479934 458632 482006 458688
rect 482062 458632 482067 458688
rect 479934 458630 482067 458632
rect 46657 458418 46723 458421
rect 46657 458416 60076 458418
rect 46657 458360 46662 458416
rect 46718 458360 60076 458416
rect 479934 458388 479994 458630
rect 482001 458627 482067 458630
rect 46657 458358 60076 458360
rect 46657 458355 46723 458358
rect 583520 458146 584960 458236
rect 509190 458086 584960 458146
rect 482093 458010 482159 458013
rect 479934 458008 482159 458010
rect 479934 457952 482098 458008
rect 482154 457952 482159 458008
rect 479934 457950 482159 457952
rect 46238 457812 46244 457876
rect 46308 457874 46314 457876
rect 46308 457814 60076 457874
rect 479934 457844 479994 457950
rect 482093 457947 482159 457950
rect 46308 457812 46314 457814
rect 482001 457602 482067 457605
rect 479934 457600 482067 457602
rect 479934 457544 482006 457600
rect 482062 457544 482067 457600
rect 479934 457542 482067 457544
rect 46790 457268 46796 457332
rect 46860 457330 46866 457332
rect 46860 457270 60076 457330
rect 479934 457300 479994 457542
rect 482001 457539 482067 457542
rect 500217 457466 500283 457469
rect 508037 457466 508103 457469
rect 509190 457466 509250 458086
rect 583520 457996 584960 458086
rect 500217 457464 509250 457466
rect 500217 457408 500222 457464
rect 500278 457408 508042 457464
rect 508098 457408 509250 457464
rect 500217 457406 509250 457408
rect 500217 457403 500283 457406
rect 508037 457403 508103 457406
rect 46860 457268 46866 457270
rect 46422 456860 46428 456924
rect 46492 456922 46498 456924
rect 46565 456922 46631 456925
rect 46492 456920 46631 456922
rect 46492 456864 46570 456920
rect 46626 456864 46631 456920
rect 46492 456862 46631 456864
rect 46492 456860 46498 456862
rect 46565 456859 46631 456862
rect 48221 456786 48287 456789
rect 48221 456784 60076 456786
rect 48221 456728 48226 456784
rect 48282 456728 60076 456784
rect 48221 456726 60076 456728
rect 48221 456723 48287 456726
rect 479934 456650 479994 456756
rect 482093 456650 482159 456653
rect 479934 456648 482159 456650
rect 479934 456592 482098 456648
rect 482154 456592 482159 456648
rect 479934 456590 482159 456592
rect 482093 456587 482159 456590
rect 484342 456378 484348 456380
rect 479934 456318 484348 456378
rect 50838 456180 50844 456244
rect 50908 456242 50914 456244
rect 50908 456182 60076 456242
rect 479934 456212 479994 456318
rect 484342 456316 484348 456318
rect 484412 456316 484418 456380
rect 50908 456180 50914 456182
rect 485814 455834 485820 455836
rect 479934 455774 485820 455834
rect 48129 455698 48195 455701
rect 48129 455696 60076 455698
rect 48129 455640 48134 455696
rect 48190 455640 60076 455696
rect 479934 455668 479994 455774
rect 485814 455772 485820 455774
rect 485884 455772 485890 455836
rect 48129 455638 60076 455640
rect 48129 455635 48195 455638
rect 482093 455290 482159 455293
rect 479934 455288 482159 455290
rect 479934 455232 482098 455288
rect 482154 455232 482159 455288
rect 479934 455230 482159 455232
rect 48446 455092 48452 455156
rect 48516 455154 48522 455156
rect 48516 455094 60076 455154
rect 479934 455124 479994 455230
rect 482093 455227 482159 455230
rect 48516 455092 48522 455094
rect 482001 454882 482067 454885
rect 479934 454880 482067 454882
rect 479934 454824 482006 454880
rect 482062 454824 482067 454880
rect 479934 454822 482067 454824
rect 59670 454548 59676 454612
rect 59740 454610 59746 454612
rect 59740 454550 60076 454610
rect 479934 454580 479994 454822
rect 482001 454819 482067 454822
rect 59740 454548 59746 454550
rect 479934 454142 480270 454202
rect 48630 454004 48636 454068
rect 48700 454066 48706 454068
rect 48700 454006 60076 454066
rect 479934 454036 479994 454142
rect 480210 454066 480270 454142
rect 485998 454066 486004 454068
rect 480210 454006 486004 454066
rect 48700 454004 48706 454006
rect 485998 454004 486004 454006
rect 486068 454004 486074 454068
rect 482093 453794 482159 453797
rect 479934 453792 482159 453794
rect 479934 453736 482098 453792
rect 482154 453736 482159 453792
rect 479934 453734 482159 453736
rect 52310 453460 52316 453524
rect 52380 453522 52386 453524
rect 52380 453462 60076 453522
rect 479934 453492 479994 453734
rect 482093 453731 482159 453734
rect 52380 453460 52386 453462
rect 479425 453250 479491 453253
rect 479382 453248 479491 453250
rect 479382 453192 479430 453248
rect 479486 453192 479491 453248
rect 479382 453187 479491 453192
rect 48078 452916 48084 452980
rect 48148 452978 48154 452980
rect 48148 452918 60076 452978
rect 479382 452948 479442 453187
rect 48148 452916 48154 452918
rect 482093 452570 482159 452573
rect 479934 452568 482159 452570
rect 479934 452512 482098 452568
rect 482154 452512 482159 452568
rect 479934 452510 482159 452512
rect 47526 452372 47532 452436
rect 47596 452434 47602 452436
rect 47596 452374 60076 452434
rect 479934 452404 479994 452510
rect 482093 452507 482159 452510
rect 47596 452372 47602 452374
rect 47710 451828 47716 451892
rect 47780 451890 47786 451892
rect 47780 451830 60076 451890
rect 47780 451828 47786 451830
rect 479374 451828 479380 451892
rect 479444 451828 479450 451892
rect 482093 451618 482159 451621
rect 479934 451616 482159 451618
rect 479934 451560 482098 451616
rect 482154 451560 482159 451616
rect 479934 451558 482159 451560
rect 58382 451284 58388 451348
rect 58452 451346 58458 451348
rect 58452 451286 60076 451346
rect 479934 451316 479994 451558
rect 482093 451555 482159 451558
rect 58452 451284 58458 451286
rect 34278 450740 34284 450804
rect 34348 450802 34354 450804
rect 34348 450742 60076 450802
rect 34348 450740 34354 450742
rect 479934 450666 479994 450772
rect 483422 450666 483428 450668
rect 479934 450606 483428 450666
rect 483422 450604 483428 450606
rect 483492 450604 483498 450668
rect 39614 450196 39620 450260
rect 39684 450258 39690 450260
rect 39684 450198 60076 450258
rect 39684 450196 39690 450198
rect 479934 450122 479994 450228
rect 487286 450122 487292 450124
rect 479934 450062 487292 450122
rect 487286 450060 487292 450062
rect 487356 450060 487362 450124
rect 479517 449986 479583 449989
rect 482185 449986 482251 449989
rect 479517 449984 482251 449986
rect 479517 449928 479522 449984
rect 479578 449928 482190 449984
rect 482246 449928 482251 449984
rect 479517 449926 482251 449928
rect 479517 449923 479583 449926
rect 482185 449923 482251 449926
rect 482185 449850 482251 449853
rect 479934 449848 482251 449850
rect 479934 449792 482190 449848
rect 482246 449792 482251 449848
rect 479934 449790 482251 449792
rect -960 449578 480 449668
rect 37222 449652 37228 449716
rect 37292 449714 37298 449716
rect 37292 449654 60076 449714
rect 479934 449684 479994 449790
rect 482185 449787 482251 449790
rect 37292 449652 37298 449654
rect 3550 449578 3556 449580
rect -960 449518 3556 449578
rect -960 449428 480 449518
rect 3550 449516 3556 449518
rect 3620 449516 3626 449580
rect 482093 449442 482159 449445
rect 479934 449440 482159 449442
rect 479934 449384 482098 449440
rect 482154 449384 482159 449440
rect 479934 449382 482159 449384
rect 58566 449108 58572 449172
rect 58636 449170 58642 449172
rect 58636 449110 60076 449170
rect 479934 449140 479994 449382
rect 482093 449379 482159 449382
rect 58636 449108 58642 449110
rect 482185 448898 482251 448901
rect 479934 448896 482251 448898
rect 479934 448840 482190 448896
rect 482246 448840 482251 448896
rect 479934 448838 482251 448840
rect 31518 448564 31524 448628
rect 31588 448626 31594 448628
rect 31588 448566 60076 448626
rect 479934 448596 479994 448838
rect 482185 448835 482251 448838
rect 31588 448564 31594 448566
rect 482185 448354 482251 448357
rect 479934 448352 482251 448354
rect 479934 448296 482190 448352
rect 482246 448296 482251 448352
rect 479934 448294 482251 448296
rect 30230 448020 30236 448084
rect 30300 448082 30306 448084
rect 30300 448022 60076 448082
rect 479934 448052 479994 448294
rect 482185 448291 482251 448294
rect 30300 448020 30306 448022
rect 482093 447946 482159 447949
rect 480210 447944 482159 447946
rect 480210 447888 482098 447944
rect 482154 447888 482159 447944
rect 480210 447886 482159 447888
rect 480210 447810 480270 447886
rect 482093 447883 482159 447886
rect 479934 447750 480270 447810
rect 31150 447476 31156 447540
rect 31220 447538 31226 447540
rect 31220 447478 60076 447538
rect 479934 447508 479994 447750
rect 31220 447476 31226 447478
rect 55990 446932 55996 446996
rect 56060 446994 56066 446996
rect 482185 446994 482251 446997
rect 56060 446934 60076 446994
rect 480210 446992 482251 446994
rect 56060 446932 56066 446934
rect 479934 446858 479994 446964
rect 480210 446936 482190 446992
rect 482246 446936 482251 446992
rect 480210 446934 482251 446936
rect 480210 446858 480270 446934
rect 482185 446931 482251 446934
rect 479934 446798 480270 446858
rect 482001 446722 482067 446725
rect 479934 446720 482067 446722
rect 479934 446664 482006 446720
rect 482062 446664 482067 446720
rect 479934 446662 482067 446664
rect 47894 446388 47900 446452
rect 47964 446450 47970 446452
rect 47964 446390 60076 446450
rect 479934 446420 479994 446662
rect 482001 446659 482067 446662
rect 47964 446388 47970 446390
rect 482093 446178 482159 446181
rect 479934 446176 482159 446178
rect 479934 446120 482098 446176
rect 482154 446120 482159 446176
rect 479934 446118 482159 446120
rect 32990 445844 32996 445908
rect 33060 445906 33066 445908
rect 33060 445846 60076 445906
rect 479934 445876 479994 446118
rect 482093 446115 482159 446118
rect 33060 445844 33066 445846
rect 482185 445498 482251 445501
rect 479934 445496 482251 445498
rect 479934 445440 482190 445496
rect 482246 445440 482251 445496
rect 479934 445438 482251 445440
rect 46606 445300 46612 445364
rect 46676 445362 46682 445364
rect 46676 445302 60076 445362
rect 479934 445332 479994 445438
rect 482185 445435 482251 445438
rect 46676 445300 46682 445302
rect 482093 445226 482159 445229
rect 480210 445224 482159 445226
rect 480210 445168 482098 445224
rect 482154 445168 482159 445224
rect 480210 445166 482159 445168
rect 480210 445090 480270 445166
rect 482093 445163 482159 445166
rect 479934 445030 480270 445090
rect 59118 444756 59124 444820
rect 59188 444818 59194 444820
rect 59188 444758 60076 444818
rect 479934 444788 479994 445030
rect 59188 444756 59194 444758
rect 583520 444668 584960 444908
rect 34094 444212 34100 444276
rect 34164 444274 34170 444276
rect 482185 444274 482251 444277
rect 34164 444214 60076 444274
rect 480210 444272 482251 444274
rect 34164 444212 34170 444214
rect 479934 444138 479994 444244
rect 480210 444216 482190 444272
rect 482246 444216 482251 444272
rect 480210 444214 482251 444216
rect 480210 444138 480270 444214
rect 482185 444211 482251 444214
rect 479934 444078 480270 444138
rect 482093 444002 482159 444005
rect 479934 444000 482159 444002
rect 479934 443944 482098 444000
rect 482154 443944 482159 444000
rect 479934 443942 482159 443944
rect 57646 443668 57652 443732
rect 57716 443730 57722 443732
rect 57716 443670 60076 443730
rect 479934 443700 479994 443942
rect 482093 443939 482159 443942
rect 57716 443668 57722 443670
rect 32622 443124 32628 443188
rect 32692 443186 32698 443188
rect 499614 443186 499620 443188
rect 32692 443126 60076 443186
rect 32692 443124 32698 443126
rect 479934 443050 479994 443156
rect 480210 443126 499620 443186
rect 480210 443050 480270 443126
rect 499614 443124 499620 443126
rect 499684 443124 499690 443188
rect 479934 442990 480270 443050
rect 482185 442778 482251 442781
rect 479934 442776 482251 442778
rect 479934 442720 482190 442776
rect 482246 442720 482251 442776
rect 479934 442718 482251 442720
rect 58934 442580 58940 442644
rect 59004 442642 59010 442644
rect 59004 442582 60076 442642
rect 479934 442612 479994 442718
rect 482185 442715 482251 442718
rect 59004 442580 59010 442582
rect 37406 442036 37412 442100
rect 37476 442098 37482 442100
rect 511022 442098 511028 442100
rect 37476 442038 60076 442098
rect 37476 442036 37482 442038
rect 479934 441962 479994 442068
rect 480210 442038 511028 442098
rect 480210 441962 480270 442038
rect 511022 442036 511028 442038
rect 511092 442036 511098 442100
rect 479934 441902 480270 441962
rect 36854 441492 36860 441556
rect 36924 441554 36930 441556
rect 510838 441554 510844 441556
rect 36924 441494 60076 441554
rect 36924 441492 36930 441494
rect 479934 441418 479994 441524
rect 480210 441494 510844 441554
rect 480210 441418 480270 441494
rect 510838 441492 510844 441494
rect 510908 441492 510914 441556
rect 479934 441358 480270 441418
rect 482093 441282 482159 441285
rect 479934 441280 482159 441282
rect 479934 441224 482098 441280
rect 482154 441224 482159 441280
rect 479934 441222 482159 441224
rect 35566 440948 35572 441012
rect 35636 441010 35642 441012
rect 35636 440950 60076 441010
rect 479934 440980 479994 441222
rect 482093 441219 482159 441222
rect 35636 440948 35642 440950
rect 482185 440738 482251 440741
rect 479934 440736 482251 440738
rect 479934 440680 482190 440736
rect 482246 440680 482251 440736
rect 479934 440678 482251 440680
rect 31334 440404 31340 440468
rect 31404 440466 31410 440468
rect 31404 440406 60076 440466
rect 479934 440436 479994 440678
rect 482185 440675 482251 440678
rect 31404 440404 31410 440406
rect 482185 440058 482251 440061
rect 479934 440056 482251 440058
rect 479934 440000 482190 440056
rect 482246 440000 482251 440056
rect 479934 439998 482251 440000
rect 32806 439860 32812 439924
rect 32876 439922 32882 439924
rect 32876 439862 60076 439922
rect 479934 439892 479994 439998
rect 482185 439995 482251 439998
rect 32876 439860 32882 439862
rect 53598 439316 53604 439380
rect 53668 439378 53674 439380
rect 494278 439378 494284 439380
rect 53668 439318 60076 439378
rect 53668 439316 53674 439318
rect 479934 439242 479994 439348
rect 480210 439318 494284 439378
rect 480210 439242 480270 439318
rect 494278 439316 494284 439318
rect 494348 439316 494354 439380
rect 479934 439182 480270 439242
rect 37038 438772 37044 438836
rect 37108 438834 37114 438836
rect 482185 438834 482251 438837
rect 37108 438774 60076 438834
rect 480210 438832 482251 438834
rect 37108 438772 37114 438774
rect 479934 438698 479994 438804
rect 480210 438776 482190 438832
rect 482246 438776 482251 438832
rect 480210 438774 482251 438776
rect 480210 438698 480270 438774
rect 482185 438771 482251 438774
rect 479934 438638 480270 438698
rect 482093 438562 482159 438565
rect 479934 438560 482159 438562
rect 479934 438504 482098 438560
rect 482154 438504 482159 438560
rect 479934 438502 482159 438504
rect 35750 438228 35756 438292
rect 35820 438290 35826 438292
rect 35820 438230 60076 438290
rect 479934 438260 479994 438502
rect 482093 438499 482159 438502
rect 35820 438228 35826 438230
rect 50337 437746 50403 437749
rect 490465 437746 490531 437749
rect 50337 437744 60076 437746
rect 50337 437688 50342 437744
rect 50398 437688 60076 437744
rect 480210 437744 490531 437746
rect 50337 437686 60076 437688
rect 50337 437683 50403 437686
rect 479934 437610 479994 437716
rect 480210 437688 490470 437744
rect 490526 437688 490531 437744
rect 480210 437686 490531 437688
rect 480210 437610 480270 437686
rect 490465 437683 490531 437686
rect 479934 437550 480270 437610
rect 34237 437202 34303 437205
rect 34237 437200 60076 437202
rect 34237 437144 34242 437200
rect 34298 437144 60076 437200
rect 34237 437142 60076 437144
rect 34237 437139 34303 437142
rect 479934 437066 479994 437172
rect 483749 437066 483815 437069
rect 479934 437064 483815 437066
rect 479934 437008 483754 437064
rect 483810 437008 483815 437064
rect 479934 437006 483815 437008
rect 483749 437003 483815 437006
rect -960 436508 480 436748
rect 49141 436658 49207 436661
rect 49141 436656 60076 436658
rect 49141 436600 49146 436656
rect 49202 436600 60076 436656
rect 49141 436598 60076 436600
rect 49141 436595 49207 436598
rect 479934 436522 479994 436628
rect 484761 436522 484827 436525
rect 479934 436520 484827 436522
rect 479934 436464 484766 436520
rect 484822 436464 484827 436520
rect 479934 436462 484827 436464
rect 484761 436459 484827 436462
rect 60181 436386 60247 436389
rect 60181 436384 60290 436386
rect 60181 436328 60186 436384
rect 60242 436328 60290 436384
rect 60181 436323 60290 436328
rect 60230 436084 60290 436323
rect 483657 436250 483723 436253
rect 479934 436248 483723 436250
rect 479934 436192 483662 436248
rect 483718 436192 483723 436248
rect 479934 436190 483723 436192
rect 479934 436084 479994 436190
rect 483657 436187 483723 436190
rect 48957 435570 49023 435573
rect 48957 435568 60076 435570
rect 48957 435512 48962 435568
rect 49018 435512 60076 435568
rect 48957 435510 60076 435512
rect 48957 435507 49023 435510
rect 479934 435434 479994 435540
rect 486325 435434 486391 435437
rect 479934 435432 486391 435434
rect 479934 435376 486330 435432
rect 486386 435376 486391 435432
rect 479934 435374 486391 435376
rect 486325 435371 486391 435374
rect 50245 435026 50311 435029
rect 50245 435024 60076 435026
rect 50245 434968 50250 435024
rect 50306 434968 60076 435024
rect 50245 434966 60076 434968
rect 50245 434963 50311 434966
rect 479934 434890 479994 434996
rect 484945 434890 485011 434893
rect 479934 434888 485011 434890
rect 479934 434832 484950 434888
rect 485006 434832 485011 434888
rect 479934 434830 485011 434832
rect 484945 434827 485011 434830
rect 49049 434482 49115 434485
rect 490373 434482 490439 434485
rect 49049 434480 60076 434482
rect 49049 434424 49054 434480
rect 49110 434424 60076 434480
rect 480210 434480 490439 434482
rect 49049 434422 60076 434424
rect 49049 434419 49115 434422
rect 479934 434346 479994 434452
rect 480210 434424 490378 434480
rect 490434 434424 490439 434480
rect 480210 434422 490439 434424
rect 480210 434346 480270 434422
rect 490373 434419 490439 434422
rect 479934 434286 480270 434346
rect 52913 433938 52979 433941
rect 52913 433936 60076 433938
rect 52913 433880 52918 433936
rect 52974 433880 60076 433936
rect 52913 433878 60076 433880
rect 52913 433875 52979 433878
rect 479934 433802 479994 433908
rect 486601 433802 486667 433805
rect 479934 433800 486667 433802
rect 479934 433744 486606 433800
rect 486662 433744 486667 433800
rect 479934 433742 486667 433744
rect 486601 433739 486667 433742
rect 486417 433530 486483 433533
rect 479934 433528 486483 433530
rect 479934 433472 486422 433528
rect 486478 433472 486483 433528
rect 479934 433470 486483 433472
rect 49509 433394 49575 433397
rect 49509 433392 60076 433394
rect 49509 433336 49514 433392
rect 49570 433336 60076 433392
rect 479934 433364 479994 433470
rect 486417 433467 486483 433470
rect 49509 433334 60076 433336
rect 49509 433331 49575 433334
rect 49233 432850 49299 432853
rect 49233 432848 60076 432850
rect 49233 432792 49238 432848
rect 49294 432792 60076 432848
rect 49233 432790 60076 432792
rect 49233 432787 49299 432790
rect 479934 432714 479994 432820
rect 485037 432714 485103 432717
rect 479934 432712 485103 432714
rect 479934 432656 485042 432712
rect 485098 432656 485103 432712
rect 479934 432654 485103 432656
rect 485037 432651 485103 432654
rect 51533 432306 51599 432309
rect 51533 432304 60076 432306
rect 51533 432248 51538 432304
rect 51594 432248 60076 432304
rect 51533 432246 60076 432248
rect 51533 432243 51599 432246
rect 479934 432170 479994 432276
rect 483565 432170 483631 432173
rect 479934 432168 483631 432170
rect 479934 432112 483570 432168
rect 483626 432112 483631 432168
rect 479934 432110 483631 432112
rect 483565 432107 483631 432110
rect 49417 431762 49483 431765
rect 49417 431760 60076 431762
rect 49417 431704 49422 431760
rect 49478 431704 60076 431760
rect 49417 431702 60076 431704
rect 49417 431699 49483 431702
rect 479934 431626 479994 431732
rect 486509 431626 486575 431629
rect 479934 431624 486575 431626
rect 479934 431568 486514 431624
rect 486570 431568 486575 431624
rect 479934 431566 486575 431568
rect 486509 431563 486575 431566
rect 580625 431626 580691 431629
rect 583520 431626 584960 431716
rect 580625 431624 584960 431626
rect 580625 431568 580630 431624
rect 580686 431568 584960 431624
rect 580625 431566 584960 431568
rect 580625 431563 580691 431566
rect 583520 431476 584960 431566
rect 50061 431218 50127 431221
rect 50061 431216 60076 431218
rect 50061 431160 50066 431216
rect 50122 431160 60076 431216
rect 50061 431158 60076 431160
rect 50061 431155 50127 431158
rect 479934 431082 479994 431188
rect 484393 431082 484459 431085
rect 479934 431080 484459 431082
rect 479934 431024 484398 431080
rect 484454 431024 484459 431080
rect 479934 431022 484459 431024
rect 484393 431019 484459 431022
rect 483473 430810 483539 430813
rect 479934 430808 483539 430810
rect 479934 430752 483478 430808
rect 483534 430752 483539 430808
rect 479934 430750 483539 430752
rect 57697 430674 57763 430677
rect 57697 430672 60076 430674
rect 57697 430616 57702 430672
rect 57758 430616 60076 430672
rect 479934 430644 479994 430750
rect 483473 430747 483539 430750
rect 57697 430614 60076 430616
rect 57697 430611 57763 430614
rect 60089 430402 60155 430405
rect 60046 430400 60155 430402
rect 60046 430344 60094 430400
rect 60150 430344 60155 430400
rect 60046 430339 60155 430344
rect 60046 430100 60106 430339
rect 479934 429994 479994 430100
rect 484669 429994 484735 429997
rect 479934 429992 484735 429994
rect 479934 429936 484674 429992
rect 484730 429936 484735 429992
rect 479934 429934 484735 429936
rect 484669 429931 484735 429934
rect 60273 429858 60339 429861
rect 60230 429856 60339 429858
rect 60230 429800 60278 429856
rect 60334 429800 60339 429856
rect 60230 429795 60339 429800
rect 60230 429556 60290 429795
rect 479934 429450 479994 429556
rect 484485 429450 484551 429453
rect 479934 429448 484551 429450
rect 479934 429392 484490 429448
rect 484546 429392 484551 429448
rect 479934 429390 484551 429392
rect 484485 429387 484551 429390
rect 58893 429042 58959 429045
rect 58893 429040 60076 429042
rect 58893 428984 58898 429040
rect 58954 428984 60076 429040
rect 58893 428982 60076 428984
rect 58893 428979 58959 428982
rect 479934 428906 479994 429012
rect 484577 428906 484643 428909
rect 479934 428904 484643 428906
rect 479934 428848 484582 428904
rect 484638 428848 484643 428904
rect 479934 428846 484643 428848
rect 484577 428843 484643 428846
rect 34329 428498 34395 428501
rect 34329 428496 60076 428498
rect 34329 428440 34334 428496
rect 34390 428440 60076 428496
rect 34329 428438 60076 428440
rect 34329 428435 34395 428438
rect 479934 428362 479994 428468
rect 483381 428362 483447 428365
rect 479934 428360 483447 428362
rect 479934 428304 483386 428360
rect 483442 428304 483447 428360
rect 479934 428302 483447 428304
rect 483381 428299 483447 428302
rect 484853 428090 484919 428093
rect 479934 428088 484919 428090
rect 479934 428032 484858 428088
rect 484914 428032 484919 428088
rect 479934 428030 484919 428032
rect 36721 427954 36787 427957
rect 36721 427952 60076 427954
rect 36721 427896 36726 427952
rect 36782 427896 60076 427952
rect 479934 427924 479994 428030
rect 484853 428027 484919 428030
rect 36721 427894 60076 427896
rect 36721 427891 36787 427894
rect 34145 427410 34211 427413
rect 501229 427410 501295 427413
rect 34145 427408 60076 427410
rect 34145 427352 34150 427408
rect 34206 427352 60076 427408
rect 480210 427408 501295 427410
rect 34145 427350 60076 427352
rect 34145 427347 34211 427350
rect 479934 427274 479994 427380
rect 480210 427352 501234 427408
rect 501290 427352 501295 427408
rect 480210 427350 501295 427352
rect 480210 427274 480270 427350
rect 501229 427347 501295 427350
rect 479934 427214 480270 427274
rect 42425 426866 42491 426869
rect 42425 426864 60076 426866
rect 42425 426808 42430 426864
rect 42486 426808 60076 426864
rect 42425 426806 60076 426808
rect 42425 426803 42491 426806
rect 479934 426730 479994 426836
rect 483197 426730 483263 426733
rect 479934 426728 483263 426730
rect 479934 426672 483202 426728
rect 483258 426672 483263 426728
rect 479934 426670 483263 426672
rect 483197 426667 483263 426670
rect 35525 426322 35591 426325
rect 35525 426320 60076 426322
rect 35525 426264 35530 426320
rect 35586 426264 60076 426320
rect 35525 426262 60076 426264
rect 35525 426259 35591 426262
rect 479934 426186 479994 426292
rect 483289 426186 483355 426189
rect 479934 426184 483355 426186
rect 479934 426128 483294 426184
rect 483350 426128 483355 426184
rect 479934 426126 483355 426128
rect 483289 426123 483355 426126
rect 51625 425778 51691 425781
rect 51625 425776 60076 425778
rect 51625 425720 51630 425776
rect 51686 425720 60076 425776
rect 51625 425718 60076 425720
rect 51625 425715 51691 425718
rect 479934 425642 479994 425748
rect 489177 425642 489243 425645
rect 479934 425640 489243 425642
rect 479934 425584 489182 425640
rect 489238 425584 489243 425640
rect 479934 425582 489243 425584
rect 489177 425579 489243 425582
rect 47393 425234 47459 425237
rect 490281 425234 490347 425237
rect 47393 425232 60076 425234
rect 47393 425176 47398 425232
rect 47454 425176 60076 425232
rect 480210 425232 490347 425234
rect 47393 425174 60076 425176
rect 47393 425171 47459 425174
rect 479934 425098 479994 425204
rect 480210 425176 490286 425232
rect 490342 425176 490347 425232
rect 480210 425174 490347 425176
rect 480210 425098 480270 425174
rect 490281 425171 490347 425174
rect 479934 425038 480270 425098
rect 482829 424826 482895 424829
rect 479934 424824 482895 424826
rect 479934 424768 482834 424824
rect 482890 424768 482895 424824
rect 479934 424766 482895 424768
rect 47669 424690 47735 424693
rect 47669 424688 60076 424690
rect 47669 424632 47674 424688
rect 47730 424632 60076 424688
rect 479934 424660 479994 424766
rect 482829 424763 482895 424766
rect 47669 424630 60076 424632
rect 47669 424627 47735 424630
rect 482185 424554 482251 424557
rect 480210 424552 482251 424554
rect 480210 424496 482190 424552
rect 482246 424496 482251 424552
rect 480210 424494 482251 424496
rect 480210 424418 480270 424494
rect 482185 424491 482251 424494
rect 479934 424358 480270 424418
rect 47761 424146 47827 424149
rect 47761 424144 60076 424146
rect 47761 424088 47766 424144
rect 47822 424088 60076 424144
rect 479934 424116 479994 424358
rect 47761 424086 60076 424088
rect 47761 424083 47827 424086
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 47945 423602 48011 423605
rect 47945 423600 60076 423602
rect 47945 423544 47950 423600
rect 48006 423544 60076 423600
rect 47945 423542 60076 423544
rect 47945 423539 48011 423542
rect 479934 423466 479994 423572
rect 482829 423466 482895 423469
rect 479934 423464 482895 423466
rect 479934 423408 482834 423464
rect 482890 423408 482895 423464
rect 479934 423406 482895 423408
rect 482829 423403 482895 423406
rect 482829 423330 482895 423333
rect 479934 423328 482895 423330
rect 479934 423272 482834 423328
rect 482890 423272 482895 423328
rect 479934 423270 482895 423272
rect 50521 423058 50587 423061
rect 50521 423056 60076 423058
rect 50521 423000 50526 423056
rect 50582 423000 60076 423056
rect 479934 423028 479994 423270
rect 482829 423267 482895 423270
rect 50521 422998 60076 423000
rect 50521 422995 50587 422998
rect 48865 422514 48931 422517
rect 492121 422514 492187 422517
rect 48865 422512 60076 422514
rect 48865 422456 48870 422512
rect 48926 422456 60076 422512
rect 480210 422512 492187 422514
rect 48865 422454 60076 422456
rect 48865 422451 48931 422454
rect 479934 422378 479994 422484
rect 480210 422456 492126 422512
rect 492182 422456 492187 422512
rect 480210 422454 492187 422456
rect 480210 422378 480270 422454
rect 492121 422451 492187 422454
rect 479934 422318 480270 422378
rect 486233 422106 486299 422109
rect 479934 422104 486299 422106
rect 479934 422048 486238 422104
rect 486294 422048 486299 422104
rect 479934 422046 486299 422048
rect 49325 421970 49391 421973
rect 49325 421968 60076 421970
rect 49325 421912 49330 421968
rect 49386 421912 60076 421968
rect 479934 421940 479994 422046
rect 486233 422043 486299 422046
rect 49325 421910 60076 421912
rect 49325 421907 49391 421910
rect 483841 421562 483907 421565
rect 479934 421560 483907 421562
rect 479934 421504 483846 421560
rect 483902 421504 483907 421560
rect 479934 421502 483907 421504
rect 50705 421426 50771 421429
rect 50705 421424 60076 421426
rect 50705 421368 50710 421424
rect 50766 421368 60076 421424
rect 479934 421396 479994 421502
rect 483841 421499 483907 421502
rect 50705 421366 60076 421368
rect 50705 421363 50771 421366
rect 50429 420882 50495 420885
rect 50429 420880 60076 420882
rect 50429 420824 50434 420880
rect 50490 420824 60076 420880
rect 50429 420822 60076 420824
rect 50429 420819 50495 420822
rect 479934 420746 479994 420852
rect 483238 420746 483244 420748
rect 479934 420686 483244 420746
rect 483238 420684 483244 420686
rect 483308 420684 483314 420748
rect 40769 420338 40835 420341
rect 499941 420338 500007 420341
rect 40769 420336 60076 420338
rect 40769 420280 40774 420336
rect 40830 420280 60076 420336
rect 480210 420336 500007 420338
rect 40769 420278 60076 420280
rect 40769 420275 40835 420278
rect 479934 420202 479994 420308
rect 480210 420280 499946 420336
rect 500002 420280 500007 420336
rect 480210 420278 500007 420280
rect 480210 420202 480270 420278
rect 499941 420275 500007 420278
rect 479934 420142 480270 420202
rect 483606 420140 483612 420204
rect 483676 420202 483682 420204
rect 543406 420202 543412 420204
rect 483676 420142 543412 420202
rect 483676 420140 483682 420142
rect 543406 420140 543412 420142
rect 543476 420140 543482 420204
rect 56225 419794 56291 419797
rect 498561 419794 498627 419797
rect 56225 419792 60076 419794
rect 56225 419736 56230 419792
rect 56286 419736 60076 419792
rect 480210 419792 498627 419794
rect 56225 419734 60076 419736
rect 56225 419731 56291 419734
rect 479934 419658 479994 419764
rect 480210 419736 498566 419792
rect 498622 419736 498627 419792
rect 480210 419734 498627 419736
rect 480210 419658 480270 419734
rect 498561 419731 498627 419734
rect 479934 419598 480270 419658
rect 55857 419250 55923 419253
rect 499757 419250 499823 419253
rect 55857 419248 60076 419250
rect 55857 419192 55862 419248
rect 55918 419192 60076 419248
rect 480210 419248 499823 419250
rect 55857 419190 60076 419192
rect 55857 419187 55923 419190
rect 479934 419114 479994 419220
rect 480210 419192 499762 419248
rect 499818 419192 499823 419248
rect 480210 419190 499823 419192
rect 480210 419114 480270 419190
rect 499757 419187 499823 419190
rect 479934 419054 480270 419114
rect 39481 418706 39547 418709
rect 495617 418706 495683 418709
rect 39481 418704 60076 418706
rect 39481 418648 39486 418704
rect 39542 418648 60076 418704
rect 480210 418704 495683 418706
rect 39481 418646 60076 418648
rect 39481 418643 39547 418646
rect 479934 418570 479994 418676
rect 480210 418648 495622 418704
rect 495678 418648 495683 418704
rect 480210 418646 495683 418648
rect 480210 418570 480270 418646
rect 495617 418643 495683 418646
rect 479934 418510 480270 418570
rect 558126 418236 558132 418300
rect 558196 418298 558202 418300
rect 583520 418298 584960 418388
rect 558196 418238 584960 418298
rect 558196 418236 558202 418238
rect 46381 418162 46447 418165
rect 46381 418160 60076 418162
rect 46381 418104 46386 418160
rect 46442 418104 60076 418160
rect 583520 418148 584960 418238
rect 46381 418102 60076 418104
rect 46381 418099 46447 418102
rect 479934 418026 479994 418132
rect 482829 418026 482895 418029
rect 479934 418024 482895 418026
rect 479934 417968 482834 418024
rect 482890 417968 482895 418024
rect 479934 417966 482895 417968
rect 482829 417963 482895 417966
rect 51717 417618 51783 417621
rect 491569 417618 491635 417621
rect 51717 417616 60076 417618
rect 51717 417560 51722 417616
rect 51778 417560 60076 417616
rect 480210 417616 491635 417618
rect 51717 417558 60076 417560
rect 51717 417555 51783 417558
rect 479934 417482 479994 417588
rect 480210 417560 491574 417616
rect 491630 417560 491635 417616
rect 480210 417558 491635 417560
rect 480210 417482 480270 417558
rect 491569 417555 491635 417558
rect 479934 417422 480270 417482
rect 482185 417346 482251 417349
rect 479934 417344 482251 417346
rect 479934 417288 482190 417344
rect 482246 417288 482251 417344
rect 479934 417286 482251 417288
rect 46289 417074 46355 417077
rect 46289 417072 60076 417074
rect 46289 417016 46294 417072
rect 46350 417016 60076 417072
rect 479934 417044 479994 417286
rect 482185 417283 482251 417286
rect 46289 417014 60076 417016
rect 46289 417011 46355 417014
rect 482829 416666 482895 416669
rect 479934 416664 482895 416666
rect 479934 416608 482834 416664
rect 482890 416608 482895 416664
rect 479934 416606 482895 416608
rect 42374 416468 42380 416532
rect 42444 416530 42450 416532
rect 42444 416470 60076 416530
rect 479934 416500 479994 416606
rect 482829 416603 482895 416606
rect 42444 416468 42450 416470
rect 44030 415924 44036 415988
rect 44100 415986 44106 415988
rect 498142 415986 498148 415988
rect 44100 415926 60076 415986
rect 44100 415924 44106 415926
rect 479934 415850 479994 415956
rect 480210 415926 498148 415986
rect 480210 415850 480270 415926
rect 498142 415924 498148 415926
rect 498212 415924 498218 415988
rect 479934 415790 480270 415850
rect 479934 415518 480270 415578
rect 43294 415380 43300 415444
rect 43364 415442 43370 415444
rect 43364 415382 60076 415442
rect 479934 415412 479994 415518
rect 480210 415442 480270 415518
rect 495801 415442 495867 415445
rect 480210 415440 495867 415442
rect 480210 415384 495806 415440
rect 495862 415384 495867 415440
rect 480210 415382 495867 415384
rect 43364 415380 43370 415382
rect 495801 415379 495867 415382
rect 482829 415170 482895 415173
rect 479934 415168 482895 415170
rect 479934 415112 482834 415168
rect 482890 415112 482895 415168
rect 479934 415110 482895 415112
rect 43846 414836 43852 414900
rect 43916 414898 43922 414900
rect 43916 414838 60076 414898
rect 479934 414868 479994 415110
rect 482829 415107 482895 415110
rect 43916 414836 43922 414838
rect 482185 414626 482251 414629
rect 479934 414624 482251 414626
rect 479934 414568 482190 414624
rect 482246 414568 482251 414624
rect 479934 414566 482251 414568
rect 44950 414292 44956 414356
rect 45020 414354 45026 414356
rect 45020 414294 60076 414354
rect 479934 414324 479994 414566
rect 482185 414563 482251 414566
rect 45020 414292 45026 414294
rect 479934 413886 480270 413946
rect 46422 413748 46428 413812
rect 46492 413810 46498 413812
rect 46492 413750 60076 413810
rect 479934 413780 479994 413886
rect 480210 413810 480270 413886
rect 482829 413810 482895 413813
rect 480210 413808 482895 413810
rect 480210 413752 482834 413808
rect 482890 413752 482895 413808
rect 480210 413750 482895 413752
rect 46492 413748 46498 413750
rect 482829 413747 482895 413750
rect 482185 413674 482251 413677
rect 480210 413672 482251 413674
rect 480210 413616 482190 413672
rect 482246 413616 482251 413672
rect 480210 413614 482251 413616
rect 480210 413538 480270 413614
rect 482185 413611 482251 413614
rect 479934 413478 480270 413538
rect 42558 413204 42564 413268
rect 42628 413266 42634 413268
rect 42628 413206 60076 413266
rect 479934 413236 479994 413478
rect 42628 413204 42634 413206
rect 481081 412994 481147 412997
rect 479934 412992 481147 412994
rect 479934 412936 481086 412992
rect 481142 412936 481147 412992
rect 479934 412934 481147 412936
rect 55949 412722 56015 412725
rect 55949 412720 60076 412722
rect 55949 412664 55954 412720
rect 56010 412664 60076 412720
rect 479934 412692 479994 412934
rect 481081 412931 481147 412934
rect 55949 412662 60076 412664
rect 55949 412659 56015 412662
rect 482829 412450 482895 412453
rect 479934 412448 482895 412450
rect 479934 412392 482834 412448
rect 482890 412392 482895 412448
rect 479934 412390 482895 412392
rect 53005 412178 53071 412181
rect 53005 412176 60076 412178
rect 53005 412120 53010 412176
rect 53066 412120 60076 412176
rect 479934 412148 479994 412390
rect 482829 412387 482895 412390
rect 53005 412118 60076 412120
rect 53005 412115 53071 412118
rect 479609 411906 479675 411909
rect 479566 411904 479675 411906
rect 479566 411848 479614 411904
rect 479670 411848 479675 411904
rect 479566 411843 479675 411848
rect 54477 411634 54543 411637
rect 54477 411632 60076 411634
rect 54477 411576 54482 411632
rect 54538 411576 60076 411632
rect 479566 411604 479626 411843
rect 54477 411574 60076 411576
rect 54477 411571 54543 411574
rect 39573 411090 39639 411093
rect 482185 411090 482251 411093
rect 39573 411088 60076 411090
rect 39573 411032 39578 411088
rect 39634 411032 60076 411088
rect 480210 411088 482251 411090
rect 39573 411030 60076 411032
rect 39573 411027 39639 411030
rect 479934 410954 479994 411060
rect 480210 411032 482190 411088
rect 482246 411032 482251 411088
rect 480210 411030 482251 411032
rect 480210 410954 480270 411030
rect 482185 411027 482251 411030
rect 479934 410894 480270 410954
rect 482185 410818 482251 410821
rect 479934 410816 482251 410818
rect 479934 410760 482190 410816
rect 482246 410760 482251 410816
rect 479934 410758 482251 410760
rect -960 410546 480 410636
rect 3734 410546 3740 410548
rect -960 410486 3740 410546
rect -960 410396 480 410486
rect 3734 410484 3740 410486
rect 3804 410484 3810 410548
rect 53097 410546 53163 410549
rect 53097 410544 60076 410546
rect 53097 410488 53102 410544
rect 53158 410488 60076 410544
rect 479934 410516 479994 410758
rect 482185 410755 482251 410758
rect 53097 410486 60076 410488
rect 53097 410483 53163 410486
rect 482829 410410 482895 410413
rect 480210 410408 482895 410410
rect 480210 410352 482834 410408
rect 482890 410352 482895 410408
rect 480210 410350 482895 410352
rect 480210 410274 480270 410350
rect 482829 410347 482895 410350
rect 479934 410214 480270 410274
rect 2998 409940 3004 410004
rect 3068 410002 3074 410004
rect 4061 410002 4127 410005
rect 3068 410000 4127 410002
rect 3068 409944 4066 410000
rect 4122 409944 4127 410000
rect 3068 409942 4127 409944
rect 3068 409940 3074 409942
rect 4061 409939 4127 409942
rect 54385 410002 54451 410005
rect 54385 410000 60076 410002
rect 54385 409944 54390 410000
rect 54446 409944 60076 410000
rect 479934 409972 479994 410214
rect 54385 409942 60076 409944
rect 54385 409939 54451 409942
rect 482829 409594 482895 409597
rect 479934 409592 482895 409594
rect 479934 409536 482834 409592
rect 482890 409536 482895 409592
rect 479934 409534 482895 409536
rect 53189 409458 53255 409461
rect 53189 409456 60076 409458
rect 53189 409400 53194 409456
rect 53250 409400 60076 409456
rect 479934 409428 479994 409534
rect 482829 409531 482895 409534
rect 53189 409398 60076 409400
rect 53189 409395 53255 409398
rect 40861 408914 40927 408917
rect 40861 408912 60076 408914
rect 40861 408856 40866 408912
rect 40922 408856 60076 408912
rect 40861 408854 60076 408856
rect 40861 408851 40927 408854
rect 479934 408778 479994 408884
rect 487705 408778 487771 408781
rect 479934 408776 487771 408778
rect 479934 408720 487710 408776
rect 487766 408720 487771 408776
rect 479934 408718 487771 408720
rect 487705 408715 487771 408718
rect 479934 408446 480270 408506
rect 42517 408370 42583 408373
rect 42517 408368 60076 408370
rect 42517 408312 42522 408368
rect 42578 408312 60076 408368
rect 479934 408340 479994 408446
rect 480210 408370 480270 408446
rect 482185 408370 482251 408373
rect 480210 408368 482251 408370
rect 42517 408310 60076 408312
rect 480210 408312 482190 408368
rect 482246 408312 482251 408368
rect 480210 408310 482251 408312
rect 42517 408307 42583 408310
rect 482185 408307 482251 408310
rect 480989 408234 481055 408237
rect 480210 408232 481055 408234
rect 480210 408176 480994 408232
rect 481050 408176 481055 408232
rect 480210 408174 481055 408176
rect 480210 408098 480270 408174
rect 480989 408171 481055 408174
rect 479934 408038 480270 408098
rect 41045 407826 41111 407829
rect 41045 407824 60076 407826
rect 41045 407768 41050 407824
rect 41106 407768 60076 407824
rect 479934 407796 479994 408038
rect 41045 407766 60076 407768
rect 41045 407763 41111 407766
rect 482829 407554 482895 407557
rect 479934 407552 482895 407554
rect 479934 407496 482834 407552
rect 482890 407496 482895 407552
rect 479934 407494 482895 407496
rect 54753 407282 54819 407285
rect 54753 407280 60076 407282
rect 54753 407224 54758 407280
rect 54814 407224 60076 407280
rect 479934 407252 479994 407494
rect 482829 407491 482895 407494
rect 54753 407222 60076 407224
rect 54753 407219 54819 407222
rect 482829 406874 482895 406877
rect 479934 406872 482895 406874
rect 479934 406816 482834 406872
rect 482890 406816 482895 406872
rect 479934 406814 482895 406816
rect 56041 406738 56107 406741
rect 56041 406736 60076 406738
rect 56041 406680 56046 406736
rect 56102 406680 60076 406736
rect 479934 406708 479994 406814
rect 482829 406811 482895 406814
rect 56041 406678 60076 406680
rect 56041 406675 56107 406678
rect 482185 406602 482251 406605
rect 480210 406600 482251 406602
rect 480210 406544 482190 406600
rect 482246 406544 482251 406600
rect 480210 406542 482251 406544
rect 480210 406466 480270 406542
rect 482185 406539 482251 406542
rect 479934 406406 480270 406466
rect 54845 406194 54911 406197
rect 54845 406192 60076 406194
rect 54845 406136 54850 406192
rect 54906 406136 60076 406192
rect 479934 406164 479994 406406
rect 54845 406134 60076 406136
rect 54845 406131 54911 406134
rect 40953 405650 41019 405653
rect 480529 405650 480595 405653
rect 40953 405648 60076 405650
rect 40953 405592 40958 405648
rect 41014 405592 60076 405648
rect 480210 405648 480595 405650
rect 40953 405590 60076 405592
rect 40953 405587 41019 405590
rect 479934 405514 479994 405620
rect 480210 405592 480534 405648
rect 480590 405592 480595 405648
rect 480210 405590 480595 405592
rect 480210 405514 480270 405590
rect 480529 405587 480595 405590
rect 479934 405454 480270 405514
rect 479793 405242 479859 405245
rect 507853 405242 507919 405245
rect 479793 405240 509250 405242
rect 479793 405184 479798 405240
rect 479854 405184 507858 405240
rect 507914 405184 509250 405240
rect 479793 405182 509250 405184
rect 479793 405179 479859 405182
rect 507853 405179 507919 405182
rect 54661 405106 54727 405109
rect 498377 405106 498443 405109
rect 54661 405104 60076 405106
rect 54661 405048 54666 405104
rect 54722 405048 60076 405104
rect 480210 405104 498443 405106
rect 54661 405046 60076 405048
rect 54661 405043 54727 405046
rect 479934 404970 479994 405076
rect 480210 405048 498382 405104
rect 498438 405048 498443 405104
rect 480210 405046 498443 405048
rect 480210 404970 480270 405046
rect 498377 405043 498443 405046
rect 479934 404910 480270 404970
rect 509190 404970 509250 405182
rect 583520 404970 584960 405060
rect 509190 404910 584960 404970
rect 482829 404834 482895 404837
rect 479934 404832 482895 404834
rect 479934 404776 482834 404832
rect 482890 404776 482895 404832
rect 583520 404820 584960 404910
rect 479934 404774 482895 404776
rect 54569 404562 54635 404565
rect 54569 404560 60076 404562
rect 54569 404504 54574 404560
rect 54630 404504 60076 404560
rect 479934 404532 479994 404774
rect 482829 404771 482895 404774
rect 54569 404502 60076 404504
rect 54569 404499 54635 404502
rect 480621 404290 480687 404293
rect 479934 404288 480687 404290
rect 479934 404232 480626 404288
rect 480682 404232 480687 404288
rect 479934 404230 480687 404232
rect 56409 404018 56475 404021
rect 56409 404016 60076 404018
rect 56409 403960 56414 404016
rect 56470 403960 60076 404016
rect 479934 403988 479994 404230
rect 480621 404227 480687 404230
rect 56409 403958 60076 403960
rect 56409 403955 56475 403958
rect 480805 403746 480871 403749
rect 479934 403744 480871 403746
rect 479934 403688 480810 403744
rect 480866 403688 480871 403744
rect 479934 403686 480871 403688
rect 45185 403474 45251 403477
rect 45185 403472 60076 403474
rect 45185 403416 45190 403472
rect 45246 403416 60076 403472
rect 479934 403444 479994 403686
rect 480805 403683 480871 403686
rect 45185 403414 60076 403416
rect 45185 403411 45251 403414
rect 479609 403066 479675 403069
rect 481766 403066 481772 403068
rect 479609 403064 481772 403066
rect 479609 403008 479614 403064
rect 479670 403008 481772 403064
rect 479609 403006 481772 403008
rect 479609 403003 479675 403006
rect 481766 403004 481772 403006
rect 481836 403004 481842 403068
rect 41137 402930 41203 402933
rect 480713 402930 480779 402933
rect 41137 402928 60076 402930
rect 41137 402872 41142 402928
rect 41198 402872 60076 402928
rect 480210 402928 480779 402930
rect 41137 402870 60076 402872
rect 41137 402867 41203 402870
rect 479934 402794 479994 402900
rect 480210 402872 480718 402928
rect 480774 402872 480779 402928
rect 480210 402870 480779 402872
rect 480210 402794 480270 402870
rect 480713 402867 480779 402870
rect 479934 402734 480270 402794
rect 480897 402658 480963 402661
rect 479934 402656 480963 402658
rect 479934 402600 480902 402656
rect 480958 402600 480963 402656
rect 479934 402598 480963 402600
rect 44081 402386 44147 402389
rect 44081 402384 60076 402386
rect 44081 402328 44086 402384
rect 44142 402328 60076 402384
rect 479934 402356 479994 402598
rect 480897 402595 480963 402598
rect 44081 402326 60076 402328
rect 44081 402323 44147 402326
rect 482829 402114 482895 402117
rect 479934 402112 482895 402114
rect 479934 402056 482834 402112
rect 482890 402056 482895 402112
rect 479934 402054 482895 402056
rect 43805 401842 43871 401845
rect 43805 401840 60076 401842
rect 43805 401784 43810 401840
rect 43866 401784 60076 401840
rect 479934 401812 479994 402054
rect 482829 402051 482895 402054
rect 43805 401782 60076 401784
rect 43805 401779 43871 401782
rect 482829 401434 482895 401437
rect 479934 401432 482895 401434
rect 479934 401376 482834 401432
rect 482890 401376 482895 401432
rect 479934 401374 482895 401376
rect 56317 401298 56383 401301
rect 56317 401296 60076 401298
rect 56317 401240 56322 401296
rect 56378 401240 60076 401296
rect 479934 401268 479994 401374
rect 482829 401371 482895 401374
rect 56317 401238 60076 401240
rect 56317 401235 56383 401238
rect 482829 401026 482895 401029
rect 479934 401024 482895 401026
rect 479934 400968 482834 401024
rect 482890 400968 482895 401024
rect 479934 400966 482895 400968
rect 51901 400754 51967 400757
rect 51901 400752 60076 400754
rect 51901 400696 51906 400752
rect 51962 400696 60076 400752
rect 479934 400724 479994 400966
rect 482829 400963 482895 400966
rect 51901 400694 60076 400696
rect 51901 400691 51967 400694
rect 51809 400210 51875 400213
rect 51809 400208 60076 400210
rect 51809 400152 51814 400208
rect 51870 400152 60076 400208
rect 51809 400150 60076 400152
rect 51809 400147 51875 400150
rect 479934 400074 479994 400180
rect 486366 400074 486372 400076
rect 479934 400014 486372 400074
rect 486366 400012 486372 400014
rect 486436 400012 486442 400076
rect 482829 399938 482895 399941
rect 479934 399936 482895 399938
rect 479934 399880 482834 399936
rect 482890 399880 482895 399936
rect 479934 399878 482895 399880
rect 41229 399666 41295 399669
rect 41229 399664 60076 399666
rect 41229 399608 41234 399664
rect 41290 399608 60076 399664
rect 479934 399636 479994 399878
rect 482829 399875 482895 399878
rect 41229 399606 60076 399608
rect 41229 399603 41295 399606
rect 482185 399394 482251 399397
rect 479934 399392 482251 399394
rect 479934 399336 482190 399392
rect 482246 399336 482251 399392
rect 479934 399334 482251 399336
rect 39665 399122 39731 399125
rect 39665 399120 60076 399122
rect 39665 399064 39670 399120
rect 39726 399064 60076 399120
rect 479934 399092 479994 399334
rect 482185 399331 482251 399334
rect 39665 399062 60076 399064
rect 39665 399059 39731 399062
rect 482829 398714 482895 398717
rect 479934 398712 482895 398714
rect 479934 398656 482834 398712
rect 482890 398656 482895 398712
rect 479934 398654 482895 398656
rect 38469 398578 38535 398581
rect 38469 398576 60076 398578
rect 38469 398520 38474 398576
rect 38530 398520 60076 398576
rect 479934 398548 479994 398654
rect 482829 398651 482895 398654
rect 38469 398518 60076 398520
rect 38469 398515 38535 398518
rect 482001 398442 482067 398445
rect 480210 398440 482067 398442
rect 480210 398384 482006 398440
rect 482062 398384 482067 398440
rect 480210 398382 482067 398384
rect 480210 398306 480270 398382
rect 482001 398379 482067 398382
rect 479934 398246 480270 398306
rect 2814 398108 2820 398172
rect 2884 398170 2890 398172
rect 3969 398170 4035 398173
rect 2884 398168 4035 398170
rect 2884 398112 3974 398168
rect 4030 398112 4035 398168
rect 2884 398110 4035 398112
rect 2884 398108 2890 398110
rect 3969 398107 4035 398110
rect 48037 398034 48103 398037
rect 48037 398032 60076 398034
rect 48037 397976 48042 398032
rect 48098 397976 60076 398032
rect 479934 398004 479994 398246
rect 48037 397974 60076 397976
rect 48037 397971 48103 397974
rect 482185 397762 482251 397765
rect 479934 397760 482251 397762
rect 479934 397704 482190 397760
rect 482246 397704 482251 397760
rect 479934 397702 482251 397704
rect -960 397490 480 397580
rect 3918 397490 3924 397492
rect -960 397430 3924 397490
rect -960 397340 480 397430
rect 3918 397428 3924 397430
rect 3988 397428 3994 397492
rect 53373 397490 53439 397493
rect 53373 397488 60076 397490
rect 53373 397432 53378 397488
rect 53434 397432 60076 397488
rect 479934 397460 479994 397702
rect 482185 397699 482251 397702
rect 53373 397430 60076 397432
rect 53373 397427 53439 397430
rect 482829 397218 482895 397221
rect 479934 397216 482895 397218
rect 479934 397160 482834 397216
rect 482890 397160 482895 397216
rect 479934 397158 482895 397160
rect 39757 396946 39823 396949
rect 39757 396944 60076 396946
rect 39757 396888 39762 396944
rect 39818 396888 60076 396944
rect 479934 396916 479994 397158
rect 482829 397155 482895 397158
rect 39757 396886 60076 396888
rect 39757 396883 39823 396886
rect 482185 396674 482251 396677
rect 479934 396672 482251 396674
rect 479934 396616 482190 396672
rect 482246 396616 482251 396672
rect 479934 396614 482251 396616
rect 54937 396402 55003 396405
rect 54937 396400 60076 396402
rect 54937 396344 54942 396400
rect 54998 396344 60076 396400
rect 479934 396372 479994 396614
rect 482185 396611 482251 396614
rect 54937 396342 60076 396344
rect 54937 396339 55003 396342
rect 479934 395934 480270 395994
rect 43897 395858 43963 395861
rect 43897 395856 60076 395858
rect 43897 395800 43902 395856
rect 43958 395800 60076 395856
rect 479934 395828 479994 395934
rect 480210 395858 480270 395934
rect 482829 395858 482895 395861
rect 480210 395856 482895 395858
rect 43897 395798 60076 395800
rect 480210 395800 482834 395856
rect 482890 395800 482895 395856
rect 480210 395798 482895 395800
rect 43897 395795 43963 395798
rect 482829 395795 482895 395798
rect 482185 395722 482251 395725
rect 480210 395720 482251 395722
rect 480210 395664 482190 395720
rect 482246 395664 482251 395720
rect 480210 395662 482251 395664
rect 480210 395586 480270 395662
rect 482185 395659 482251 395662
rect 479934 395526 480270 395586
rect 28901 395314 28967 395317
rect 28901 395312 60076 395314
rect 28901 395256 28906 395312
rect 28962 395256 60076 395312
rect 479934 395284 479994 395526
rect 28901 395254 60076 395256
rect 28901 395251 28967 395254
rect 489310 394906 489316 394908
rect 479934 394846 489316 394906
rect 45277 394770 45343 394773
rect 45277 394768 60076 394770
rect 45277 394712 45282 394768
rect 45338 394712 60076 394768
rect 479934 394740 479994 394846
rect 489310 394844 489316 394846
rect 489380 394844 489386 394908
rect 45277 394710 60076 394712
rect 45277 394707 45343 394710
rect 482829 394362 482895 394365
rect 479934 394360 482895 394362
rect 479934 394304 482834 394360
rect 482890 394304 482895 394360
rect 479934 394302 482895 394304
rect 46841 394226 46907 394229
rect 46841 394224 60076 394226
rect 46841 394168 46846 394224
rect 46902 394168 60076 394224
rect 479934 394196 479994 394302
rect 482829 394299 482895 394302
rect 46841 394166 60076 394168
rect 46841 394163 46907 394166
rect 482185 393954 482251 393957
rect 479934 393952 482251 393954
rect 479934 393896 482190 393952
rect 482246 393896 482251 393952
rect 479934 393894 482251 393896
rect 45461 393682 45527 393685
rect 45461 393680 60076 393682
rect 45461 393624 45466 393680
rect 45522 393624 60076 393680
rect 479934 393652 479994 393894
rect 482185 393891 482251 393894
rect 45461 393622 60076 393624
rect 45461 393619 45527 393622
rect 482829 393274 482895 393277
rect 479934 393272 482895 393274
rect 479934 393216 482834 393272
rect 482890 393216 482895 393272
rect 479934 393214 482895 393216
rect 45369 393138 45435 393141
rect 45369 393136 60076 393138
rect 45369 393080 45374 393136
rect 45430 393080 60076 393136
rect 479934 393108 479994 393214
rect 482829 393211 482895 393214
rect 45369 393078 60076 393080
rect 45369 393075 45435 393078
rect 482921 392866 482987 392869
rect 479934 392864 482987 392866
rect 479934 392808 482926 392864
rect 482982 392808 482987 392864
rect 479934 392806 482987 392808
rect 57329 392594 57395 392597
rect 57329 392592 60076 392594
rect 57329 392536 57334 392592
rect 57390 392536 60076 392592
rect 479934 392564 479994 392806
rect 482921 392803 482987 392806
rect 57329 392534 60076 392536
rect 57329 392531 57395 392534
rect 482093 392322 482159 392325
rect 479934 392320 482159 392322
rect 479934 392264 482098 392320
rect 482154 392264 482159 392320
rect 479934 392262 482159 392264
rect 37181 392050 37247 392053
rect 37181 392048 60076 392050
rect 37181 391992 37186 392048
rect 37242 391992 60076 392048
rect 479934 392020 479994 392262
rect 482093 392259 482159 392262
rect 37181 391990 60076 391992
rect 37181 391987 37247 391990
rect 482921 391642 482987 391645
rect 479934 391640 482987 391642
rect 479934 391584 482926 391640
rect 482982 391584 482987 391640
rect 583520 391628 584960 391868
rect 479934 391582 482987 391584
rect 35801 391506 35867 391509
rect 35801 391504 60076 391506
rect 35801 391448 35806 391504
rect 35862 391448 60076 391504
rect 479934 391476 479994 391582
rect 482921 391579 482987 391582
rect 35801 391446 60076 391448
rect 35801 391443 35867 391446
rect 482829 391234 482895 391237
rect 479934 391232 482895 391234
rect 479934 391176 482834 391232
rect 482890 391176 482895 391232
rect 479934 391174 482895 391176
rect 34421 390962 34487 390965
rect 34421 390960 60076 390962
rect 34421 390904 34426 390960
rect 34482 390904 60076 390960
rect 479934 390932 479994 391174
rect 482829 391171 482895 391174
rect 34421 390902 60076 390904
rect 34421 390899 34487 390902
rect 31661 390418 31727 390421
rect 482921 390418 482987 390421
rect 31661 390416 60076 390418
rect 31661 390360 31666 390416
rect 31722 390360 60076 390416
rect 480210 390416 482987 390418
rect 31661 390358 60076 390360
rect 31661 390355 31727 390358
rect 479934 390282 479994 390388
rect 480210 390360 482926 390416
rect 482982 390360 482987 390416
rect 480210 390358 482987 390360
rect 480210 390282 480270 390358
rect 482921 390355 482987 390358
rect 479934 390222 480270 390282
rect 94129 390146 94195 390149
rect 500217 390146 500283 390149
rect 94129 390144 500283 390146
rect 94129 390088 94134 390144
rect 94190 390088 500222 390144
rect 500278 390088 500283 390144
rect 94129 390086 500283 390088
rect 94129 390083 94195 390086
rect 500217 390083 500283 390086
rect 59169 389194 59235 389197
rect 476113 389194 476179 389197
rect 479517 389194 479583 389197
rect 59169 389192 59370 389194
rect 59169 389136 59174 389192
rect 59230 389136 59370 389192
rect 59169 389134 59370 389136
rect 59169 389131 59235 389134
rect 59310 389058 59370 389134
rect 476113 389192 479583 389194
rect 476113 389136 476118 389192
rect 476174 389136 479522 389192
rect 479578 389136 479583 389192
rect 476113 389134 479583 389136
rect 476113 389131 476179 389134
rect 479517 389131 479583 389134
rect 60733 389058 60799 389061
rect 59310 389056 60799 389058
rect 59310 389000 60738 389056
rect 60794 389000 60799 389056
rect 59310 388998 60799 389000
rect 60733 388995 60799 388998
rect 97257 389058 97323 389061
rect 503069 389058 503135 389061
rect 97257 389056 503135 389058
rect 97257 389000 97262 389056
rect 97318 389000 503074 389056
rect 503130 389000 503135 389056
rect 97257 388998 503135 389000
rect 97257 388995 97323 388998
rect 503069 388995 503135 388998
rect 101305 388922 101371 388925
rect 503805 388922 503871 388925
rect 101305 388920 503871 388922
rect 101305 388864 101310 388920
rect 101366 388864 503810 388920
rect 503866 388864 503871 388920
rect 101305 388862 503871 388864
rect 101305 388859 101371 388862
rect 503805 388859 503871 388862
rect 90541 388786 90607 388789
rect 473169 388786 473235 388789
rect 90541 388784 473235 388786
rect 90541 388728 90546 388784
rect 90602 388728 473174 388784
rect 473230 388728 473235 388784
rect 90541 388726 473235 388728
rect 90541 388723 90607 388726
rect 473169 388723 473235 388726
rect 473353 388786 473419 388789
rect 479558 388786 479564 388788
rect 473353 388784 479564 388786
rect 473353 388728 473358 388784
rect 473414 388728 479564 388784
rect 473353 388726 479564 388728
rect 473353 388723 473419 388726
rect 479558 388724 479564 388726
rect 479628 388724 479634 388788
rect 166257 388650 166323 388653
rect 545113 388650 545179 388653
rect 166257 388648 545179 388650
rect 166257 388592 166262 388648
rect 166318 388592 545118 388648
rect 545174 388592 545179 388648
rect 166257 388590 545179 388592
rect 166257 388587 166323 388590
rect 545113 388587 545179 388590
rect 234521 388514 234587 388517
rect 473261 388514 473327 388517
rect 234521 388512 473327 388514
rect 234521 388456 234526 388512
rect 234582 388456 473266 388512
rect 473322 388456 473327 388512
rect 234521 388454 473327 388456
rect 234521 388451 234587 388454
rect 473261 388451 473327 388454
rect 473537 388514 473603 388517
rect 476113 388514 476179 388517
rect 473537 388512 476179 388514
rect 473537 388456 473542 388512
rect 473598 388456 476118 388512
rect 476174 388456 476179 388512
rect 473537 388454 476179 388456
rect 473537 388451 473603 388454
rect 476113 388451 476179 388454
rect 235533 388378 235599 388381
rect 482185 388378 482251 388381
rect 235533 388376 482251 388378
rect 235533 388320 235538 388376
rect 235594 388320 482190 388376
rect 482246 388320 482251 388376
rect 235533 388318 482251 388320
rect 235533 388315 235599 388318
rect 482185 388315 482251 388318
rect 473169 388242 473235 388245
rect 479793 388242 479859 388245
rect 473169 388240 479859 388242
rect 473169 388184 473174 388240
rect 473230 388184 479798 388240
rect 479854 388184 479859 388240
rect 473169 388182 479859 388184
rect 473169 388179 473235 388182
rect 479793 388179 479859 388182
rect 231761 387834 231827 387837
rect 474641 387834 474707 387837
rect 231761 387832 474707 387834
rect 231761 387776 231766 387832
rect 231822 387776 474646 387832
rect 474702 387776 474707 387832
rect 231761 387774 474707 387776
rect 231761 387771 231827 387774
rect 474641 387771 474707 387774
rect 60641 387698 60707 387701
rect 122833 387698 122899 387701
rect 60641 387696 122899 387698
rect 60641 387640 60646 387696
rect 60702 387640 122838 387696
rect 122894 387640 122899 387696
rect 60641 387638 122899 387640
rect 60641 387635 60707 387638
rect 122833 387635 122899 387638
rect 249885 387698 249951 387701
rect 348877 387698 348943 387701
rect 249885 387696 348943 387698
rect 249885 387640 249890 387696
rect 249946 387640 348882 387696
rect 348938 387640 348943 387696
rect 249885 387638 348943 387640
rect 249885 387635 249951 387638
rect 348877 387635 348943 387638
rect 452929 387698 452995 387701
rect 482277 387698 482343 387701
rect 452929 387696 482343 387698
rect 452929 387640 452934 387696
rect 452990 387640 482282 387696
rect 482338 387640 482343 387696
rect 452929 387638 482343 387640
rect 452929 387635 452995 387638
rect 482277 387635 482343 387638
rect 55070 387500 55076 387564
rect 55140 387562 55146 387564
rect 125593 387562 125659 387565
rect 126421 387562 126487 387565
rect 55140 387560 126487 387562
rect 55140 387504 125598 387560
rect 125654 387504 126426 387560
rect 126482 387504 126487 387560
rect 55140 387502 126487 387504
rect 55140 387500 55146 387502
rect 125593 387499 125659 387502
rect 126421 387499 126487 387502
rect 251909 387562 251975 387565
rect 356053 387562 356119 387565
rect 251909 387560 356119 387562
rect 251909 387504 251914 387560
rect 251970 387504 356058 387560
rect 356114 387504 356119 387560
rect 251909 387502 356119 387504
rect 251909 387499 251975 387502
rect 356053 387499 356119 387502
rect 417417 387562 417483 387565
rect 449341 387562 449407 387565
rect 417417 387560 449407 387562
rect 417417 387504 417422 387560
rect 417478 387504 449346 387560
rect 449402 387504 449407 387560
rect 417417 387502 449407 387504
rect 417417 387499 417483 387502
rect 449341 387499 449407 387502
rect 60457 387426 60523 387429
rect 62113 387426 62179 387429
rect 129733 387426 129799 387429
rect 60457 387424 62179 387426
rect 60457 387368 60462 387424
rect 60518 387368 62118 387424
rect 62174 387368 62179 387424
rect 60457 387366 62179 387368
rect 60457 387363 60523 387366
rect 62113 387363 62179 387366
rect 64830 387424 129799 387426
rect 64830 387368 129738 387424
rect 129794 387368 129799 387424
rect 64830 387366 129799 387368
rect 59261 387290 59327 387293
rect 64830 387290 64890 387366
rect 129733 387363 129799 387366
rect 150433 387426 150499 387429
rect 158713 387426 158779 387429
rect 150433 387424 158779 387426
rect 150433 387368 150438 387424
rect 150494 387368 158718 387424
rect 158774 387368 158779 387424
rect 150433 387366 158779 387368
rect 150433 387363 150499 387366
rect 158713 387363 158779 387366
rect 239213 387426 239279 387429
rect 259177 387426 259243 387429
rect 239213 387424 259243 387426
rect 239213 387368 239218 387424
rect 239274 387368 259182 387424
rect 259238 387368 259243 387424
rect 239213 387366 259243 387368
rect 239213 387363 239279 387366
rect 259177 387363 259243 387366
rect 270125 387426 270191 387429
rect 420637 387426 420703 387429
rect 270125 387424 420703 387426
rect 270125 387368 270130 387424
rect 270186 387368 420642 387424
rect 420698 387368 420703 387424
rect 270125 387366 420703 387368
rect 270125 387363 270191 387366
rect 420637 387363 420703 387366
rect 59261 387288 64890 387290
rect 59261 387232 59266 387288
rect 59322 387232 64890 387288
rect 59261 387230 64890 387232
rect 119337 387290 119403 387293
rect 270401 387290 270467 387293
rect 119337 387288 270467 387290
rect 119337 387232 119342 387288
rect 119398 387232 270406 387288
rect 270462 387232 270467 387288
rect 119337 387230 270467 387232
rect 59261 387227 59327 387230
rect 119337 387227 119403 387230
rect 270401 387227 270467 387230
rect 273161 387290 273227 387293
rect 431401 387290 431467 387293
rect 273161 387288 431467 387290
rect 273161 387232 273166 387288
rect 273222 387232 431406 387288
rect 431462 387232 431467 387288
rect 273161 387230 431467 387232
rect 273161 387227 273227 387230
rect 431401 387227 431467 387230
rect 55673 387154 55739 387157
rect 106181 387154 106247 387157
rect 55673 387152 106247 387154
rect 55673 387096 55678 387152
rect 55734 387096 106186 387152
rect 106242 387096 106247 387152
rect 55673 387094 106247 387096
rect 55673 387091 55739 387094
rect 106181 387091 106247 387094
rect 115289 387154 115355 387157
rect 274633 387154 274699 387157
rect 115289 387152 274699 387154
rect 115289 387096 115294 387152
rect 115350 387096 274638 387152
rect 274694 387096 274699 387152
rect 115289 387094 274699 387096
rect 115289 387091 115355 387094
rect 274633 387091 274699 387094
rect 392577 387154 392643 387157
rect 442165 387154 442231 387157
rect 392577 387152 442231 387154
rect 392577 387096 392582 387152
rect 392638 387096 442170 387152
rect 442226 387096 442231 387152
rect 392577 387094 442231 387096
rect 392577 387091 392643 387094
rect 442165 387091 442231 387094
rect 62573 387018 62639 387021
rect 90541 387018 90607 387021
rect 62573 387016 90607 387018
rect 62573 386960 62578 387016
rect 62634 386960 90546 387016
rect 90602 386960 90607 387016
rect 62573 386958 90607 386960
rect 62573 386955 62639 386958
rect 90541 386955 90607 386958
rect 108389 387018 108455 387021
rect 272517 387018 272583 387021
rect 108389 387016 272583 387018
rect 108389 386960 108394 387016
rect 108450 386960 272522 387016
rect 272578 386960 272583 387016
rect 108389 386958 272583 386960
rect 108389 386955 108455 386958
rect 272517 386955 272583 386958
rect 275185 387018 275251 387021
rect 438577 387018 438643 387021
rect 275185 387016 438643 387018
rect 275185 386960 275190 387016
rect 275246 386960 438582 387016
rect 438638 386960 438643 387016
rect 275185 386958 438643 386960
rect 275185 386955 275251 386958
rect 438577 386955 438643 386958
rect 60917 386882 60983 386885
rect 86953 386882 87019 386885
rect 115841 386882 115907 386885
rect 60917 386880 115907 386882
rect 60917 386824 60922 386880
rect 60978 386824 86958 386880
rect 87014 386824 115846 386880
rect 115902 386824 115907 386880
rect 60917 386822 115907 386824
rect 60917 386819 60983 386822
rect 86953 386819 87019 386822
rect 115841 386819 115907 386822
rect 124121 386882 124187 386885
rect 150433 386882 150499 386885
rect 151537 386882 151603 386885
rect 124121 386880 151603 386882
rect 124121 386824 124126 386880
rect 124182 386824 150438 386880
rect 150494 386824 151542 386880
rect 151598 386824 151603 386880
rect 124121 386822 151603 386824
rect 124121 386819 124187 386822
rect 150433 386819 150499 386822
rect 151537 386819 151603 386822
rect 236453 386882 236519 386885
rect 237649 386882 237715 386885
rect 236453 386880 237715 386882
rect 236453 386824 236458 386880
rect 236514 386824 237654 386880
rect 237710 386824 237715 386880
rect 236453 386822 237715 386824
rect 236453 386819 236519 386822
rect 237649 386819 237715 386822
rect 239029 386882 239095 386885
rect 244825 386882 244891 386885
rect 239029 386880 244891 386882
rect 239029 386824 239034 386880
rect 239090 386824 244830 386880
rect 244886 386824 244891 386880
rect 239029 386822 244891 386824
rect 239029 386819 239095 386822
rect 244825 386819 244891 386822
rect 256049 386882 256115 386885
rect 341701 386882 341767 386885
rect 256049 386880 341767 386882
rect 256049 386824 256054 386880
rect 256110 386824 341706 386880
rect 341762 386824 341767 386880
rect 256049 386822 341767 386824
rect 256049 386819 256115 386822
rect 341701 386819 341767 386822
rect 454677 386882 454743 386885
rect 456517 386882 456583 386885
rect 454677 386880 456583 386882
rect 454677 386824 454682 386880
rect 454738 386824 456522 386880
rect 456578 386824 456583 386880
rect 454677 386822 456583 386824
rect 454677 386819 454743 386822
rect 456517 386819 456583 386822
rect 105629 386746 105695 386749
rect 118693 386746 118759 386749
rect 105629 386744 118759 386746
rect 105629 386688 105634 386744
rect 105690 386688 118698 386744
rect 118754 386688 118759 386744
rect 105629 386686 118759 386688
rect 105629 386683 105695 386686
rect 118693 386683 118759 386686
rect 134517 386746 134583 386749
rect 179413 386746 179479 386749
rect 180241 386746 180307 386749
rect 134517 386744 180307 386746
rect 134517 386688 134522 386744
rect 134578 386688 179418 386744
rect 179474 386688 180246 386744
rect 180302 386688 180307 386744
rect 134517 386686 180307 386688
rect 134517 386683 134583 386686
rect 179413 386683 179479 386686
rect 180241 386683 180307 386686
rect 258717 386746 258783 386749
rect 334525 386746 334591 386749
rect 258717 386744 334591 386746
rect 258717 386688 258722 386744
rect 258778 386688 334530 386744
rect 334586 386688 334591 386744
rect 258717 386686 334591 386688
rect 258717 386683 258783 386686
rect 334525 386683 334591 386686
rect 95693 386610 95759 386613
rect 108297 386610 108363 386613
rect 95693 386608 108363 386610
rect 95693 386552 95698 386608
rect 95754 386552 108302 386608
rect 108358 386552 108363 386608
rect 95693 386550 108363 386552
rect 95693 386547 95759 386550
rect 108297 386547 108363 386550
rect 135897 386610 135963 386613
rect 183829 386610 183895 386613
rect 184841 386610 184907 386613
rect 135897 386608 184907 386610
rect 135897 386552 135902 386608
rect 135958 386552 183834 386608
rect 183890 386552 184846 386608
rect 184902 386552 184907 386608
rect 135897 386550 184907 386552
rect 135897 386547 135963 386550
rect 183829 386547 183895 386550
rect 184841 386547 184907 386550
rect 57789 386474 57855 386477
rect 132585 386474 132651 386477
rect 133597 386474 133663 386477
rect 57789 386472 133663 386474
rect 57789 386416 57794 386472
rect 57850 386416 132590 386472
rect 132646 386416 133602 386472
rect 133658 386416 133663 386472
rect 57789 386414 133663 386416
rect 57789 386411 57855 386414
rect 132585 386411 132651 386414
rect 133597 386411 133663 386414
rect 137277 386474 137343 386477
rect 186957 386474 187023 386477
rect 137277 386472 187023 386474
rect 137277 386416 137282 386472
rect 137338 386416 186962 386472
rect 187018 386416 187023 386472
rect 137277 386414 187023 386416
rect 137277 386411 137343 386414
rect 186957 386411 187023 386414
rect 112069 386338 112135 386341
rect 112437 386338 112503 386341
rect 482829 386338 482895 386341
rect 112069 386336 482895 386338
rect 112069 386280 112074 386336
rect 112130 386280 112442 386336
rect 112498 386280 482834 386336
rect 482890 386280 482895 386336
rect 112069 386278 482895 386280
rect 112069 386275 112135 386278
rect 112437 386275 112503 386278
rect 482829 386275 482895 386278
rect 184841 386202 184907 386205
rect 531957 386202 532023 386205
rect 184841 386200 532023 386202
rect 184841 386144 184846 386200
rect 184902 386144 531962 386200
rect 532018 386144 532023 386200
rect 184841 386142 532023 386144
rect 184841 386139 184907 386142
rect 531957 386139 532023 386142
rect 477493 386066 477559 386069
rect 479701 386066 479767 386069
rect 477493 386064 479767 386066
rect 477493 386008 477498 386064
rect 477554 386008 479706 386064
rect 479762 386008 479767 386064
rect 477493 386006 479767 386008
rect 477493 386003 477559 386006
rect 479701 386003 479767 386006
rect 67541 385658 67607 385661
rect 101305 385658 101371 385661
rect 67541 385656 101371 385658
rect 67541 385600 67546 385656
rect 67602 385600 101310 385656
rect 101366 385600 101371 385656
rect 67541 385598 101371 385600
rect 67541 385595 67607 385598
rect 101305 385595 101371 385598
rect 173157 384978 173223 384981
rect 546677 384978 546743 384981
rect 173157 384976 546743 384978
rect 173157 384920 173162 384976
rect 173218 384920 546682 384976
rect 546738 384920 546743 384976
rect 173157 384918 546743 384920
rect 173157 384915 173223 384918
rect 546677 384915 546743 384918
rect 179413 384842 179479 384845
rect 546585 384842 546651 384845
rect 179413 384840 546651 384842
rect 179413 384784 179418 384840
rect 179474 384784 546590 384840
rect 546646 384784 546651 384840
rect 179413 384782 546651 384784
rect 179413 384779 179479 384782
rect 546585 384779 546651 384782
rect 471237 384706 471303 384709
rect 473261 384706 473327 384709
rect 471237 384704 473327 384706
rect 471237 384648 471242 384704
rect 471298 384648 473266 384704
rect 473322 384648 473327 384704
rect 471237 384646 473327 384648
rect 471237 384643 471303 384646
rect 473261 384643 473327 384646
rect -960 384284 480 384524
rect 282177 384434 282243 384437
rect 541341 384434 541407 384437
rect 282177 384432 541407 384434
rect 282177 384376 282182 384432
rect 282238 384376 541346 384432
rect 541402 384376 541407 384432
rect 282177 384374 541407 384376
rect 282177 384371 282243 384374
rect 541341 384371 541407 384374
rect 3550 384236 3556 384300
rect 3620 384298 3626 384300
rect 210366 384298 210372 384300
rect 3620 384238 210372 384298
rect 3620 384236 3626 384238
rect 210366 384236 210372 384238
rect 210436 384236 210442 384300
rect 239806 384236 239812 384300
rect 239876 384298 239882 384300
rect 452929 384298 452995 384301
rect 239876 384296 452995 384298
rect 239876 384240 452934 384296
rect 452990 384240 452995 384296
rect 239876 384238 452995 384240
rect 239876 384236 239882 384238
rect 452929 384235 452995 384238
rect 60733 383754 60799 383757
rect 60733 383752 62130 383754
rect 60733 383696 60738 383752
rect 60794 383696 62130 383752
rect 60733 383694 62130 383696
rect 60733 383691 60799 383694
rect 62070 383618 62130 383694
rect 63493 383618 63559 383621
rect 62070 383616 63559 383618
rect 62070 383560 63498 383616
rect 63554 383560 63559 383616
rect 62070 383558 63559 383560
rect 63493 383555 63559 383558
rect 169017 383618 169083 383621
rect 543733 383618 543799 383621
rect 169017 383616 543799 383618
rect 169017 383560 169022 383616
rect 169078 383560 543738 383616
rect 543794 383560 543799 383616
rect 169017 383558 543799 383560
rect 169017 383555 169083 383558
rect 543733 383555 543799 383558
rect 186957 383482 187023 383485
rect 536097 383482 536163 383485
rect 186957 383480 536163 383482
rect 186957 383424 186962 383480
rect 187018 383424 536102 383480
rect 536158 383424 536163 383480
rect 186957 383422 536163 383424
rect 186957 383419 187023 383422
rect 536097 383419 536163 383422
rect 233141 383346 233207 383349
rect 482737 383346 482803 383349
rect 233141 383344 482803 383346
rect 233141 383288 233146 383344
rect 233202 383288 482742 383344
rect 482798 383288 482803 383344
rect 233141 383286 482803 383288
rect 233141 383283 233207 383286
rect 482737 383283 482803 383286
rect 282269 383210 282335 383213
rect 541157 383210 541223 383213
rect 282269 383208 541223 383210
rect 282269 383152 282274 383208
rect 282330 383152 541162 383208
rect 541218 383152 541223 383208
rect 282269 383150 541223 383152
rect 282269 383147 282335 383150
rect 541157 383147 541223 383150
rect 233049 383074 233115 383077
rect 505921 383074 505987 383077
rect 233049 383072 505987 383074
rect 233049 383016 233054 383072
rect 233110 383016 505926 383072
rect 505982 383016 505987 383072
rect 233049 383014 505987 383016
rect 233049 383011 233115 383014
rect 505921 383011 505987 383014
rect 3969 382938 4035 382941
rect 214649 382938 214715 382941
rect 3969 382936 214715 382938
rect 3969 382880 3974 382936
rect 4030 382880 214654 382936
rect 214710 382880 214715 382936
rect 3969 382878 214715 382880
rect 3969 382875 4035 382878
rect 214649 382875 214715 382878
rect 231577 382938 231643 382941
rect 508681 382938 508747 382941
rect 231577 382936 508747 382938
rect 231577 382880 231582 382936
rect 231638 382880 508686 382936
rect 508742 382880 508747 382936
rect 231577 382878 508747 382880
rect 231577 382875 231643 382878
rect 508681 382875 508747 382878
rect 239622 382740 239628 382804
rect 239692 382802 239698 382804
rect 305821 382802 305887 382805
rect 239692 382800 305887 382802
rect 239692 382744 305826 382800
rect 305882 382744 305887 382800
rect 239692 382742 305887 382744
rect 239692 382740 239698 382742
rect 305821 382739 305887 382742
rect 469213 382802 469279 382805
rect 477493 382802 477559 382805
rect 469213 382800 477559 382802
rect 469213 382744 469218 382800
rect 469274 382744 477498 382800
rect 477554 382744 477559 382800
rect 469213 382742 477559 382744
rect 469213 382739 469279 382742
rect 477493 382739 477559 382742
rect 257981 381714 258047 381717
rect 377581 381714 377647 381717
rect 257981 381712 377647 381714
rect 257981 381656 257986 381712
rect 258042 381656 377586 381712
rect 377642 381656 377647 381712
rect 257981 381654 377647 381656
rect 257981 381651 258047 381654
rect 377581 381651 377647 381654
rect 3918 381516 3924 381580
rect 3988 381578 3994 381580
rect 206134 381578 206140 381580
rect 3988 381518 206140 381578
rect 3988 381516 3994 381518
rect 206134 381516 206140 381518
rect 206204 381516 206210 381580
rect 282126 381516 282132 381580
rect 282196 381578 282202 381580
rect 541198 381578 541204 381580
rect 282196 381518 541204 381578
rect 282196 381516 282202 381518
rect 541198 381516 541204 381518
rect 541268 381516 541274 381580
rect 541249 381034 541315 381037
rect 541382 381034 541388 381036
rect 541249 381032 541388 381034
rect 541249 380976 541254 381032
rect 541310 380976 541388 381032
rect 541249 380974 541388 380976
rect 541249 380971 541315 380974
rect 541382 380972 541388 380974
rect 541452 380972 541458 381036
rect 232957 380898 233023 380901
rect 510061 380898 510127 380901
rect 232957 380896 510127 380898
rect 232957 380840 232962 380896
rect 233018 380840 510066 380896
rect 510122 380840 510127 380896
rect 232957 380838 510127 380840
rect 232957 380835 233023 380838
rect 510061 380835 510127 380838
rect 228909 380762 228975 380765
rect 512821 380762 512887 380765
rect 228909 380760 512887 380762
rect 228909 380704 228914 380760
rect 228970 380704 512826 380760
rect 512882 380704 512887 380760
rect 228909 380702 512887 380704
rect 228909 380699 228975 380702
rect 512821 380699 512887 380702
rect 230381 380626 230447 380629
rect 515581 380626 515647 380629
rect 230381 380624 515647 380626
rect 230381 380568 230386 380624
rect 230442 380568 515586 380624
rect 515642 380568 515647 380624
rect 230381 380566 515647 380568
rect 230381 380563 230447 380566
rect 515581 380563 515647 380566
rect 231669 380490 231735 380493
rect 516961 380490 517027 380493
rect 231669 380488 517027 380490
rect 231669 380432 231674 380488
rect 231730 380432 516966 380488
rect 517022 380432 517027 380488
rect 231669 380430 517027 380432
rect 231669 380427 231735 380430
rect 516961 380427 517027 380430
rect 228725 380354 228791 380357
rect 514201 380354 514267 380357
rect 228725 380352 514267 380354
rect 228725 380296 228730 380352
rect 228786 380296 514206 380352
rect 514262 380296 514267 380352
rect 228725 380294 514267 380296
rect 228725 380291 228791 380294
rect 514201 380291 514267 380294
rect 228817 380218 228883 380221
rect 519721 380218 519787 380221
rect 228817 380216 519787 380218
rect 228817 380160 228822 380216
rect 228878 380160 519726 380216
rect 519782 380160 519787 380216
rect 228817 380158 519787 380160
rect 228817 380155 228883 380158
rect 519721 380155 519787 380158
rect 234429 380082 234495 380085
rect 500401 380082 500467 380085
rect 234429 380080 500467 380082
rect 234429 380024 234434 380080
rect 234490 380024 500406 380080
rect 500462 380024 500467 380080
rect 234429 380022 500467 380024
rect 234429 380019 234495 380022
rect 500401 380019 500467 380022
rect 281758 379476 281764 379540
rect 281828 379538 281834 379540
rect 282821 379538 282887 379541
rect 281828 379536 282887 379538
rect 281828 379480 282826 379536
rect 282882 379480 282887 379536
rect 281828 379478 282887 379480
rect 281828 379476 281834 379478
rect 282821 379475 282887 379478
rect 271229 378858 271295 378861
rect 417049 378858 417115 378861
rect 271229 378856 417115 378858
rect 271229 378800 271234 378856
rect 271290 378800 417054 378856
rect 417110 378800 417115 378856
rect 271229 378798 417115 378800
rect 271229 378795 271295 378798
rect 417049 378795 417115 378798
rect 230197 378722 230263 378725
rect 528001 378722 528067 378725
rect 230197 378720 528067 378722
rect 230197 378664 230202 378720
rect 230258 378664 528006 378720
rect 528062 378664 528067 378720
rect 230197 378662 528067 378664
rect 230197 378659 230263 378662
rect 528001 378659 528067 378662
rect 236126 378388 236132 378452
rect 236196 378450 236202 378452
rect 583520 378450 584960 378540
rect 236196 378390 584960 378450
rect 236196 378388 236202 378390
rect 583520 378300 584960 378390
rect 3734 377980 3740 378044
rect 3804 378042 3810 378044
rect 284334 378042 284340 378044
rect 3804 377982 284340 378042
rect 3804 377980 3810 377982
rect 284334 377980 284340 377982
rect 284404 377980 284410 378044
rect 467097 378042 467163 378045
rect 469213 378042 469279 378045
rect 467097 378040 469279 378042
rect 467097 377984 467102 378040
rect 467158 377984 469218 378040
rect 469274 377984 469279 378040
rect 467097 377982 469279 377984
rect 467097 377979 467163 377982
rect 469213 377979 469279 377982
rect 235073 377906 235139 377909
rect 525241 377906 525307 377909
rect 235073 377904 525307 377906
rect 235073 377848 235078 377904
rect 235134 377848 525246 377904
rect 525302 377848 525307 377904
rect 235073 377846 525307 377848
rect 235073 377843 235139 377846
rect 525241 377843 525307 377846
rect 232865 377770 232931 377773
rect 522481 377770 522547 377773
rect 232865 377768 522547 377770
rect 232865 377712 232870 377768
rect 232926 377712 522486 377768
rect 522542 377712 522547 377768
rect 232865 377710 522547 377712
rect 232865 377707 232931 377710
rect 522481 377707 522547 377710
rect 233693 377634 233759 377637
rect 523861 377634 523927 377637
rect 233693 377632 523927 377634
rect 233693 377576 233698 377632
rect 233754 377576 523866 377632
rect 523922 377576 523927 377632
rect 233693 377574 523927 377576
rect 233693 377571 233759 377574
rect 523861 377571 523927 377574
rect 230289 377498 230355 377501
rect 521101 377498 521167 377501
rect 230289 377496 521167 377498
rect 230289 377440 230294 377496
rect 230350 377440 521106 377496
rect 521162 377440 521167 377496
rect 230289 377438 521167 377440
rect 230289 377435 230355 377438
rect 521101 377435 521167 377438
rect 228633 377362 228699 377365
rect 526621 377362 526687 377365
rect 228633 377360 526687 377362
rect 228633 377304 228638 377360
rect 228694 377304 526626 377360
rect 526682 377304 526687 377360
rect 228633 377302 526687 377304
rect 228633 377299 228699 377302
rect 526621 377299 526687 377302
rect 260005 377226 260071 377229
rect 384757 377226 384823 377229
rect 260005 377224 384823 377226
rect 260005 377168 260010 377224
rect 260066 377168 384762 377224
rect 384818 377168 384823 377224
rect 260005 377166 384823 377168
rect 260005 377163 260071 377166
rect 384757 377163 384823 377166
rect 231485 376818 231551 376821
rect 260741 376818 260807 376821
rect 231485 376816 260807 376818
rect 231485 376760 231490 376816
rect 231546 376760 260746 376816
rect 260802 376760 260807 376816
rect 231485 376758 260807 376760
rect 231485 376755 231551 376758
rect 260741 376755 260807 376758
rect 281942 376756 281948 376820
rect 282012 376818 282018 376820
rect 282821 376818 282887 376821
rect 282012 376816 282887 376818
rect 282012 376760 282826 376816
rect 282882 376760 282887 376816
rect 282012 376758 282887 376760
rect 282012 376756 282018 376758
rect 282821 376755 282887 376758
rect 271137 376274 271203 376277
rect 424225 376274 424291 376277
rect 271137 376272 424291 376274
rect 271137 376216 271142 376272
rect 271198 376216 424230 376272
rect 424286 376216 424291 376272
rect 271137 376214 424291 376216
rect 271137 376211 271203 376214
rect 424225 376211 424291 376214
rect 4061 376138 4127 376141
rect 282913 376138 282979 376141
rect 4061 376136 282979 376138
rect 4061 376080 4066 376136
rect 4122 376080 282918 376136
rect 282974 376080 282979 376136
rect 4061 376078 282979 376080
rect 4061 376075 4127 376078
rect 282913 376075 282979 376078
rect 238569 376002 238635 376005
rect 533521 376002 533587 376005
rect 238569 376000 533587 376002
rect 238569 375944 238574 376000
rect 238630 375944 533526 376000
rect 533582 375944 533587 376000
rect 238569 375942 533587 375944
rect 238569 375939 238635 375942
rect 533521 375939 533587 375942
rect 63493 375458 63559 375461
rect 65057 375458 65123 375461
rect 63493 375456 65123 375458
rect 63493 375400 63498 375456
rect 63554 375400 65062 375456
rect 65118 375400 65123 375456
rect 63493 375398 65123 375400
rect 63493 375395 63559 375398
rect 65057 375395 65123 375398
rect 467833 375458 467899 375461
rect 471237 375458 471303 375461
rect 467833 375456 471303 375458
rect 467833 375400 467838 375456
rect 467894 375400 471242 375456
rect 471298 375400 471303 375456
rect 467833 375398 471303 375400
rect 467833 375395 467899 375398
rect 471237 375395 471303 375398
rect 235441 374778 235507 374781
rect 492990 374778 492996 374780
rect 235441 374776 492996 374778
rect 235441 374720 235446 374776
rect 235502 374720 492996 374776
rect 235441 374718 492996 374720
rect 235441 374715 235507 374718
rect 492990 374716 492996 374718
rect 493060 374716 493066 374780
rect 229001 374642 229067 374645
rect 503161 374642 503227 374645
rect 229001 374640 503227 374642
rect 229001 374584 229006 374640
rect 229062 374584 503166 374640
rect 503222 374584 503227 374640
rect 229001 374582 503227 374584
rect 229001 374579 229067 374582
rect 503161 374579 503227 374582
rect 261017 373418 261083 373421
rect 388345 373418 388411 373421
rect 261017 373416 388411 373418
rect 261017 373360 261022 373416
rect 261078 373360 388350 373416
rect 388406 373360 388411 373416
rect 261017 373358 388411 373360
rect 261017 373355 261083 373358
rect 388345 373355 388411 373358
rect 65885 373282 65951 373285
rect 97257 373282 97323 373285
rect 65885 373280 97323 373282
rect 65885 373224 65890 373280
rect 65946 373224 97262 373280
rect 97318 373224 97323 373280
rect 65885 373222 97323 373224
rect 65885 373219 65951 373222
rect 97257 373219 97323 373222
rect 235758 373220 235764 373284
rect 235828 373282 235834 373284
rect 580257 373282 580323 373285
rect 235828 373280 580323 373282
rect 235828 373224 580262 373280
rect 580318 373224 580323 373280
rect 235828 373222 580323 373224
rect 235828 373220 235834 373222
rect 580257 373219 580323 373222
rect 97349 371922 97415 371925
rect 166257 371922 166323 371925
rect 84150 371920 166323 371922
rect 84150 371864 97354 371920
rect 97410 371864 166262 371920
rect 166318 371864 166323 371920
rect 84150 371862 166323 371864
rect -960 371378 480 371468
rect 84150 371378 84210 371862
rect 97349 371859 97415 371862
rect 166257 371859 166323 371862
rect 258993 371922 259059 371925
rect 381169 371922 381235 371925
rect 258993 371920 381235 371922
rect 258993 371864 258998 371920
rect 259054 371864 381174 371920
rect 381230 371864 381235 371920
rect 258993 371862 381235 371864
rect 258993 371859 259059 371862
rect 381169 371859 381235 371862
rect 465073 371514 465139 371517
rect 467097 371514 467163 371517
rect 465073 371512 467163 371514
rect 465073 371456 465078 371512
rect 465134 371456 467102 371512
rect 467158 371456 467163 371512
rect 465073 371454 467163 371456
rect 465073 371451 465139 371454
rect 467097 371451 467163 371454
rect 467833 371378 467899 371381
rect -960 371318 84210 371378
rect 465030 371376 467899 371378
rect 465030 371320 467838 371376
rect 467894 371320 467899 371376
rect 465030 371318 467899 371320
rect -960 371228 480 371318
rect 464337 371242 464403 371245
rect 465030 371242 465090 371318
rect 467833 371315 467899 371318
rect 464337 371240 465090 371242
rect 464337 371184 464342 371240
rect 464398 371184 465090 371240
rect 464337 371182 465090 371184
rect 464337 371179 464403 371182
rect 264237 370698 264303 370701
rect 395521 370698 395587 370701
rect 264237 370696 395587 370698
rect 264237 370640 264242 370696
rect 264298 370640 395526 370696
rect 395582 370640 395587 370696
rect 264237 370638 395587 370640
rect 264237 370635 264303 370638
rect 395521 370635 395587 370638
rect 3366 370500 3372 370564
rect 3436 370562 3442 370564
rect 282862 370562 282868 370564
rect 3436 370502 282868 370562
rect 3436 370500 3442 370502
rect 282862 370500 282868 370502
rect 282932 370500 282938 370564
rect 65057 369746 65123 369749
rect 70301 369746 70367 369749
rect 65057 369744 70367 369746
rect 65057 369688 65062 369744
rect 65118 369688 70306 369744
rect 70362 369688 70367 369744
rect 65057 369686 70367 369688
rect 65057 369683 65123 369686
rect 70301 369683 70367 369686
rect 254945 369338 255011 369341
rect 366817 369338 366883 369341
rect 254945 369336 366883 369338
rect 254945 369280 254950 369336
rect 255006 369280 366822 369336
rect 366878 369280 366883 369336
rect 254945 369278 366883 369280
rect 254945 369275 255011 369278
rect 366817 369275 366883 369278
rect 236821 369202 236887 369205
rect 518341 369202 518407 369205
rect 236821 369200 518407 369202
rect 236821 369144 236826 369200
rect 236882 369144 518346 369200
rect 518402 369144 518407 369200
rect 236821 369142 518407 369144
rect 236821 369139 236887 369142
rect 518341 369139 518407 369142
rect 237925 369066 237991 369069
rect 523677 369066 523743 369069
rect 237925 369064 523743 369066
rect 237925 369008 237930 369064
rect 237986 369008 523682 369064
rect 523738 369008 523743 369064
rect 237925 369006 523743 369008
rect 237925 369003 237991 369006
rect 523677 369003 523743 369006
rect 462957 368386 463023 368389
rect 464981 368386 465047 368389
rect 462957 368384 465047 368386
rect 462957 368328 462962 368384
rect 463018 368328 464986 368384
rect 465042 368328 465047 368384
rect 462957 368326 465047 368328
rect 462957 368323 463023 368326
rect 464981 368323 465047 368326
rect 253933 367706 253999 367709
rect 363229 367706 363295 367709
rect 253933 367704 363295 367706
rect 253933 367648 253938 367704
rect 253994 367648 363234 367704
rect 363290 367648 363295 367704
rect 253933 367646 363295 367648
rect 253933 367643 253999 367646
rect 363229 367643 363295 367646
rect 70393 366346 70459 366349
rect 77937 366346 78003 366349
rect 70393 366344 78003 366346
rect 70393 366288 70398 366344
rect 70454 366288 77942 366344
rect 77998 366288 78003 366344
rect 70393 366286 78003 366288
rect 70393 366283 70459 366286
rect 77937 366283 78003 366286
rect 265065 366346 265131 366349
rect 402697 366346 402763 366349
rect 265065 366344 402763 366346
rect 265065 366288 265070 366344
rect 265126 366288 402702 366344
rect 402758 366288 402763 366344
rect 265065 366286 402763 366288
rect 265065 366283 265131 366286
rect 402697 366283 402763 366286
rect 267089 365122 267155 365125
rect 409873 365122 409939 365125
rect 267089 365120 409939 365122
rect 267089 365064 267094 365120
rect 267150 365064 409878 365120
rect 409934 365064 409939 365120
rect 267089 365062 409939 365064
rect 267089 365059 267155 365062
rect 409873 365059 409939 365062
rect 580390 365060 580396 365124
rect 580460 365122 580466 365124
rect 583520 365122 584960 365212
rect 580460 365062 584960 365122
rect 580460 365060 580466 365062
rect 233877 364986 233943 364989
rect 501781 364986 501847 364989
rect 233877 364984 501847 364986
rect 233877 364928 233882 364984
rect 233938 364928 501786 364984
rect 501842 364928 501847 364984
rect 583520 364972 584960 365062
rect 233877 364926 501847 364928
rect 233877 364923 233943 364926
rect 501781 364923 501847 364926
rect 241789 363762 241855 363765
rect 454677 363762 454743 363765
rect 241789 363760 454743 363762
rect 241789 363704 241794 363760
rect 241850 363704 454682 363760
rect 454738 363704 454743 363760
rect 241789 363702 454743 363704
rect 241789 363699 241855 363702
rect 454677 363699 454743 363702
rect 83457 363626 83523 363629
rect 497457 363626 497523 363629
rect 83457 363624 497523 363626
rect 83457 363568 83462 363624
rect 83518 363568 497462 363624
rect 497518 363568 497523 363624
rect 83457 363566 497523 363568
rect 83457 363563 83523 363566
rect 497457 363563 497523 363566
rect 234245 362538 234311 362541
rect 295057 362538 295123 362541
rect 234245 362536 295123 362538
rect 234245 362480 234250 362536
rect 234306 362480 295062 362536
rect 295118 362480 295123 362536
rect 234245 362478 295123 362480
rect 234245 362475 234311 362478
rect 295057 362475 295123 362478
rect 273897 362402 273963 362405
rect 427813 362402 427879 362405
rect 273897 362400 427879 362402
rect 273897 362344 273902 362400
rect 273958 362344 427818 362400
rect 427874 362344 427879 362400
rect 273897 362342 427879 362344
rect 273897 362339 273963 362342
rect 427813 362339 427879 362342
rect 236729 362266 236795 362269
rect 511441 362266 511507 362269
rect 236729 362264 511507 362266
rect 236729 362208 236734 362264
rect 236790 362208 511446 362264
rect 511502 362208 511507 362264
rect 236729 362206 511507 362208
rect 236729 362203 236795 362206
rect 511441 362203 511507 362206
rect 234337 361042 234403 361045
rect 284293 361042 284359 361045
rect 234337 361040 284359 361042
rect 234337 360984 234342 361040
rect 234398 360984 284298 361040
rect 284354 360984 284359 361040
rect 234337 360982 284359 360984
rect 234337 360979 234403 360982
rect 284293 360979 284359 360982
rect 266997 360906 267063 360909
rect 406285 360906 406351 360909
rect 266997 360904 406351 360906
rect 266997 360848 267002 360904
rect 267058 360848 406290 360904
rect 406346 360848 406351 360904
rect 266997 360846 406351 360848
rect 266997 360843 267063 360846
rect 406285 360843 406351 360846
rect 262857 359546 262923 359549
rect 391933 359546 391999 359549
rect 262857 359544 391999 359546
rect 262857 359488 262862 359544
rect 262918 359488 391938 359544
rect 391994 359488 391999 359544
rect 262857 359486 391999 359488
rect 262857 359483 262923 359486
rect 391933 359483 391999 359486
rect 235349 359410 235415 359413
rect 499021 359410 499087 359413
rect 235349 359408 499087 359410
rect 235349 359352 235354 359408
rect 235410 359352 499026 359408
rect 499082 359352 499087 359408
rect 235349 359350 499087 359352
rect 235349 359347 235415 359350
rect 499021 359347 499087 359350
rect 462957 359002 463023 359005
rect 460890 359000 463023 359002
rect 460890 358944 462962 359000
rect 463018 358944 463023 359000
rect 460890 358942 463023 358944
rect 459553 358730 459619 358733
rect 460890 358730 460950 358942
rect 462957 358939 463023 358942
rect 459553 358728 460950 358730
rect 459553 358672 459558 358728
rect 459614 358672 460950 358728
rect 459553 358670 460950 358672
rect 459553 358667 459619 358670
rect -960 358458 480 358548
rect 294454 358458 294460 358460
rect -960 358398 294460 358458
rect -960 358308 480 358398
rect 294454 358396 294460 358398
rect 294524 358396 294530 358460
rect 246297 358050 246363 358053
rect 327349 358050 327415 358053
rect 246297 358048 327415 358050
rect 246297 357992 246302 358048
rect 246358 357992 327354 358048
rect 327410 357992 327415 358048
rect 246297 357990 327415 357992
rect 246297 357987 246363 357990
rect 327349 357987 327415 357990
rect 462313 357370 462379 357373
rect 464337 357370 464403 357373
rect 462313 357368 464403 357370
rect 462313 357312 462318 357368
rect 462374 357312 464342 357368
rect 464398 357312 464403 357368
rect 462313 357310 464403 357312
rect 462313 357307 462379 357310
rect 464337 357307 464403 357310
rect 234153 356962 234219 356965
rect 309409 356962 309475 356965
rect 234153 356960 309475 356962
rect 234153 356904 234158 356960
rect 234214 356904 309414 356960
rect 309470 356904 309475 356960
rect 234153 356902 309475 356904
rect 234153 356899 234219 356902
rect 309409 356899 309475 356902
rect 274173 356826 274239 356829
rect 434989 356826 435055 356829
rect 274173 356824 435055 356826
rect 274173 356768 274178 356824
rect 274234 356768 434994 356824
rect 435050 356768 435055 356824
rect 274173 356766 435055 356768
rect 274173 356763 274239 356766
rect 434989 356763 435055 356766
rect 235809 356690 235875 356693
rect 580625 356690 580691 356693
rect 235809 356688 580691 356690
rect 235809 356632 235814 356688
rect 235870 356632 580630 356688
rect 580686 356632 580691 356688
rect 235809 356630 580691 356632
rect 235809 356627 235875 356630
rect 580625 356627 580691 356630
rect 458173 356010 458239 356013
rect 459553 356010 459619 356013
rect 458173 356008 459619 356010
rect 458173 355952 458178 356008
rect 458234 355952 459558 356008
rect 459614 355952 459619 356008
rect 458173 355950 459619 355952
rect 458173 355947 458239 355950
rect 459553 355947 459619 355950
rect 239438 355404 239444 355468
rect 239508 355466 239514 355468
rect 320173 355466 320239 355469
rect 239508 355464 320239 355466
rect 239508 355408 320178 355464
rect 320234 355408 320239 355464
rect 239508 355406 320239 355408
rect 239508 355404 239514 355406
rect 320173 355403 320239 355406
rect 237281 355330 237347 355333
rect 474457 355330 474523 355333
rect 237281 355328 474523 355330
rect 237281 355272 237286 355328
rect 237342 355272 474462 355328
rect 474518 355272 474523 355328
rect 237281 355270 474523 355272
rect 237281 355267 237347 355270
rect 474457 355267 474523 355270
rect 235257 354106 235323 354109
rect 496261 354106 496327 354109
rect 235257 354104 496327 354106
rect 235257 354048 235262 354104
rect 235318 354048 496266 354104
rect 496322 354048 496327 354104
rect 235257 354046 496327 354048
rect 235257 354043 235323 354046
rect 496261 354043 496327 354046
rect 237189 353970 237255 353973
rect 580441 353970 580507 353973
rect 237189 353968 580507 353970
rect 237189 353912 237194 353968
rect 237250 353912 580446 353968
rect 580502 353912 580507 353968
rect 237189 353910 580507 353912
rect 237189 353907 237255 353910
rect 580441 353907 580507 353910
rect 233969 352610 234035 352613
rect 312997 352610 313063 352613
rect 233969 352608 313063 352610
rect 233969 352552 233974 352608
rect 234030 352552 313002 352608
rect 313058 352552 313063 352608
rect 233969 352550 313063 352552
rect 233969 352547 234035 352550
rect 312997 352547 313063 352550
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 233785 351386 233851 351389
rect 316585 351386 316651 351389
rect 233785 351384 316651 351386
rect 233785 351328 233790 351384
rect 233846 351328 316590 351384
rect 316646 351328 316651 351384
rect 233785 351326 316651 351328
rect 233785 351323 233851 351326
rect 316585 351323 316651 351326
rect 238477 351250 238543 351253
rect 530761 351250 530827 351253
rect 238477 351248 530827 351250
rect 238477 351192 238482 351248
rect 238538 351192 530766 351248
rect 530822 351192 530827 351248
rect 238477 351190 530827 351192
rect 238477 351187 238543 351190
rect 530761 351187 530827 351190
rect 237005 351114 237071 351117
rect 580533 351114 580599 351117
rect 237005 351112 580599 351114
rect 237005 351056 237010 351112
rect 237066 351056 580538 351112
rect 580594 351056 580599 351112
rect 237005 351054 580599 351056
rect 237005 351051 237071 351054
rect 580533 351051 580599 351054
rect 458909 350434 458975 350437
rect 462313 350434 462379 350437
rect 458909 350432 462379 350434
rect 458909 350376 458914 350432
rect 458970 350376 462318 350432
rect 462374 350376 462379 350432
rect 458909 350374 462379 350376
rect 458909 350371 458975 350374
rect 462313 350371 462379 350374
rect 235165 350026 235231 350029
rect 496854 350026 496860 350028
rect 235165 350024 496860 350026
rect 235165 349968 235170 350024
rect 235226 349968 496860 350024
rect 235165 349966 496860 349968
rect 235165 349963 235231 349966
rect 496854 349964 496860 349966
rect 496924 349964 496930 350028
rect 238518 349828 238524 349892
rect 238588 349890 238594 349892
rect 529197 349890 529263 349893
rect 238588 349888 529263 349890
rect 238588 349832 529202 349888
rect 529258 349832 529263 349888
rect 238588 349830 529263 349832
rect 238588 349828 238594 349830
rect 529197 349827 529263 349830
rect 237230 349692 237236 349756
rect 237300 349754 237306 349756
rect 580206 349754 580212 349756
rect 237300 349694 580212 349754
rect 237300 349692 237306 349694
rect 580206 349692 580212 349694
rect 580276 349692 580282 349756
rect 235901 348530 235967 348533
rect 463693 348530 463759 348533
rect 235901 348528 463759 348530
rect 235901 348472 235906 348528
rect 235962 348472 463698 348528
rect 463754 348472 463759 348528
rect 235901 348470 463759 348472
rect 235901 348467 235967 348470
rect 463693 348467 463759 348470
rect 238334 348332 238340 348396
rect 238404 348394 238410 348396
rect 534901 348394 534967 348397
rect 238404 348392 534967 348394
rect 238404 348336 534906 348392
rect 534962 348336 534967 348392
rect 238404 348334 534967 348336
rect 238404 348332 238410 348334
rect 534901 348331 534967 348334
rect 77937 347714 78003 347717
rect 78857 347714 78923 347717
rect 77937 347712 78923 347714
rect 77937 347656 77942 347712
rect 77998 347656 78862 347712
rect 78918 347656 78923 347712
rect 77937 347654 78923 347656
rect 77937 347651 78003 347654
rect 78857 347651 78923 347654
rect 456793 347714 456859 347717
rect 458909 347714 458975 347717
rect 456793 347712 458975 347714
rect 456793 347656 456798 347712
rect 456854 347656 458914 347712
rect 458970 347656 458975 347712
rect 456793 347654 458975 347656
rect 456793 347651 456859 347654
rect 458909 347651 458975 347654
rect 239254 347108 239260 347172
rect 239324 347170 239330 347172
rect 536281 347170 536347 347173
rect 239324 347168 536347 347170
rect 239324 347112 536286 347168
rect 536342 347112 536347 347168
rect 239324 347110 536347 347112
rect 239324 347108 239330 347110
rect 536281 347107 536347 347110
rect 69013 347034 69079 347037
rect 507945 347034 508011 347037
rect 69013 347032 508011 347034
rect 69013 346976 69018 347032
rect 69074 346976 507950 347032
rect 508006 346976 508011 347032
rect 69013 346974 508011 346976
rect 69013 346971 69079 346974
rect 507945 346971 508011 346974
rect 239581 346082 239647 346085
rect 273529 346082 273595 346085
rect 239581 346080 273595 346082
rect 239581 346024 239586 346080
rect 239642 346024 273534 346080
rect 273590 346024 273595 346080
rect 239581 346022 273595 346024
rect 239581 346019 239647 346022
rect 273529 346019 273595 346022
rect 238017 345946 238083 345949
rect 302233 345946 302299 345949
rect 238017 345944 302299 345946
rect 238017 345888 238022 345944
rect 238078 345888 302238 345944
rect 302294 345888 302299 345944
rect 238017 345886 302299 345888
rect 238017 345883 238083 345886
rect 302233 345883 302299 345886
rect 238150 345748 238156 345812
rect 238220 345810 238226 345812
rect 494094 345810 494100 345812
rect 238220 345750 494100 345810
rect 238220 345748 238226 345750
rect 494094 345748 494100 345750
rect 494164 345748 494170 345812
rect 236545 345674 236611 345677
rect 504541 345674 504607 345677
rect 236545 345672 504607 345674
rect 236545 345616 236550 345672
rect 236606 345616 504546 345672
rect 504602 345616 504607 345672
rect 236545 345614 504607 345616
rect 236545 345611 236611 345614
rect 504541 345611 504607 345614
rect -960 345402 480 345492
rect 230974 345402 230980 345404
rect -960 345342 230980 345402
rect -960 345252 480 345342
rect 230974 345340 230980 345342
rect 231044 345340 231050 345404
rect 242709 344994 242775 344997
rect 323761 344994 323827 344997
rect 242709 344992 323827 344994
rect 242709 344936 242714 344992
rect 242770 344936 323766 344992
rect 323822 344936 323827 344992
rect 242709 344934 323827 344936
rect 242709 344931 242775 344934
rect 323761 344931 323827 344934
rect 252921 344858 252987 344861
rect 359641 344858 359707 344861
rect 252921 344856 359707 344858
rect 252921 344800 252926 344856
rect 252982 344800 359646 344856
rect 359702 344800 359707 344856
rect 252921 344798 359707 344800
rect 252921 344795 252987 344798
rect 359641 344795 359707 344798
rect 78857 344722 78923 344725
rect 86861 344722 86927 344725
rect 78857 344720 86927 344722
rect 78857 344664 78862 344720
rect 78918 344664 86866 344720
rect 86922 344664 86927 344720
rect 78857 344662 86927 344664
rect 78857 344659 78923 344662
rect 86861 344659 86927 344662
rect 255957 344722 256023 344725
rect 370405 344722 370471 344725
rect 255957 344720 370471 344722
rect 255957 344664 255962 344720
rect 256018 344664 370410 344720
rect 370466 344664 370471 344720
rect 255957 344662 370471 344664
rect 255957 344659 256023 344662
rect 370405 344659 370471 344662
rect 48078 344524 48084 344588
rect 48148 344586 48154 344588
rect 253197 344586 253263 344589
rect 48148 344584 253263 344586
rect 48148 344528 253202 344584
rect 253258 344528 253263 344584
rect 48148 344526 253263 344528
rect 48148 344524 48154 344526
rect 253197 344523 253263 344526
rect 256969 344586 257035 344589
rect 373993 344586 374059 344589
rect 256969 344584 374059 344586
rect 256969 344528 256974 344584
rect 257030 344528 373998 344584
rect 374054 344528 374059 344584
rect 256969 344526 374059 344528
rect 256969 344523 257035 344526
rect 373993 344523 374059 344526
rect 231158 344388 231164 344452
rect 231228 344450 231234 344452
rect 256693 344450 256759 344453
rect 231228 344448 256759 344450
rect 231228 344392 256698 344448
rect 256754 344392 256759 344448
rect 231228 344390 256759 344392
rect 231228 344388 231234 344390
rect 256693 344387 256759 344390
rect 264053 344450 264119 344453
rect 399109 344450 399175 344453
rect 264053 344448 399175 344450
rect 264053 344392 264058 344448
rect 264114 344392 399114 344448
rect 399170 344392 399175 344448
rect 264053 344390 399175 344392
rect 264053 344387 264119 344390
rect 399109 344387 399175 344390
rect 239489 344314 239555 344317
rect 266353 344314 266419 344317
rect 239489 344312 266419 344314
rect 239489 344256 239494 344312
rect 239550 344256 266358 344312
rect 266414 344256 266419 344312
rect 239489 344254 266419 344256
rect 239489 344251 239555 344254
rect 266353 344251 266419 344254
rect 268101 344314 268167 344317
rect 413461 344314 413527 344317
rect 268101 344312 413527 344314
rect 268101 344256 268106 344312
rect 268162 344256 413466 344312
rect 413522 344256 413527 344312
rect 268101 344254 413527 344256
rect 268101 344251 268167 344254
rect 413461 344251 413527 344254
rect 224350 344116 224356 344180
rect 224420 344178 224426 344180
rect 255313 344178 255379 344181
rect 224420 344176 255379 344178
rect 224420 344120 255318 344176
rect 255374 344120 255379 344176
rect 224420 344118 255379 344120
rect 224420 344116 224426 344118
rect 255313 344115 255379 344118
rect 230054 343980 230060 344044
rect 230124 344042 230130 344044
rect 263593 344042 263659 344045
rect 230124 344040 263659 344042
rect 230124 343984 263598 344040
rect 263654 343984 263659 344040
rect 230124 343982 263659 343984
rect 230124 343980 230130 343982
rect 263593 343979 263659 343982
rect 229870 343844 229876 343908
rect 229940 343906 229946 343908
rect 285990 343906 285996 343908
rect 229940 343846 285996 343906
rect 229940 343844 229946 343846
rect 285990 343844 285996 343846
rect 286060 343844 286066 343908
rect 235625 343770 235691 343773
rect 242801 343770 242867 343773
rect 235625 343768 242867 343770
rect 235625 343712 235630 343768
rect 235686 343712 242806 343768
rect 242862 343712 242867 343768
rect 235625 343710 242867 343712
rect 235625 343707 235691 343710
rect 242801 343707 242867 343710
rect 227478 343572 227484 343636
rect 227548 343634 227554 343636
rect 247033 343634 247099 343637
rect 227548 343632 247099 343634
rect 227548 343576 247038 343632
rect 247094 343576 247099 343632
rect 227548 343574 247099 343576
rect 227548 343572 227554 343574
rect 247033 343571 247099 343574
rect 224902 343436 224908 343500
rect 224972 343498 224978 343500
rect 251081 343498 251147 343501
rect 224972 343496 251147 343498
rect 224972 343440 251086 343496
rect 251142 343440 251147 343496
rect 224972 343438 251147 343440
rect 224972 343436 224978 343438
rect 251081 343435 251147 343438
rect 250897 343362 250963 343365
rect 352465 343362 352531 343365
rect 250897 343360 352531 343362
rect 250897 343304 250902 343360
rect 250958 343304 352470 343360
rect 352526 343304 352531 343360
rect 250897 343302 352531 343304
rect 250897 343299 250963 343302
rect 352465 343299 352531 343302
rect 245837 343226 245903 343229
rect 258717 343226 258783 343229
rect 245837 343224 258783 343226
rect 245837 343168 245842 343224
rect 245898 343168 258722 343224
rect 258778 343168 258783 343224
rect 245837 343166 258783 343168
rect 245837 343163 245903 343166
rect 258717 343163 258783 343166
rect 276197 343226 276263 343229
rect 392577 343226 392643 343229
rect 276197 343224 392643 343226
rect 276197 343168 276202 343224
rect 276258 343168 392582 343224
rect 392638 343168 392643 343224
rect 276197 343166 392643 343168
rect 276197 343163 276263 343166
rect 392577 343163 392643 343166
rect 227110 343028 227116 343092
rect 227180 343090 227186 343092
rect 245653 343090 245719 343093
rect 227180 343088 245719 343090
rect 227180 343032 245658 343088
rect 245714 343032 245719 343088
rect 227180 343030 245719 343032
rect 227180 343028 227186 343030
rect 245653 343027 245719 343030
rect 247861 343090 247927 343093
rect 256049 343090 256115 343093
rect 247861 343088 256115 343090
rect 247861 343032 247866 343088
rect 247922 343032 256054 343088
rect 256110 343032 256115 343088
rect 247861 343030 256115 343032
rect 247861 343027 247927 343030
rect 256049 343027 256115 343030
rect 278221 343090 278287 343093
rect 417417 343090 417483 343093
rect 278221 343088 417483 343090
rect 278221 343032 278226 343088
rect 278282 343032 417422 343088
rect 417478 343032 417483 343088
rect 278221 343030 417483 343032
rect 278221 343027 278287 343030
rect 417417 343027 417483 343030
rect 239397 342954 239463 342957
rect 269941 342954 270007 342957
rect 239397 342952 270007 342954
rect 239397 342896 239402 342952
rect 239458 342896 269946 342952
rect 270002 342896 270007 342952
rect 239397 342894 270007 342896
rect 239397 342891 239463 342894
rect 269941 342891 270007 342894
rect 279233 342954 279299 342957
rect 482461 342954 482527 342957
rect 279233 342952 482527 342954
rect 279233 342896 279238 342952
rect 279294 342896 482466 342952
rect 482522 342896 482527 342952
rect 279233 342894 482527 342896
rect 279233 342891 279299 342894
rect 482461 342891 482527 342894
rect 244825 342818 244891 342821
rect 330937 342818 331003 342821
rect 244825 342816 331003 342818
rect 244825 342760 244830 342816
rect 244886 342760 330942 342816
rect 330998 342760 331003 342816
rect 244825 342758 331003 342760
rect 244825 342755 244891 342758
rect 330937 342755 331003 342758
rect 223246 342620 223252 342684
rect 223316 342682 223322 342684
rect 243537 342682 243603 342685
rect 223316 342680 243603 342682
rect 223316 342624 243542 342680
rect 243598 342624 243603 342680
rect 223316 342622 243603 342624
rect 223316 342620 223322 342622
rect 243537 342619 243603 342622
rect 248873 342682 248939 342685
rect 345289 342682 345355 342685
rect 248873 342680 345355 342682
rect 248873 342624 248878 342680
rect 248934 342624 345294 342680
rect 345350 342624 345355 342680
rect 248873 342622 345355 342624
rect 248873 342619 248939 342622
rect 345289 342619 345355 342622
rect 224534 342484 224540 342548
rect 224604 342546 224610 342548
rect 244273 342546 244339 342549
rect 224604 342544 244339 342546
rect 224604 342488 244278 342544
rect 244334 342488 244339 342544
rect 224604 342486 244339 342488
rect 224604 342484 224610 342486
rect 244273 342483 244339 342486
rect 246849 342546 246915 342549
rect 338113 342546 338179 342549
rect 246849 342544 338179 342546
rect 246849 342488 246854 342544
rect 246910 342488 338118 342544
rect 338174 342488 338179 342544
rect 246849 342486 338179 342488
rect 246849 342483 246915 342486
rect 338113 342483 338179 342486
rect 222929 342410 222995 342413
rect 226333 342410 226399 342413
rect 222929 342408 226399 342410
rect 222929 342352 222934 342408
rect 222990 342352 226338 342408
rect 226394 342352 226399 342408
rect 222929 342350 226399 342352
rect 222929 342347 222995 342350
rect 226333 342347 226399 342350
rect 227294 342348 227300 342412
rect 227364 342410 227370 342412
rect 249701 342410 249767 342413
rect 227364 342408 249767 342410
rect 227364 342352 249706 342408
rect 249762 342352 249767 342408
rect 227364 342350 249767 342352
rect 227364 342348 227370 342350
rect 249701 342347 249767 342350
rect 224166 342212 224172 342276
rect 224236 342274 224242 342276
rect 226609 342274 226675 342277
rect 224236 342272 226675 342274
rect 224236 342216 226614 342272
rect 226670 342216 226675 342272
rect 224236 342214 226675 342216
rect 224236 342212 224242 342214
rect 226609 342211 226675 342214
rect 227621 342274 227687 342277
rect 240041 342274 240107 342277
rect 227621 342272 240107 342274
rect 227621 342216 227626 342272
rect 227682 342216 240046 342272
rect 240102 342216 240107 342272
rect 227621 342214 240107 342216
rect 227621 342211 227687 342214
rect 240041 342211 240107 342214
rect 243813 342274 243879 342277
rect 246297 342274 246363 342277
rect 243813 342272 246363 342274
rect 243813 342216 243818 342272
rect 243874 342216 246302 342272
rect 246358 342216 246363 342272
rect 243813 342214 246363 342216
rect 243813 342211 243879 342214
rect 246297 342211 246363 342214
rect 262029 342274 262095 342277
rect 262857 342274 262923 342277
rect 262029 342272 262923 342274
rect 262029 342216 262034 342272
rect 262090 342216 262862 342272
rect 262918 342216 262923 342272
rect 262029 342214 262923 342216
rect 262029 342211 262095 342214
rect 262857 342211 262923 342214
rect 263041 342274 263107 342277
rect 264237 342274 264303 342277
rect 263041 342272 264303 342274
rect 263041 342216 263046 342272
rect 263102 342216 264242 342272
rect 264298 342216 264303 342272
rect 263041 342214 264303 342216
rect 263041 342211 263107 342214
rect 264237 342211 264303 342214
rect 269113 342274 269179 342277
rect 271229 342274 271295 342277
rect 269113 342272 271295 342274
rect 269113 342216 269118 342272
rect 269174 342216 271234 342272
rect 271290 342216 271295 342272
rect 269113 342214 271295 342216
rect 269113 342211 269179 342214
rect 271229 342211 271295 342214
rect 272149 342274 272215 342277
rect 273897 342274 273963 342277
rect 272149 342272 273963 342274
rect 272149 342216 272154 342272
rect 272210 342216 273902 342272
rect 273958 342216 273963 342272
rect 272149 342214 273963 342216
rect 272149 342211 272215 342214
rect 273897 342211 273963 342214
rect 29494 342076 29500 342140
rect 29564 342138 29570 342140
rect 227713 342138 227779 342141
rect 29564 342136 227779 342138
rect 29564 342080 227718 342136
rect 227774 342080 227779 342136
rect 29564 342078 227779 342080
rect 29564 342076 29570 342078
rect 227713 342075 227779 342078
rect 86861 342002 86927 342005
rect 90357 342002 90423 342005
rect 86861 342000 90423 342002
rect 86861 341944 86866 342000
rect 86922 341944 90362 342000
rect 90418 341944 90423 342000
rect 86861 341942 90423 341944
rect 86861 341939 86927 341942
rect 90357 341939 90423 341942
rect 222878 341940 222884 342004
rect 222948 342002 222954 342004
rect 285622 342002 285628 342004
rect 222948 341942 285628 342002
rect 222948 341940 222954 341942
rect 285622 341940 285628 341942
rect 285692 341940 285698 342004
rect 32397 341866 32463 341869
rect 225045 341866 225111 341869
rect 32397 341864 225111 341866
rect 32397 341808 32402 341864
rect 32458 341808 225050 341864
rect 225106 341808 225111 341864
rect 32397 341806 225111 341808
rect 32397 341803 32463 341806
rect 225045 341803 225111 341806
rect 226190 341804 226196 341868
rect 226260 341866 226266 341868
rect 284518 341866 284524 341868
rect 226260 341806 284524 341866
rect 226260 341804 226266 341806
rect 284518 341804 284524 341806
rect 284588 341804 284594 341868
rect 33041 341730 33107 341733
rect 225137 341730 225203 341733
rect 33041 341728 225203 341730
rect 33041 341672 33046 341728
rect 33102 341672 225142 341728
rect 225198 341672 225203 341728
rect 33041 341670 225203 341672
rect 33041 341667 33107 341670
rect 225137 341667 225203 341670
rect 239121 341730 239187 341733
rect 255589 341730 255655 341733
rect 239121 341728 255655 341730
rect 239121 341672 239126 341728
rect 239182 341672 255594 341728
rect 255650 341672 255655 341728
rect 239121 341670 255655 341672
rect 239121 341667 239187 341670
rect 255589 341667 255655 341670
rect 30281 341594 30347 341597
rect 224953 341594 225019 341597
rect 30281 341592 225019 341594
rect 30281 341536 30286 341592
rect 30342 341536 224958 341592
rect 225014 341536 225019 341592
rect 30281 341534 225019 341536
rect 30281 341531 30347 341534
rect 224953 341531 225019 341534
rect 238201 341594 238267 341597
rect 280705 341594 280771 341597
rect 238201 341592 280771 341594
rect 238201 341536 238206 341592
rect 238262 341536 280710 341592
rect 280766 341536 280771 341592
rect 238201 341534 280771 341536
rect 238201 341531 238267 341534
rect 280705 341531 280771 341534
rect 225781 341458 225847 341461
rect 237373 341458 237439 341461
rect 225781 341456 237439 341458
rect 225781 341400 225786 341456
rect 225842 341400 237378 341456
rect 237434 341400 237439 341456
rect 225781 341398 237439 341400
rect 225781 341395 225847 341398
rect 237373 341395 237439 341398
rect 237741 341458 237807 341461
rect 277117 341458 277183 341461
rect 237741 341456 277183 341458
rect 237741 341400 237746 341456
rect 237802 341400 277122 341456
rect 277178 341400 277183 341456
rect 237741 341398 277183 341400
rect 237741 341395 237807 341398
rect 277117 341395 277183 341398
rect 223062 341260 223068 341324
rect 223132 341322 223138 341324
rect 251030 341322 251036 341324
rect 223132 341262 251036 341322
rect 223132 341260 223138 341262
rect 251030 341260 251036 341262
rect 251100 341260 251106 341324
rect 225965 341186 226031 341189
rect 280889 341186 280955 341189
rect 225965 341184 280955 341186
rect 225965 341128 225970 341184
rect 226026 341128 280894 341184
rect 280950 341128 280955 341184
rect 225965 341126 280955 341128
rect 225965 341123 226031 341126
rect 280889 341123 280955 341126
rect 228357 341050 228423 341053
rect 237465 341050 237531 341053
rect 228357 341048 237531 341050
rect 228357 340992 228362 341048
rect 228418 340992 237470 341048
rect 237526 340992 237531 341048
rect 228357 340990 237531 340992
rect 228357 340987 228423 340990
rect 237465 340987 237531 340990
rect 223205 340914 223271 340917
rect 227805 340914 227871 340917
rect 223205 340912 227871 340914
rect 223205 340856 223210 340912
rect 223266 340856 227810 340912
rect 227866 340856 227871 340912
rect 223205 340854 227871 340856
rect 223205 340851 223271 340854
rect 227805 340851 227871 340854
rect 228173 340914 228239 340917
rect 240041 340914 240107 340917
rect 228173 340912 240107 340914
rect 228173 340856 228178 340912
rect 228234 340856 240046 340912
rect 240102 340856 240107 340912
rect 228173 340854 240107 340856
rect 228173 340851 228239 340854
rect 240041 340851 240107 340854
rect 226149 340778 226215 340781
rect 239949 340778 240015 340781
rect 226149 340776 240015 340778
rect 226149 340720 226154 340776
rect 226210 340720 239954 340776
rect 240010 340720 240015 340776
rect 226149 340718 240015 340720
rect 226149 340715 226215 340718
rect 239949 340715 240015 340718
rect 239305 340642 239371 340645
rect 262765 340642 262831 340645
rect 239305 340640 262831 340642
rect 239305 340584 239310 340640
rect 239366 340584 262770 340640
rect 262826 340584 262831 340640
rect 239305 340582 262831 340584
rect 239305 340579 239371 340582
rect 262765 340579 262831 340582
rect 239673 340506 239739 340509
rect 248505 340506 248571 340509
rect 239673 340504 248571 340506
rect 239673 340448 239678 340504
rect 239734 340448 248510 340504
rect 248566 340448 248571 340504
rect 239673 340446 248571 340448
rect 239673 340443 239739 340446
rect 248505 340443 248571 340446
rect 251030 340444 251036 340508
rect 251100 340506 251106 340508
rect 285806 340506 285812 340508
rect 251100 340446 285812 340506
rect 251100 340444 251106 340446
rect 285806 340444 285812 340446
rect 285876 340444 285882 340508
rect 228541 340370 228607 340373
rect 237465 340370 237531 340373
rect 228541 340368 237531 340370
rect 228541 340312 228546 340368
rect 228602 340312 237470 340368
rect 237526 340312 237531 340368
rect 228541 340310 237531 340312
rect 228541 340307 228607 340310
rect 237465 340307 237531 340310
rect 238201 340370 238267 340373
rect 287881 340370 287947 340373
rect 238201 340368 287947 340370
rect 238201 340312 238206 340368
rect 238262 340312 287886 340368
rect 287942 340312 287947 340368
rect 238201 340310 287947 340312
rect 238201 340307 238267 340310
rect 287881 340307 287947 340310
rect 238109 340234 238175 340237
rect 291469 340234 291535 340237
rect 238109 340232 291535 340234
rect 238109 340176 238114 340232
rect 238170 340176 291474 340232
rect 291530 340176 291535 340232
rect 238109 340174 291535 340176
rect 238109 340171 238175 340174
rect 291469 340171 291535 340174
rect 225597 340098 225663 340101
rect 237373 340098 237439 340101
rect 225597 340096 237439 340098
rect 225597 340040 225602 340096
rect 225658 340040 237378 340096
rect 237434 340040 237439 340096
rect 225597 340038 237439 340040
rect 225597 340035 225663 340038
rect 237373 340035 237439 340038
rect 237833 340098 237899 340101
rect 298645 340098 298711 340101
rect 237833 340096 298711 340098
rect 237833 340040 237838 340096
rect 237894 340040 298650 340096
rect 298706 340040 298711 340096
rect 237833 340038 298711 340040
rect 237833 340035 237899 340038
rect 298645 340035 298711 340038
rect 226926 339900 226932 339964
rect 226996 339962 227002 339964
rect 240041 339962 240107 339965
rect 252185 339962 252251 339965
rect 226996 339960 240107 339962
rect 226996 339904 240046 339960
rect 240102 339904 240107 339960
rect 226996 339902 240107 339904
rect 226996 339900 227002 339902
rect 240041 339899 240107 339902
rect 248370 339960 252251 339962
rect 248370 339904 252190 339960
rect 252246 339904 252251 339960
rect 248370 339902 252251 339904
rect 225413 339826 225479 339829
rect 239857 339826 239923 339829
rect 225413 339824 239923 339826
rect 225413 339768 225418 339824
rect 225474 339768 239862 339824
rect 239918 339768 239923 339824
rect 225413 339766 239923 339768
rect 225413 339763 225479 339766
rect 239857 339763 239923 339766
rect 240041 339826 240107 339829
rect 248370 339826 248430 339902
rect 252185 339899 252251 339902
rect 240041 339824 248430 339826
rect 240041 339768 240046 339824
rect 240102 339768 248430 339824
rect 240041 339766 248430 339768
rect 240041 339763 240107 339766
rect 228265 339690 228331 339693
rect 237557 339690 237623 339693
rect 228265 339688 237623 339690
rect 228265 339632 228270 339688
rect 228326 339632 237562 339688
rect 237618 339632 237623 339688
rect 228265 339630 237623 339632
rect 228265 339627 228331 339630
rect 237557 339627 237623 339630
rect 222694 339492 222700 339556
rect 222764 339554 222770 339556
rect 287094 339554 287100 339556
rect 222764 339494 287100 339554
rect 222764 339492 222770 339494
rect 287094 339492 287100 339494
rect 287164 339492 287170 339556
rect 238661 339418 238727 339421
rect 241237 339418 241303 339421
rect 238661 339416 241303 339418
rect 238661 339360 238666 339416
rect 238722 339360 241242 339416
rect 241298 339360 241303 339416
rect 238661 339358 241303 339360
rect 238661 339355 238727 339358
rect 241237 339355 241303 339358
rect 453297 339418 453363 339421
rect 456793 339418 456859 339421
rect 453297 339416 456859 339418
rect 453297 339360 453302 339416
rect 453358 339360 456798 339416
rect 456854 339360 456859 339416
rect 453297 339358 456859 339360
rect 453297 339355 453363 339358
rect 456793 339355 456859 339358
rect 231025 338874 231091 338877
rect 280654 338874 280660 338876
rect 231025 338872 280660 338874
rect 231025 338816 231030 338872
rect 231086 338816 280660 338872
rect 231025 338814 280660 338816
rect 231025 338811 231091 338814
rect 280654 338812 280660 338814
rect 280724 338812 280730 338876
rect 282361 338874 282427 338877
rect 539777 338874 539843 338877
rect 282361 338872 539843 338874
rect 282361 338816 282366 338872
rect 282422 338816 539782 338872
rect 539838 338816 539843 338872
rect 282361 338814 539843 338816
rect 282361 338811 282427 338814
rect 539777 338811 539843 338814
rect 65425 338738 65491 338741
rect 490046 338738 490052 338740
rect 65425 338736 490052 338738
rect 65425 338680 65430 338736
rect 65486 338680 490052 338736
rect 65425 338678 490052 338680
rect 65425 338675 65491 338678
rect 490046 338676 490052 338678
rect 490116 338676 490122 338740
rect 230933 338602 230999 338605
rect 280521 338602 280587 338605
rect 230933 338600 280587 338602
rect 230933 338544 230938 338600
rect 230994 338544 280526 338600
rect 280582 338544 280587 338600
rect 230933 338542 280587 338544
rect 230933 338539 230999 338542
rect 280521 338539 280587 338542
rect 227529 338466 227595 338469
rect 280153 338466 280219 338469
rect 227529 338464 280219 338466
rect 227529 338408 227534 338464
rect 227590 338408 280158 338464
rect 280214 338408 280219 338464
rect 583520 338452 584960 338692
rect 227529 338406 280219 338408
rect 227529 338403 227595 338406
rect 280153 338403 280219 338406
rect 228214 338268 228220 338332
rect 228284 338330 228290 338332
rect 284702 338330 284708 338332
rect 228284 338270 284708 338330
rect 228284 338268 228290 338270
rect 284702 338268 284708 338270
rect 284772 338268 284778 338332
rect 228398 338132 228404 338196
rect 228468 338194 228474 338196
rect 290590 338194 290596 338196
rect 228468 338134 290596 338194
rect 228468 338132 228474 338134
rect 290590 338132 290596 338134
rect 290660 338132 290666 338196
rect 233734 337588 233740 337652
rect 233804 337650 233810 337652
rect 281574 337650 281580 337652
rect 233804 337590 281580 337650
rect 233804 337588 233810 337590
rect 281574 337588 281580 337590
rect 281644 337588 281650 337652
rect 238385 337514 238451 337517
rect 238385 337512 239690 337514
rect 238385 337456 238390 337512
rect 238446 337456 239690 337512
rect 238385 337454 239690 337456
rect 238385 337451 238451 337454
rect 239630 337310 239690 337454
rect 295926 337316 295932 337380
rect 295996 337378 296002 337380
rect 580390 337378 580396 337380
rect 295996 337318 580396 337378
rect 295996 337316 296002 337318
rect 580390 337316 580396 337318
rect 580460 337316 580466 337380
rect 239630 337250 240212 337310
rect 238518 336228 238524 336292
rect 238588 336290 238594 336292
rect 238588 336230 239690 336290
rect 238588 336228 238594 336230
rect 239630 336222 239690 336230
rect 239630 336162 240212 336222
rect 287646 335956 287652 336020
rect 287716 336018 287722 336020
rect 542670 336018 542676 336020
rect 287716 335958 542676 336018
rect 287716 335956 287722 335958
rect 542670 335956 542676 335958
rect 542740 335956 542746 336020
rect 239254 335140 239260 335204
rect 239324 335202 239330 335204
rect 239324 335142 239690 335202
rect 239324 335140 239330 335142
rect 239630 335134 239690 335142
rect 239630 335074 240212 335134
rect 239814 333986 240212 334046
rect 238334 333916 238340 333980
rect 238404 333978 238410 333980
rect 239814 333978 239874 333986
rect 238404 333918 239874 333978
rect 238404 333916 238410 333918
rect 237649 333298 237715 333301
rect 239029 333298 239095 333301
rect 237649 333296 239095 333298
rect 237649 333240 237654 333296
rect 237710 333240 239034 333296
rect 239090 333240 239095 333296
rect 237649 333238 239095 333240
rect 237649 333235 237715 333238
rect 239029 333235 239095 333238
rect 298686 333236 298692 333300
rect 298756 333298 298762 333300
rect 543590 333298 543596 333300
rect 298756 333238 543596 333298
rect 298756 333236 298762 333238
rect 543590 333236 543596 333238
rect 543660 333236 543666 333300
rect 238569 333026 238635 333029
rect 238569 333024 239690 333026
rect 238569 332968 238574 333024
rect 238630 332968 239690 333024
rect 238569 332966 239690 332968
rect 238569 332963 238635 332966
rect 239630 332958 239690 332966
rect 239630 332898 240212 332958
rect 90357 332618 90423 332621
rect 91737 332618 91803 332621
rect 90357 332616 91803 332618
rect 90357 332560 90362 332616
rect 90418 332560 91742 332616
rect 91798 332560 91803 332616
rect 90357 332558 91803 332560
rect 90357 332555 90423 332558
rect 91737 332555 91803 332558
rect 447777 332482 447843 332485
rect 453297 332482 453363 332485
rect 447777 332480 453363 332482
rect -960 332196 480 332436
rect 447777 332424 447782 332480
rect 447838 332424 453302 332480
rect 453358 332424 453363 332480
rect 447777 332422 453363 332424
rect 447777 332419 447843 332422
rect 453297 332419 453363 332422
rect 237925 331938 237991 331941
rect 237925 331936 239690 331938
rect 237925 331880 237930 331936
rect 237986 331880 239690 331936
rect 237925 331878 239690 331880
rect 237925 331875 237991 331878
rect 239630 331870 239690 331878
rect 239630 331810 240212 331870
rect 282453 331802 282519 331805
rect 539593 331802 539659 331805
rect 282453 331800 539659 331802
rect 282453 331744 282458 331800
rect 282514 331744 539598 331800
rect 539654 331744 539659 331800
rect 282453 331742 539659 331744
rect 282453 331739 282519 331742
rect 539593 331739 539659 331742
rect 237925 331122 237991 331125
rect 239213 331122 239279 331125
rect 237925 331120 239279 331122
rect 237925 331064 237930 331120
rect 237986 331064 239218 331120
rect 239274 331064 239279 331120
rect 237925 331062 239279 331064
rect 237925 331059 237991 331062
rect 239213 331059 239279 331062
rect 238477 330850 238543 330853
rect 238477 330848 239690 330850
rect 238477 330792 238482 330848
rect 238538 330792 239690 330848
rect 238477 330790 239690 330792
rect 238477 330787 238543 330790
rect 239630 330782 239690 330790
rect 239630 330722 240212 330782
rect 282545 330442 282611 330445
rect 539685 330442 539751 330445
rect 282545 330440 539751 330442
rect 282545 330384 282550 330440
rect 282606 330384 539690 330440
rect 539746 330384 539751 330440
rect 282545 330382 539751 330384
rect 282545 330379 282611 330382
rect 539685 330379 539751 330382
rect 236453 329762 236519 329765
rect 238017 329762 238083 329765
rect 236453 329760 238083 329762
rect 236453 329704 236458 329760
rect 236514 329704 238022 329760
rect 238078 329704 238083 329760
rect 236453 329702 238083 329704
rect 236453 329699 236519 329702
rect 238017 329699 238083 329702
rect 239630 329634 240212 329694
rect 231485 329626 231551 329629
rect 239630 329626 239690 329634
rect 231485 329624 239690 329626
rect 231485 329568 231490 329624
rect 231546 329568 239690 329624
rect 231485 329566 239690 329568
rect 231485 329563 231551 329566
rect 536046 328810 536052 328812
rect 230197 328674 230263 328677
rect 279926 328674 279986 328780
rect 287010 328750 536052 328810
rect 287010 328674 287070 328750
rect 536046 328748 536052 328750
rect 536116 328748 536122 328812
rect 230197 328672 239690 328674
rect 230197 328616 230202 328672
rect 230258 328616 239690 328672
rect 230197 328614 239690 328616
rect 279926 328614 287070 328674
rect 230197 328611 230263 328614
rect 239630 328606 239690 328614
rect 239630 328546 240212 328606
rect 538438 327994 538444 327996
rect 279926 327858 279986 327964
rect 287010 327934 538444 327994
rect 287010 327858 287070 327934
rect 538438 327932 538444 327934
rect 538508 327932 538514 327996
rect 279926 327798 287070 327858
rect 228633 327586 228699 327589
rect 228633 327584 239690 327586
rect 228633 327528 228638 327584
rect 228694 327528 239690 327584
rect 228633 327526 239690 327528
rect 228633 327523 228699 327526
rect 239630 327518 239690 327526
rect 239630 327458 240212 327518
rect 279926 327254 287070 327314
rect 279926 327148 279986 327254
rect 287010 327178 287070 327254
rect 530526 327178 530532 327180
rect 287010 327118 530532 327178
rect 530526 327116 530532 327118
rect 530596 327116 530602 327180
rect 456057 327042 456123 327045
rect 457437 327042 457503 327045
rect 456057 327040 457503 327042
rect 456057 326984 456062 327040
rect 456118 326984 457442 327040
rect 457498 326984 457503 327040
rect 456057 326982 457503 326984
rect 456057 326979 456123 326982
rect 457437 326979 457503 326982
rect 235073 326498 235139 326501
rect 235073 326496 239690 326498
rect 235073 326440 235078 326496
rect 235134 326440 239690 326496
rect 235073 326438 239690 326440
rect 235073 326435 235139 326438
rect 239630 326430 239690 326438
rect 239630 326370 240212 326430
rect 533286 326362 533292 326364
rect 279926 326226 279986 326332
rect 287010 326302 533292 326362
rect 287010 326226 287070 326302
rect 533286 326300 533292 326302
rect 533356 326300 533362 326364
rect 279926 326166 287070 326226
rect 501454 325546 501460 325548
rect 233693 325410 233759 325413
rect 279926 325410 279986 325516
rect 287010 325486 501460 325546
rect 287010 325410 287070 325486
rect 501454 325484 501460 325486
rect 501524 325484 501530 325548
rect 233693 325408 239690 325410
rect 233693 325352 233698 325408
rect 233754 325352 239690 325408
rect 233693 325350 239690 325352
rect 279926 325350 287070 325410
rect 233693 325347 233759 325350
rect 239630 325342 239690 325350
rect 239630 325282 240212 325342
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect 538254 324730 538260 324732
rect 279926 324594 279986 324700
rect 287010 324670 538260 324730
rect 287010 324594 287070 324670
rect 538254 324668 538260 324670
rect 538324 324668 538330 324732
rect 279926 324534 287070 324594
rect 232865 324322 232931 324325
rect 232865 324320 239690 324322
rect 232865 324264 232870 324320
rect 232926 324264 239690 324320
rect 232865 324262 239690 324264
rect 232865 324259 232931 324262
rect 239630 324254 239690 324262
rect 239630 324194 240212 324254
rect 511206 323914 511212 323916
rect 279926 323778 279986 323884
rect 287010 323854 511212 323914
rect 287010 323778 287070 323854
rect 511206 323852 511212 323854
rect 511276 323852 511282 323916
rect 279926 323718 287070 323778
rect 91737 323642 91803 323645
rect 95877 323642 95943 323645
rect 282269 323642 282335 323645
rect 91737 323640 95943 323642
rect 91737 323584 91742 323640
rect 91798 323584 95882 323640
rect 95938 323584 95943 323640
rect 91737 323582 95943 323584
rect 91737 323579 91803 323582
rect 95877 323579 95943 323582
rect 279926 323640 282335 323642
rect 279926 323584 282274 323640
rect 282330 323584 282335 323640
rect 279926 323582 282335 323584
rect 230289 323234 230355 323237
rect 230289 323232 239690 323234
rect 230289 323176 230294 323232
rect 230350 323176 239690 323232
rect 230289 323174 239690 323176
rect 230289 323171 230355 323174
rect 239630 323166 239690 323174
rect 239630 323106 240212 323166
rect 279926 323068 279986 323582
rect 282269 323579 282335 323582
rect 541065 322282 541131 322285
rect 287010 322280 541131 322282
rect 228817 322146 228883 322149
rect 279926 322146 279986 322252
rect 287010 322224 541070 322280
rect 541126 322224 541131 322280
rect 287010 322222 541131 322224
rect 287010 322146 287070 322222
rect 541065 322219 541131 322222
rect 228817 322144 239690 322146
rect 228817 322088 228822 322144
rect 228878 322088 239690 322144
rect 228817 322086 239690 322088
rect 279926 322086 287070 322146
rect 228817 322083 228883 322086
rect 239630 322078 239690 322086
rect 239630 322018 240212 322078
rect 540973 321466 541039 321469
rect 287010 321464 541039 321466
rect 279926 321330 279986 321436
rect 287010 321408 540978 321464
rect 541034 321408 541039 321464
rect 287010 321406 541039 321408
rect 287010 321330 287070 321406
rect 540973 321403 541039 321406
rect 279926 321270 287070 321330
rect 236821 321058 236887 321061
rect 236821 321056 239690 321058
rect 236821 321000 236826 321056
rect 236882 321000 239690 321056
rect 236821 320998 239690 321000
rect 236821 320995 236887 320998
rect 239630 320990 239690 320998
rect 239630 320930 240212 320990
rect 541382 320650 541388 320652
rect 279926 320514 279986 320620
rect 287010 320590 541388 320650
rect 287010 320514 287070 320590
rect 541382 320588 541388 320590
rect 541452 320588 541458 320652
rect 279926 320454 287070 320514
rect 231669 319970 231735 319973
rect 231669 319968 239690 319970
rect 231669 319912 231674 319968
rect 231730 319912 239690 319968
rect 231669 319910 239690 319912
rect 231669 319907 231735 319910
rect 239630 319902 239690 319910
rect 239630 319842 240212 319902
rect 541014 319834 541020 319836
rect 279926 319698 279986 319804
rect 287010 319774 541020 319834
rect 287010 319698 287070 319774
rect 541014 319772 541020 319774
rect 541084 319772 541090 319836
rect 279926 319638 287070 319698
rect 282177 319562 282243 319565
rect 279926 319560 282243 319562
rect 279926 319504 282182 319560
rect 282238 319504 282243 319560
rect 279926 319502 282243 319504
rect 169017 319426 169083 319429
rect 103470 319424 169083 319426
rect -960 319290 480 319380
rect 103470 319368 169022 319424
rect 169078 319368 169083 319424
rect 103470 319366 169083 319368
rect 99005 319290 99071 319293
rect 103470 319290 103530 319366
rect 169017 319363 169083 319366
rect -960 319288 103530 319290
rect -960 319232 99010 319288
rect 99066 319232 103530 319288
rect -960 319230 103530 319232
rect -960 319140 480 319230
rect 99005 319227 99071 319230
rect 279926 318988 279986 319502
rect 282177 319499 282243 319502
rect 239814 318754 240212 318814
rect 230381 318746 230447 318749
rect 239814 318746 239874 318754
rect 230381 318744 239874 318746
rect 230381 318688 230386 318744
rect 230442 318688 239874 318744
rect 230381 318686 239874 318688
rect 454677 318746 454743 318749
rect 456057 318746 456123 318749
rect 454677 318744 456123 318746
rect 454677 318688 454682 318744
rect 454738 318688 456062 318744
rect 456118 318688 456123 318744
rect 454677 318686 456123 318688
rect 230381 318683 230447 318686
rect 454677 318683 454743 318686
rect 456057 318683 456123 318686
rect 543774 318202 543780 318204
rect 279926 318066 279986 318172
rect 287010 318142 543780 318202
rect 287010 318066 287070 318142
rect 543774 318140 543780 318142
rect 543844 318140 543850 318204
rect 279926 318006 287070 318066
rect 228725 317794 228791 317797
rect 228725 317792 239690 317794
rect 228725 317736 228730 317792
rect 228786 317736 239690 317792
rect 228725 317734 239690 317736
rect 228725 317731 228791 317734
rect 239630 317726 239690 317734
rect 239630 317666 240212 317726
rect 522430 317386 522436 317388
rect 279926 317250 279986 317356
rect 287010 317326 522436 317386
rect 287010 317250 287070 317326
rect 522430 317324 522436 317326
rect 522500 317324 522506 317388
rect 279926 317190 287070 317250
rect 282361 317114 282427 317117
rect 279926 317112 282427 317114
rect 279926 317056 282366 317112
rect 282422 317056 282427 317112
rect 279926 317054 282427 317056
rect 8109 316706 8175 316709
rect 228725 316706 228791 316709
rect 8109 316704 228791 316706
rect 8109 316648 8114 316704
rect 8170 316648 228730 316704
rect 228786 316648 228791 316704
rect 8109 316646 228791 316648
rect 8109 316643 8175 316646
rect 228725 316643 228791 316646
rect 228909 316706 228975 316709
rect 228909 316704 239690 316706
rect 228909 316648 228914 316704
rect 228970 316648 239690 316704
rect 228909 316646 239690 316648
rect 228909 316643 228975 316646
rect 239630 316638 239690 316646
rect 239630 316578 240212 316638
rect 279926 316540 279986 317054
rect 282361 317051 282427 317054
rect 539542 315754 539548 315756
rect 236729 315618 236795 315621
rect 279926 315618 279986 315724
rect 287010 315694 539548 315754
rect 287010 315618 287070 315694
rect 539542 315692 539548 315694
rect 539612 315692 539618 315756
rect 236729 315616 239690 315618
rect 236729 315560 236734 315616
rect 236790 315560 239690 315616
rect 236729 315558 239690 315560
rect 279926 315558 287070 315618
rect 236729 315555 236795 315558
rect 239630 315550 239690 315558
rect 239630 315490 240212 315550
rect 282453 315482 282519 315485
rect 279926 315480 282519 315482
rect 279926 315424 282458 315480
rect 282514 315424 282519 315480
rect 279926 315422 282519 315424
rect 279926 314908 279986 315422
rect 282453 315419 282519 315422
rect 232957 314530 233023 314533
rect 232957 314528 239690 314530
rect 232957 314472 232962 314528
rect 233018 314472 239690 314528
rect 232957 314470 239690 314472
rect 232957 314467 233023 314470
rect 239630 314462 239690 314470
rect 239630 314402 240212 314462
rect 539726 314122 539732 314124
rect 279926 313986 279986 314092
rect 287010 314062 539732 314122
rect 287010 313986 287070 314062
rect 539726 314060 539732 314062
rect 539796 314060 539802 314124
rect 279926 313926 287070 313986
rect 282545 313850 282611 313853
rect 279926 313848 282611 313850
rect 279926 313792 282550 313848
rect 282606 313792 282611 313848
rect 279926 313790 282611 313792
rect 231577 313442 231643 313445
rect 231577 313440 239690 313442
rect 231577 313384 231582 313440
rect 231638 313384 239690 313440
rect 231577 313382 239690 313384
rect 231577 313379 231643 313382
rect 239630 313374 239690 313382
rect 239630 313314 240212 313374
rect 279926 313276 279986 313790
rect 282545 313787 282611 313790
rect 539910 312490 539916 312492
rect 236913 312354 236979 312357
rect 279926 312354 279986 312460
rect 287010 312430 539916 312490
rect 287010 312354 287070 312430
rect 539910 312428 539916 312430
rect 539980 312428 539986 312492
rect 236913 312352 239690 312354
rect 236913 312296 236918 312352
rect 236974 312296 239690 312352
rect 236913 312294 239690 312296
rect 279926 312294 287070 312354
rect 236913 312291 236979 312294
rect 239630 312286 239690 312294
rect 239630 312226 240212 312286
rect 580206 312020 580212 312084
rect 580276 312082 580282 312084
rect 583520 312082 584960 312172
rect 580276 312022 584960 312082
rect 580276 312020 580282 312022
rect 95877 311946 95943 311949
rect 99373 311946 99439 311949
rect 95877 311944 99439 311946
rect 95877 311888 95882 311944
rect 95938 311888 99378 311944
rect 99434 311888 99439 311944
rect 583520 311932 584960 312022
rect 95877 311886 99439 311888
rect 95877 311883 95943 311886
rect 99373 311883 99439 311886
rect 279926 311750 281826 311810
rect 279926 311644 279986 311750
rect 281766 311676 281826 311750
rect 281758 311612 281764 311676
rect 281828 311612 281834 311676
rect 233049 311266 233115 311269
rect 233049 311264 239690 311266
rect 233049 311208 233054 311264
rect 233110 311208 239690 311264
rect 233049 311206 239690 311208
rect 233049 311203 233115 311206
rect 239630 311198 239690 311206
rect 239630 311138 240212 311198
rect 282310 311068 282316 311132
rect 282380 311130 282386 311132
rect 539358 311130 539364 311132
rect 282380 311070 539364 311130
rect 282380 311068 282386 311070
rect 539358 311068 539364 311070
rect 539428 311068 539434 311132
rect 279926 310934 282010 310994
rect 279926 310828 279986 310934
rect 281950 310860 282010 310934
rect 281942 310796 281948 310860
rect 282012 310796 282018 310860
rect 236545 310178 236611 310181
rect 236545 310176 239690 310178
rect 236545 310120 236550 310176
rect 236606 310120 239690 310176
rect 236545 310118 239690 310120
rect 236545 310115 236611 310118
rect 239630 310110 239690 310118
rect 279926 310118 282194 310178
rect 239630 310050 240212 310110
rect 279926 310012 279986 310118
rect 282134 310044 282194 310118
rect 282126 309980 282132 310044
rect 282196 309980 282202 310044
rect 279926 309302 287070 309362
rect 279926 309196 279986 309302
rect 287010 309226 287070 309302
rect 522246 309226 522252 309228
rect 287010 309166 522252 309226
rect 522246 309164 522252 309166
rect 522316 309164 522322 309228
rect 229001 309090 229067 309093
rect 229001 309088 239690 309090
rect 229001 309032 229006 309088
rect 229062 309032 239690 309088
rect 229001 309030 239690 309032
rect 229001 309027 229067 309030
rect 239630 309022 239690 309030
rect 239630 308962 240212 309022
rect 537518 308410 537524 308412
rect 279926 308274 279986 308380
rect 287010 308350 537524 308410
rect 287010 308274 287070 308350
rect 537518 308348 537524 308350
rect 537588 308348 537594 308412
rect 279926 308214 287070 308274
rect 233877 308002 233943 308005
rect 233877 308000 239690 308002
rect 233877 307944 233882 308000
rect 233938 307944 239690 308000
rect 233877 307942 239690 307944
rect 233877 307939 233943 307942
rect 239630 307934 239690 307942
rect 239630 307874 240212 307934
rect 99373 307730 99439 307733
rect 102041 307730 102107 307733
rect 99373 307728 102107 307730
rect 99373 307672 99378 307728
rect 99434 307672 102046 307728
rect 102102 307672 102107 307728
rect 99373 307670 102107 307672
rect 99373 307667 99439 307670
rect 102041 307667 102107 307670
rect 483606 307594 483612 307596
rect 279926 307458 279986 307564
rect 287010 307534 483612 307594
rect 287010 307458 287070 307534
rect 483606 307532 483612 307534
rect 483676 307532 483682 307596
rect 279926 307398 287070 307458
rect 234429 306914 234495 306917
rect 234429 306912 239690 306914
rect 234429 306856 234434 306912
rect 234490 306856 239690 306912
rect 234429 306854 239690 306856
rect 234429 306851 234495 306854
rect 239630 306846 239690 306854
rect 239630 306786 240212 306846
rect 298686 306778 298692 306780
rect 279926 306642 279986 306748
rect 287010 306718 298692 306778
rect 287010 306642 287070 306718
rect 298686 306716 298692 306718
rect 298756 306716 298762 306780
rect 279926 306582 287070 306642
rect -960 306234 480 306324
rect 228398 306234 228404 306236
rect -960 306174 228404 306234
rect -960 306084 480 306174
rect 228398 306172 228404 306174
rect 228468 306172 228474 306236
rect 279926 306038 287070 306098
rect 279926 305932 279986 306038
rect 287010 305962 287070 306038
rect 287646 305962 287652 305964
rect 287010 305902 287652 305962
rect 287646 305900 287652 305902
rect 287716 305900 287722 305964
rect 235349 305826 235415 305829
rect 235349 305824 239690 305826
rect 235349 305768 235354 305824
rect 235410 305768 239690 305824
rect 235349 305766 239690 305768
rect 235349 305763 235415 305766
rect 239630 305758 239690 305766
rect 239630 305698 240212 305758
rect 279926 305222 287070 305282
rect 279926 305116 279986 305222
rect 287010 305146 287070 305222
rect 518014 305146 518020 305148
rect 287010 305086 518020 305146
rect 518014 305084 518020 305086
rect 518084 305084 518090 305148
rect 235165 304738 235231 304741
rect 235165 304736 239690 304738
rect 235165 304680 235170 304736
rect 235226 304680 239690 304736
rect 235165 304678 239690 304680
rect 235165 304675 235231 304678
rect 239630 304670 239690 304678
rect 239630 304610 240212 304670
rect 102041 304602 102107 304605
rect 104801 304602 104867 304605
rect 102041 304600 104867 304602
rect 102041 304544 102046 304600
rect 102102 304544 104806 304600
rect 104862 304544 104867 304600
rect 102041 304542 104867 304544
rect 102041 304539 102107 304542
rect 104801 304539 104867 304542
rect 279926 304406 287070 304466
rect 279926 304300 279986 304406
rect 287010 304330 287070 304406
rect 506974 304330 506980 304332
rect 287010 304270 506980 304330
rect 506974 304268 506980 304270
rect 507044 304268 507050 304332
rect 239630 303522 240212 303582
rect 235257 303514 235323 303517
rect 239630 303514 239690 303522
rect 508446 303514 508452 303516
rect 235257 303512 239690 303514
rect 235257 303456 235262 303512
rect 235318 303456 239690 303512
rect 235257 303454 239690 303456
rect 235257 303451 235323 303454
rect 279926 303378 279986 303484
rect 287010 303454 508452 303514
rect 287010 303378 287070 303454
rect 508446 303452 508452 303454
rect 508516 303452 508522 303516
rect 279926 303318 287070 303378
rect 279926 302774 282378 302834
rect 279926 302668 279986 302774
rect 282318 302700 282378 302774
rect 282310 302636 282316 302700
rect 282380 302636 282386 302700
rect 238150 302500 238156 302564
rect 238220 302562 238226 302564
rect 238220 302502 239690 302562
rect 238220 302500 238226 302502
rect 239630 302494 239690 302502
rect 239630 302434 240212 302494
rect 279926 301958 287070 302018
rect 279926 301852 279986 301958
rect 287010 301882 287070 301958
rect 537334 301882 537340 301884
rect 287010 301822 537340 301882
rect 537334 301820 537340 301822
rect 537404 301820 537410 301884
rect 79133 301474 79199 301477
rect 125593 301474 125659 301477
rect 79133 301472 125659 301474
rect 79133 301416 79138 301472
rect 79194 301416 125598 301472
rect 125654 301416 125659 301472
rect 79133 301414 125659 301416
rect 79133 301411 79199 301414
rect 125593 301411 125659 301414
rect 235441 301474 235507 301477
rect 235441 301472 239690 301474
rect 235441 301416 235446 301472
rect 235502 301416 239690 301472
rect 235441 301414 239690 301416
rect 235441 301411 235507 301414
rect 239630 301406 239690 301414
rect 239630 301346 240212 301406
rect 279926 301142 287070 301202
rect 279926 301036 279986 301142
rect 287010 301066 287070 301142
rect 534574 301066 534580 301068
rect 287010 301006 534580 301066
rect 534574 301004 534580 301006
rect 534644 301004 534650 301068
rect 104801 300658 104867 300661
rect 109677 300658 109743 300661
rect 104801 300656 109743 300658
rect 104801 300600 104806 300656
rect 104862 300600 109682 300656
rect 109738 300600 109743 300656
rect 104801 300598 109743 300600
rect 104801 300595 104867 300598
rect 109677 300595 109743 300598
rect 235533 300386 235599 300389
rect 235533 300384 239690 300386
rect 235533 300328 235538 300384
rect 235594 300328 239690 300384
rect 235533 300326 239690 300328
rect 235533 300323 235599 300326
rect 239630 300318 239690 300326
rect 279926 300326 287070 300386
rect 239630 300258 240212 300318
rect 279926 300220 279986 300326
rect 287010 300250 287070 300326
rect 526294 300250 526300 300252
rect 287010 300190 526300 300250
rect 526294 300188 526300 300190
rect 526364 300188 526370 300252
rect 279926 299510 281090 299570
rect 279926 299404 279986 299510
rect 280889 299434 280955 299437
rect 280110 299432 280955 299434
rect 280110 299376 280894 299432
rect 280950 299376 280955 299432
rect 280110 299374 280955 299376
rect 281030 299434 281090 299510
rect 282177 299434 282243 299437
rect 281030 299432 282243 299434
rect 281030 299376 282182 299432
rect 282238 299376 282243 299432
rect 281030 299374 282243 299376
rect 236637 299298 236703 299301
rect 280110 299298 280170 299374
rect 280889 299371 280955 299374
rect 282177 299371 282243 299374
rect 236637 299296 239690 299298
rect 236637 299240 236642 299296
rect 236698 299240 239690 299296
rect 236637 299238 239690 299240
rect 236637 299235 236703 299238
rect 239630 299230 239690 299238
rect 279926 299238 280170 299298
rect 239630 299170 240212 299230
rect 59261 298754 59327 298757
rect 83457 298754 83523 298757
rect 59261 298752 83523 298754
rect 59261 298696 59266 298752
rect 59322 298696 83462 298752
rect 83518 298696 83523 298752
rect 59261 298694 83523 298696
rect 59261 298691 59327 298694
rect 83457 298691 83523 298694
rect 279926 298588 279986 299238
rect 497457 298754 497523 298757
rect 583520 298754 584960 298844
rect 497457 298752 584960 298754
rect 497457 298696 497462 298752
rect 497518 298696 584960 298752
rect 497457 298694 584960 298696
rect 497457 298691 497523 298694
rect 583520 298604 584960 298694
rect 239814 298082 240212 298142
rect 239438 298012 239444 298076
rect 239508 298074 239514 298076
rect 239814 298074 239874 298082
rect 280981 298074 281047 298077
rect 239508 298014 239874 298074
rect 279926 298072 281047 298074
rect 279926 298016 280986 298072
rect 281042 298016 281047 298072
rect 279926 298014 281047 298016
rect 239508 298012 239514 298014
rect 279926 297772 279986 298014
rect 280981 298011 281047 298014
rect 280705 297802 280771 297805
rect 280110 297800 280771 297802
rect 280110 297744 280710 297800
rect 280766 297744 280771 297800
rect 280110 297742 280771 297744
rect 280110 297666 280170 297742
rect 280705 297739 280771 297742
rect 279926 297606 280170 297666
rect 233785 297122 233851 297125
rect 233785 297120 239690 297122
rect 233785 297064 233790 297120
rect 233846 297064 239690 297120
rect 233785 297062 239690 297064
rect 233785 297059 233851 297062
rect 239630 297054 239690 297062
rect 239630 296994 240212 297054
rect 279926 296956 279986 297606
rect 280613 296442 280679 296445
rect 279926 296440 280679 296442
rect 279926 296384 280618 296440
rect 280674 296384 280679 296440
rect 279926 296382 280679 296384
rect 279926 296140 279986 296382
rect 280613 296379 280679 296382
rect 233969 296034 234035 296037
rect 280797 296034 280863 296037
rect 233969 296032 239690 296034
rect 233969 295976 233974 296032
rect 234030 295976 239690 296032
rect 233969 295974 239690 295976
rect 233969 295971 234035 295974
rect 239630 295966 239690 295974
rect 279926 296032 280863 296034
rect 279926 295976 280802 296032
rect 280858 295976 280863 296032
rect 279926 295974 280863 295976
rect 239630 295906 240212 295966
rect 109677 295354 109743 295357
rect 113817 295354 113883 295357
rect 109677 295352 113883 295354
rect 109677 295296 109682 295352
rect 109738 295296 113822 295352
rect 113878 295296 113883 295352
rect 279926 295324 279986 295974
rect 280797 295971 280863 295974
rect 109677 295294 113883 295296
rect 109677 295291 109743 295294
rect 113817 295291 113883 295294
rect 280337 295218 280403 295221
rect 279926 295216 280403 295218
rect 279926 295160 280342 295216
rect 280398 295160 280403 295216
rect 279926 295158 280403 295160
rect 234153 294946 234219 294949
rect 234153 294944 239690 294946
rect 234153 294888 234158 294944
rect 234214 294888 239690 294944
rect 234153 294886 239690 294888
rect 234153 294883 234219 294886
rect 239630 294878 239690 294886
rect 239630 294818 240212 294878
rect 279926 294508 279986 295158
rect 280337 295155 280403 295158
rect 280429 293858 280495 293861
rect 279926 293856 280495 293858
rect 279926 293800 280434 293856
rect 280490 293800 280495 293856
rect 279926 293798 280495 293800
rect 239622 293728 239628 293792
rect 239692 293790 239698 293792
rect 239692 293730 240212 293790
rect 239692 293728 239698 293730
rect 279926 293692 279986 293798
rect 280429 293795 280495 293798
rect 281717 293586 281783 293589
rect 279926 293584 281783 293586
rect 279926 293528 281722 293584
rect 281778 293528 281783 293584
rect 279926 293526 281783 293528
rect -960 293178 480 293268
rect 122046 293178 122052 293180
rect -960 293118 122052 293178
rect -960 293028 480 293118
rect 122046 293116 122052 293118
rect 122116 293116 122122 293180
rect 279926 292876 279986 293526
rect 281717 293523 281783 293526
rect 238293 292770 238359 292773
rect 238293 292768 239690 292770
rect 238293 292712 238298 292768
rect 238354 292712 239690 292768
rect 238293 292710 239690 292712
rect 238293 292707 238359 292710
rect 239630 292702 239690 292710
rect 239630 292642 240212 292702
rect 280521 292498 280587 292501
rect 279926 292496 280587 292498
rect 279926 292440 280526 292496
rect 280582 292440 280587 292496
rect 279926 292438 280587 292440
rect 279926 292060 279986 292438
rect 280521 292435 280587 292438
rect 237833 291682 237899 291685
rect 237833 291680 239690 291682
rect 237833 291624 237838 291680
rect 237894 291624 239690 291680
rect 237833 291622 239690 291624
rect 237833 291619 237899 291622
rect 239630 291614 239690 291622
rect 239630 291554 240212 291614
rect 279926 291350 280722 291410
rect 279926 291244 279986 291350
rect 280662 291276 280722 291350
rect 280654 291212 280660 291276
rect 280724 291212 280730 291276
rect 281625 291138 281691 291141
rect 279926 291136 281691 291138
rect 279926 291080 281630 291136
rect 281686 291080 281691 291136
rect 279926 291078 281691 291080
rect 234245 290594 234311 290597
rect 234245 290592 239690 290594
rect 234245 290536 234250 290592
rect 234306 290536 239690 290592
rect 234245 290534 239690 290536
rect 234245 290531 234311 290534
rect 239630 290526 239690 290534
rect 239630 290466 240212 290526
rect 279926 290428 279986 291078
rect 281625 291075 281691 291078
rect 235942 289716 235948 289780
rect 236012 289778 236018 289780
rect 237005 289778 237071 289781
rect 282177 289778 282243 289781
rect 236012 289776 237071 289778
rect 236012 289720 237010 289776
rect 237066 289720 237071 289776
rect 236012 289718 237071 289720
rect 236012 289716 236018 289718
rect 237005 289715 237071 289718
rect 279926 289776 282243 289778
rect 279926 289720 282182 289776
rect 282238 289720 282243 289776
rect 279926 289718 282243 289720
rect 236126 289580 236132 289644
rect 236196 289642 236202 289644
rect 237966 289642 237972 289644
rect 236196 289582 237972 289642
rect 236196 289580 236202 289582
rect 237966 289580 237972 289582
rect 238036 289580 238042 289644
rect 279926 289612 279986 289718
rect 282177 289715 282243 289718
rect 238109 289506 238175 289509
rect 281533 289506 281599 289509
rect 238109 289504 239690 289506
rect 238109 289448 238114 289504
rect 238170 289448 239690 289504
rect 238109 289446 239690 289448
rect 238109 289443 238175 289446
rect 239630 289438 239690 289446
rect 279926 289504 281599 289506
rect 279926 289448 281538 289504
rect 281594 289448 281599 289504
rect 279926 289446 281599 289448
rect 239630 289378 240212 289438
rect 279926 288796 279986 289446
rect 281533 289443 281599 289446
rect 238201 288418 238267 288421
rect 238201 288416 239690 288418
rect 238201 288360 238206 288416
rect 238262 288360 239690 288416
rect 238201 288358 239690 288360
rect 238201 288355 238267 288358
rect 239630 288350 239690 288358
rect 239630 288290 240212 288350
rect 282085 288282 282151 288285
rect 279926 288280 282151 288282
rect 279926 288224 282090 288280
rect 282146 288224 282151 288280
rect 279926 288222 282151 288224
rect 279926 287980 279986 288222
rect 282085 288219 282151 288222
rect 282729 288010 282795 288013
rect 280662 288008 282795 288010
rect 280662 287952 282734 288008
rect 282790 287952 282795 288008
rect 280662 287950 282795 287952
rect 280662 287874 280722 287950
rect 282729 287947 282795 287950
rect 279926 287814 280722 287874
rect 234337 287330 234403 287333
rect 234337 287328 239690 287330
rect 234337 287272 234342 287328
rect 234398 287272 239690 287328
rect 234337 287270 239690 287272
rect 234337 287267 234403 287270
rect 239630 287262 239690 287270
rect 239630 287202 240212 287262
rect 279926 287164 279986 287814
rect 282637 286650 282703 286653
rect 279926 286648 282703 286650
rect 279926 286592 282642 286648
rect 282698 286592 282703 286648
rect 279926 286590 282703 286592
rect 11646 286316 11652 286380
rect 11716 286378 11722 286380
rect 238150 286378 238156 286380
rect 11716 286318 238156 286378
rect 11716 286316 11722 286318
rect 238150 286316 238156 286318
rect 238220 286316 238226 286380
rect 279926 286348 279986 286590
rect 282637 286587 282703 286590
rect 238385 286242 238451 286245
rect 238385 286240 239690 286242
rect 238385 286184 238390 286240
rect 238446 286184 239690 286240
rect 238385 286182 239690 286184
rect 238385 286179 238451 286182
rect 239630 286174 239690 286182
rect 239630 286114 240212 286174
rect 279926 285638 281826 285698
rect 279926 285532 279986 285638
rect 281533 285562 281599 285565
rect 280110 285560 281599 285562
rect 280110 285504 281538 285560
rect 281594 285504 281599 285560
rect 280110 285502 281599 285504
rect 281766 285562 281826 285638
rect 282637 285562 282703 285565
rect 281766 285560 282703 285562
rect 281766 285504 282642 285560
rect 282698 285504 282703 285560
rect 281766 285502 282703 285504
rect 280110 285426 280170 285502
rect 281533 285499 281599 285502
rect 282637 285499 282703 285502
rect 279926 285366 280170 285426
rect 237741 285154 237807 285157
rect 237741 285152 239690 285154
rect 237741 285096 237746 285152
rect 237802 285096 239690 285152
rect 237741 285094 239690 285096
rect 237741 285091 237807 285094
rect 239630 285086 239690 285094
rect 239630 285026 240212 285086
rect 279926 284716 279986 285366
rect 583520 285276 584960 285516
rect 282085 284202 282151 284205
rect 279926 284200 282151 284202
rect 279926 284144 282090 284200
rect 282146 284144 282151 284200
rect 279926 284142 282151 284144
rect 239581 284066 239647 284069
rect 239581 284064 239690 284066
rect 239581 284008 239586 284064
rect 239642 284008 239690 284064
rect 239581 284003 239690 284008
rect 239630 283998 239690 284003
rect 239630 283938 240212 283998
rect 279926 283900 279986 284142
rect 282085 284139 282151 284142
rect 283557 283658 283623 283661
rect 279926 283656 283623 283658
rect 279926 283600 283562 283656
rect 283618 283600 283623 283656
rect 279926 283598 283623 283600
rect 279926 283084 279986 283598
rect 283557 283595 283623 283598
rect 239814 282850 240212 282910
rect 239397 282842 239463 282845
rect 239814 282842 239874 282850
rect 239397 282840 239874 282842
rect 239397 282784 239402 282840
rect 239458 282784 239874 282840
rect 239397 282782 239874 282784
rect 239397 282779 239463 282782
rect 283465 282706 283531 282709
rect 279926 282704 283531 282706
rect 279926 282648 283470 282704
rect 283526 282648 283531 282704
rect 279926 282646 283531 282648
rect 279926 282268 279986 282646
rect 283465 282643 283531 282646
rect 239489 281890 239555 281893
rect 239489 281888 239690 281890
rect 239489 281832 239494 281888
rect 239550 281832 239690 281888
rect 239489 281830 239690 281832
rect 239489 281827 239555 281830
rect 239630 281822 239690 281830
rect 239630 281762 240212 281822
rect 281993 281482 282059 281485
rect 280110 281480 282059 281482
rect 279926 281346 279986 281452
rect 280110 281424 281998 281480
rect 282054 281424 282059 281480
rect 280110 281422 282059 281424
rect 280110 281346 280170 281422
rect 281993 281419 282059 281422
rect 279926 281286 280170 281346
rect 283649 281074 283715 281077
rect 279926 281072 283715 281074
rect 279926 281016 283654 281072
rect 283710 281016 283715 281072
rect 279926 281014 283715 281016
rect 239305 280802 239371 280805
rect 239305 280800 239690 280802
rect 239305 280744 239310 280800
rect 239366 280744 239690 280800
rect 239305 280742 239690 280744
rect 239305 280739 239371 280742
rect 239630 280734 239690 280742
rect 239630 280674 240212 280734
rect 279926 280636 279986 281014
rect 283649 281011 283715 281014
rect -960 279972 480 280212
rect 283373 280122 283439 280125
rect 279926 280120 283439 280122
rect 279926 280064 283378 280120
rect 283434 280064 283439 280120
rect 279926 280062 283439 280064
rect 279926 279820 279986 280062
rect 283373 280059 283439 280062
rect 237925 279714 237991 279717
rect 281993 279714 282059 279717
rect 237925 279712 239690 279714
rect 237925 279656 237930 279712
rect 237986 279656 239690 279712
rect 237925 279654 239690 279656
rect 237925 279651 237991 279654
rect 239630 279646 239690 279654
rect 279926 279712 282059 279714
rect 279926 279656 281998 279712
rect 282054 279656 282059 279712
rect 279926 279654 282059 279656
rect 239630 279586 240212 279646
rect 279926 279004 279986 279654
rect 281993 279651 282059 279654
rect 239857 278558 239923 278561
rect 239857 278556 240212 278558
rect 239857 278500 239862 278556
rect 239918 278500 240212 278556
rect 239857 278498 240212 278500
rect 239857 278495 239923 278498
rect 279926 277810 279986 278188
rect 492581 278082 492647 278085
rect 507853 278082 507919 278085
rect 492581 278080 507919 278082
rect 492581 278024 492586 278080
rect 492642 278024 507858 278080
rect 507914 278024 507919 278080
rect 492581 278022 507919 278024
rect 492581 278019 492647 278022
rect 507853 278019 507919 278022
rect 282821 277810 282887 277813
rect 279926 277808 282887 277810
rect 279926 277752 282826 277808
rect 282882 277752 282887 277808
rect 279926 277750 282887 277752
rect 282821 277747 282887 277750
rect 239857 277470 239923 277473
rect 239857 277468 240212 277470
rect 239857 277412 239862 277468
rect 239918 277412 240212 277468
rect 239857 277410 240212 277412
rect 239857 277407 239923 277410
rect 279926 277402 280170 277410
rect 282729 277402 282795 277405
rect 279926 277400 282795 277402
rect 279926 277350 282734 277400
rect 280110 277344 282734 277350
rect 282790 277344 282795 277400
rect 280110 277342 282795 277344
rect 282729 277339 282795 277342
rect 345606 276660 345612 276724
rect 345676 276722 345682 276724
rect 580206 276722 580212 276724
rect 345676 276662 580212 276722
rect 345676 276660 345682 276662
rect 580206 276660 580212 276662
rect 580276 276660 580282 276724
rect 239673 276382 239739 276385
rect 239673 276380 240212 276382
rect 239673 276324 239678 276380
rect 239734 276324 240212 276380
rect 239673 276322 240212 276324
rect 239673 276319 239739 276322
rect 279926 276314 279986 276556
rect 282821 276314 282887 276317
rect 279926 276312 282887 276314
rect 279926 276256 282826 276312
rect 282882 276256 282887 276312
rect 279926 276254 282887 276256
rect 282821 276251 282887 276254
rect 237649 275362 237715 275365
rect 237649 275360 239690 275362
rect 237649 275304 237654 275360
rect 237710 275304 239690 275360
rect 237649 275302 239690 275304
rect 237649 275299 237715 275302
rect 239630 275294 239690 275302
rect 239630 275234 240212 275294
rect 279926 275226 279986 275740
rect 282821 275226 282887 275229
rect 279926 275224 282887 275226
rect 279926 275168 282826 275224
rect 282882 275168 282887 275224
rect 279926 275166 282887 275168
rect 282821 275163 282887 275166
rect 279926 275030 287070 275090
rect 279926 274924 279986 275030
rect 287010 274954 287070 275030
rect 288801 274954 288867 274957
rect 287010 274952 288867 274954
rect 287010 274896 288806 274952
rect 288862 274896 288867 274952
rect 287010 274894 288867 274896
rect 288801 274891 288867 274894
rect 234061 274546 234127 274549
rect 237373 274546 237439 274549
rect 234061 274544 237439 274546
rect 234061 274488 234066 274544
rect 234122 274488 237378 274544
rect 237434 274488 237439 274544
rect 234061 274486 237439 274488
rect 234061 274483 234127 274486
rect 237373 274483 237439 274486
rect 238661 274274 238727 274277
rect 238661 274272 239690 274274
rect 238661 274216 238666 274272
rect 238722 274216 239690 274272
rect 238661 274214 239690 274216
rect 238661 274211 238727 274214
rect 239630 274206 239690 274214
rect 239630 274146 240212 274206
rect 14406 273804 14412 273868
rect 14476 273866 14482 273868
rect 237414 273866 237420 273868
rect 14476 273806 237420 273866
rect 14476 273804 14482 273806
rect 237414 273804 237420 273806
rect 237484 273804 237490 273868
rect 279926 273730 279986 274108
rect 282729 273730 282795 273733
rect 279926 273728 282795 273730
rect 279926 273672 282734 273728
rect 282790 273672 282795 273728
rect 279926 273670 282795 273672
rect 282729 273667 282795 273670
rect 279926 273322 280170 273356
rect 282821 273322 282887 273325
rect 279926 273320 282887 273322
rect 279926 273296 282826 273320
rect 279926 273292 279986 273296
rect 280110 273264 282826 273296
rect 282882 273264 282887 273320
rect 280110 273262 282887 273264
rect 282821 273259 282887 273262
rect 238017 273186 238083 273189
rect 238017 273184 239690 273186
rect 238017 273128 238022 273184
rect 238078 273128 239690 273184
rect 238017 273126 239690 273128
rect 238017 273123 238083 273126
rect 239630 273118 239690 273126
rect 239630 273058 240212 273118
rect 72509 272642 72575 272645
rect 112437 272642 112503 272645
rect 72509 272640 112503 272642
rect 72509 272584 72514 272640
rect 72570 272584 112442 272640
rect 112498 272584 112503 272640
rect 72509 272582 112503 272584
rect 72509 272579 72575 272582
rect 112437 272579 112503 272582
rect 4654 272444 4660 272508
rect 4724 272506 4730 272508
rect 238518 272506 238524 272508
rect 4724 272446 238524 272506
rect 4724 272444 4730 272446
rect 238518 272444 238524 272446
rect 238588 272444 238594 272508
rect 279926 272234 279986 272476
rect 282821 272234 282887 272237
rect 279926 272232 282887 272234
rect 279926 272176 282826 272232
rect 282882 272176 282887 272232
rect 279926 272174 282887 272176
rect 282821 272171 282887 272174
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 237373 272098 237439 272101
rect 237373 272096 239690 272098
rect 237373 272040 237378 272096
rect 237434 272040 239690 272096
rect 583520 272084 584960 272174
rect 237373 272038 239690 272040
rect 237373 272035 237439 272038
rect 239630 272030 239690 272038
rect 239630 271970 240212 272030
rect 279926 271146 279986 271660
rect 282729 271146 282795 271149
rect 279926 271144 282795 271146
rect 279926 271088 282734 271144
rect 282790 271088 282795 271144
rect 279926 271086 282795 271088
rect 282729 271083 282795 271086
rect 230473 271010 230539 271013
rect 230473 271008 239690 271010
rect 230473 270952 230478 271008
rect 230534 270952 239690 271008
rect 230473 270950 239690 270952
rect 230473 270947 230539 270950
rect 239630 270942 239690 270950
rect 239630 270882 240212 270942
rect 279926 270738 279986 270844
rect 282821 270738 282887 270741
rect 279926 270736 282887 270738
rect 279926 270680 282826 270736
rect 282882 270680 282887 270736
rect 279926 270678 282887 270680
rect 282821 270675 282887 270678
rect 283189 270466 283255 270469
rect 279926 270464 283255 270466
rect 279926 270408 283194 270464
rect 283250 270408 283255 270464
rect 279926 270406 283255 270408
rect 279926 270028 279986 270406
rect 283189 270403 283255 270406
rect 442257 270466 442323 270469
rect 447777 270466 447843 270469
rect 442257 270464 447843 270466
rect 442257 270408 442262 270464
rect 442318 270408 447782 270464
rect 447838 270408 447843 270464
rect 442257 270406 447843 270408
rect 442257 270403 442323 270406
rect 447777 270403 447843 270406
rect 281901 270058 281967 270061
rect 280662 270056 281967 270058
rect 280662 270000 281906 270056
rect 281962 270000 281967 270056
rect 280662 269998 281967 270000
rect 226885 269922 226951 269925
rect 280662 269922 280722 269998
rect 281901 269995 281967 269998
rect 226885 269920 239690 269922
rect 226885 269864 226890 269920
rect 226946 269864 239690 269920
rect 226885 269862 239690 269864
rect 226885 269859 226951 269862
rect 239630 269854 239690 269862
rect 279926 269862 280722 269922
rect 239630 269794 240212 269854
rect 279926 269212 279986 269862
rect 283281 268970 283347 268973
rect 279926 268968 283347 268970
rect 279926 268912 283286 268968
rect 283342 268912 283347 268968
rect 279926 268910 283347 268912
rect 223297 268834 223363 268837
rect 223297 268832 239690 268834
rect 223297 268776 223302 268832
rect 223358 268776 239690 268832
rect 223297 268774 239690 268776
rect 223297 268771 223363 268774
rect 239630 268766 239690 268774
rect 239630 268706 240212 268766
rect 279926 268396 279986 268910
rect 283281 268907 283347 268910
rect 219709 267746 219775 267749
rect 219709 267744 239690 267746
rect 219709 267688 219714 267744
rect 219770 267688 239690 267744
rect 219709 267686 239690 267688
rect 219709 267683 219775 267686
rect 239630 267678 239690 267686
rect 279926 267686 280170 267746
rect 239630 267618 240212 267678
rect 279926 267580 279986 267686
rect 280110 267610 280170 267686
rect 281901 267610 281967 267613
rect 280110 267608 281967 267610
rect 280110 267552 281906 267608
rect 281962 267552 281967 267608
rect 280110 267550 281967 267552
rect 281901 267547 281967 267550
rect 283097 267338 283163 267341
rect 279926 267336 283163 267338
rect -960 267202 480 267292
rect 279926 267280 283102 267336
rect 283158 267280 283163 267336
rect 279926 267278 283163 267280
rect 100569 267202 100635 267205
rect -960 267200 103530 267202
rect -960 267144 100574 267200
rect 100630 267144 103530 267200
rect -960 267142 103530 267144
rect -960 267052 480 267142
rect 100569 267139 100635 267142
rect 103470 267066 103530 267142
rect 173157 267066 173223 267069
rect 103470 267064 173223 267066
rect 103470 267008 173162 267064
rect 173218 267008 173223 267064
rect 103470 267006 173223 267008
rect 173157 267003 173223 267006
rect 279926 266764 279986 267278
rect 283097 267275 283163 267278
rect 216121 266658 216187 266661
rect 216121 266656 239690 266658
rect 216121 266600 216126 266656
rect 216182 266600 239690 266656
rect 216121 266598 239690 266600
rect 216121 266595 216187 266598
rect 239630 266590 239690 266598
rect 239630 266530 240212 266590
rect 279926 266054 284586 266114
rect 279926 265948 279986 266054
rect 281809 265978 281875 265981
rect 284526 265980 284586 266054
rect 280110 265976 281875 265978
rect 280110 265920 281814 265976
rect 281870 265920 281875 265976
rect 280110 265918 281875 265920
rect 280110 265842 280170 265918
rect 281809 265915 281875 265918
rect 284518 265916 284524 265980
rect 284588 265916 284594 265980
rect 279926 265782 280170 265842
rect 64505 265570 64571 265573
rect 94129 265570 94195 265573
rect 64505 265568 94195 265570
rect 64505 265512 64510 265568
rect 64566 265512 94134 265568
rect 94190 265512 94195 265568
rect 64505 265510 94195 265512
rect 64505 265507 64571 265510
rect 94129 265507 94195 265510
rect 212533 265570 212599 265573
rect 212533 265568 239690 265570
rect 212533 265512 212538 265568
rect 212594 265512 239690 265568
rect 212533 265510 239690 265512
rect 212533 265507 212599 265510
rect 239630 265502 239690 265510
rect 239630 265442 240212 265502
rect 279926 265132 279986 265782
rect 208945 264482 209011 264485
rect 208945 264480 239690 264482
rect 208945 264424 208950 264480
rect 209006 264424 239690 264480
rect 208945 264422 239690 264424
rect 208945 264419 209011 264422
rect 239630 264414 239690 264422
rect 279926 264422 286058 264482
rect 239630 264354 240212 264414
rect 279926 264316 279986 264422
rect 285998 264348 286058 264422
rect 285990 264284 285996 264348
rect 286060 264284 286066 264348
rect 279926 263606 280538 263666
rect 102133 263530 102199 263533
rect 105537 263530 105603 263533
rect 102133 263528 105603 263530
rect 102133 263472 102138 263528
rect 102194 263472 105542 263528
rect 105598 263472 105603 263528
rect 279926 263500 279986 263606
rect 280245 263530 280311 263533
rect 280110 263528 280311 263530
rect 102133 263470 105603 263472
rect 102133 263467 102199 263470
rect 105537 263467 105603 263470
rect 280110 263472 280250 263528
rect 280306 263472 280311 263528
rect 280110 263470 280311 263472
rect 280478 263530 280538 263606
rect 284702 263530 284708 263532
rect 280478 263470 284708 263530
rect 205357 263394 205423 263397
rect 280110 263394 280170 263470
rect 280245 263467 280311 263470
rect 284702 263468 284708 263470
rect 284772 263468 284778 263532
rect 205357 263392 239690 263394
rect 205357 263336 205362 263392
rect 205418 263336 239690 263392
rect 205357 263334 239690 263336
rect 205357 263331 205423 263334
rect 239630 263326 239690 263334
rect 279926 263334 280170 263394
rect 239630 263266 240212 263326
rect 108941 263258 109007 263261
rect 138657 263258 138723 263261
rect 108941 263256 138723 263258
rect 108941 263200 108946 263256
rect 109002 263200 138662 263256
rect 138718 263200 138723 263256
rect 108941 263198 138723 263200
rect 108941 263195 109007 263198
rect 138657 263195 138723 263198
rect 105905 263122 105971 263125
rect 135897 263122 135963 263125
rect 105905 263120 135963 263122
rect 105905 263064 105910 263120
rect 105966 263064 135902 263120
rect 135958 263064 135963 263120
rect 105905 263062 135963 263064
rect 105905 263059 105971 263062
rect 135897 263059 135963 263062
rect 50981 262986 51047 262989
rect 65517 262986 65583 262989
rect 50981 262984 65583 262986
rect 50981 262928 50986 262984
rect 51042 262928 65522 262984
rect 65578 262928 65583 262984
rect 50981 262926 65583 262928
rect 50981 262923 51047 262926
rect 65517 262923 65583 262926
rect 107561 262986 107627 262989
rect 137277 262986 137343 262989
rect 107561 262984 137343 262986
rect 107561 262928 107566 262984
rect 107622 262928 137282 262984
rect 137338 262928 137343 262984
rect 107561 262926 137343 262928
rect 107561 262923 107627 262926
rect 137277 262923 137343 262926
rect 52913 262850 52979 262853
rect 69657 262850 69723 262853
rect 52913 262848 69723 262850
rect 52913 262792 52918 262848
rect 52974 262792 69662 262848
rect 69718 262792 69723 262848
rect 52913 262790 69723 262792
rect 52913 262787 52979 262790
rect 69657 262787 69723 262790
rect 104801 262850 104867 262853
rect 134517 262850 134583 262853
rect 104801 262848 134583 262850
rect 104801 262792 104806 262848
rect 104862 262792 134522 262848
rect 134578 262792 134583 262848
rect 104801 262790 134583 262792
rect 104801 262787 104867 262790
rect 134517 262787 134583 262790
rect 279926 262684 279986 263334
rect 4797 262306 4863 262309
rect 108941 262306 109007 262309
rect 4797 262304 109007 262306
rect 4797 262248 4802 262304
rect 4858 262248 108946 262304
rect 109002 262248 109007 262304
rect 4797 262246 109007 262248
rect 4797 262243 4863 262246
rect 108941 262243 109007 262246
rect 239814 262178 240212 262238
rect 201769 262170 201835 262173
rect 239814 262170 239874 262178
rect 201769 262168 239874 262170
rect 201769 262112 201774 262168
rect 201830 262112 239874 262168
rect 201769 262110 239874 262112
rect 201769 262107 201835 262110
rect 282821 262034 282887 262037
rect 279926 262032 282887 262034
rect 279926 261976 282826 262032
rect 282882 261976 282887 262032
rect 279926 261974 282887 261976
rect 279926 261868 279986 261974
rect 282821 261971 282887 261974
rect 47577 261218 47643 261221
rect 105905 261218 105971 261221
rect 47577 261216 105971 261218
rect 47577 261160 47582 261216
rect 47638 261160 105910 261216
rect 105966 261160 105971 261216
rect 47577 261158 105971 261160
rect 47577 261155 47643 261158
rect 105905 261155 105971 261158
rect 198181 261218 198247 261221
rect 198181 261216 239690 261218
rect 198181 261160 198186 261216
rect 198242 261160 239690 261216
rect 198181 261158 239690 261160
rect 198181 261155 198247 261158
rect 239630 261150 239690 261158
rect 279926 261158 281642 261218
rect 239630 261090 240212 261150
rect 40677 261082 40743 261085
rect 103789 261082 103855 261085
rect 104801 261082 104867 261085
rect 40677 261080 104867 261082
rect 40677 261024 40682 261080
rect 40738 261024 103794 261080
rect 103850 261024 104806 261080
rect 104862 261024 104867 261080
rect 279926 261052 279986 261158
rect 281582 261084 281642 261158
rect 40677 261022 104867 261024
rect 40677 261019 40743 261022
rect 103789 261019 103855 261022
rect 104801 261019 104867 261022
rect 281574 261020 281580 261084
rect 281644 261020 281650 261084
rect 35157 260946 35223 260949
rect 107561 260946 107627 260949
rect 35157 260944 107627 260946
rect 35157 260888 35162 260944
rect 35218 260888 107566 260944
rect 107622 260888 107627 260944
rect 35157 260886 107627 260888
rect 35157 260883 35223 260886
rect 107561 260883 107627 260886
rect 282545 260810 282611 260813
rect 279926 260808 282611 260810
rect 279926 260752 282550 260808
rect 282606 260752 282611 260808
rect 279926 260750 282611 260752
rect 194593 260266 194659 260269
rect 194593 260264 239690 260266
rect 194593 260208 194598 260264
rect 194654 260208 239690 260264
rect 279926 260236 279986 260750
rect 282545 260747 282611 260750
rect 194593 260206 239690 260208
rect 194593 260203 194659 260206
rect 54886 260068 54892 260132
rect 54956 260130 54962 260132
rect 238201 260130 238267 260133
rect 54956 260128 238267 260130
rect 54956 260072 238206 260128
rect 238262 260072 238267 260128
rect 54956 260070 238267 260072
rect 54956 260068 54962 260070
rect 238201 260067 238267 260070
rect 239630 260062 239690 260206
rect 239630 260002 240212 260062
rect 279926 259314 279986 259420
rect 285806 259314 285812 259316
rect 279926 259254 285812 259314
rect 285806 259252 285812 259254
rect 285876 259252 285882 259316
rect 222837 259042 222903 259045
rect 222837 259040 239690 259042
rect 222837 258984 222842 259040
rect 222898 258984 239690 259040
rect 222837 258982 239690 258984
rect 222837 258979 222903 258982
rect 239630 258974 239690 258982
rect 239630 258914 240212 258974
rect 287646 258844 287652 258908
rect 287716 258906 287722 258908
rect 583520 258906 584960 258996
rect 287716 258846 584960 258906
rect 287716 258844 287722 258846
rect 285622 258770 285628 258772
rect 279926 258710 285628 258770
rect 227478 258634 227484 258636
rect 109940 258574 227484 258634
rect 227478 258572 227484 258574
rect 227548 258572 227554 258636
rect 279926 258604 279986 258710
rect 285622 258708 285628 258710
rect 285692 258708 285698 258772
rect 583520 258756 584960 258846
rect 117957 257954 118023 257957
rect 287094 257954 287100 257956
rect 117957 257952 239690 257954
rect 117957 257896 117962 257952
rect 118018 257896 239690 257952
rect 117957 257894 239690 257896
rect 117957 257891 118023 257894
rect 239630 257886 239690 257894
rect 279926 257894 287100 257954
rect 239630 257826 240212 257886
rect 226742 257756 226748 257820
rect 226812 257818 226818 257820
rect 227621 257818 227687 257821
rect 226812 257816 227687 257818
rect 226812 257760 227626 257816
rect 227682 257760 227687 257816
rect 279926 257788 279986 257894
rect 287094 257892 287100 257894
rect 287164 257892 287170 257956
rect 226812 257758 227687 257760
rect 226812 257756 226818 257758
rect 227621 257755 227687 257758
rect 282545 257410 282611 257413
rect 279926 257408 282611 257410
rect 279926 257352 282550 257408
rect 282606 257352 282611 257408
rect 279926 257350 282611 257352
rect 227294 257002 227300 257004
rect 110462 256942 227300 257002
rect 110462 256934 110522 256942
rect 227294 256940 227300 256942
rect 227364 256940 227370 257004
rect 279926 256972 279986 257350
rect 282545 257347 282611 257350
rect 109940 256874 110522 256934
rect 178677 256866 178743 256869
rect 178677 256864 239690 256866
rect 178677 256808 178682 256864
rect 178738 256808 239690 256864
rect 178677 256806 239690 256808
rect 178677 256803 178743 256806
rect 239630 256798 239690 256806
rect 239630 256738 240212 256798
rect 226558 256668 226564 256732
rect 226628 256730 226634 256732
rect 227529 256730 227595 256733
rect 226628 256728 227595 256730
rect 226628 256672 227534 256728
rect 227590 256672 227595 256728
rect 226628 256670 227595 256672
rect 226628 256668 226634 256670
rect 227529 256667 227595 256670
rect 282821 256458 282887 256461
rect 279926 256456 282887 256458
rect 279926 256400 282826 256456
rect 282882 256400 282887 256456
rect 279926 256398 282887 256400
rect 279926 256156 279986 256398
rect 282821 256395 282887 256398
rect 280153 256050 280219 256053
rect 279926 256048 280219 256050
rect 279926 255992 280158 256048
rect 280214 255992 280219 256048
rect 279926 255990 280219 255992
rect 239630 255650 240212 255710
rect 238109 255642 238175 255645
rect 239630 255642 239690 255650
rect 238109 255640 239690 255642
rect 238109 255584 238114 255640
rect 238170 255584 239690 255640
rect 238109 255582 239690 255584
rect 238109 255579 238175 255582
rect 224902 255370 224908 255372
rect 110094 255310 224908 255370
rect 110094 255302 110154 255310
rect 224902 255308 224908 255310
rect 224972 255308 224978 255372
rect 279926 255340 279986 255990
rect 280153 255987 280219 255990
rect 109940 255242 110154 255302
rect 283005 255098 283071 255101
rect 279926 255096 283071 255098
rect 279926 255040 283010 255096
rect 283066 255040 283071 255096
rect 279926 255038 283071 255040
rect 123477 254690 123543 254693
rect 123477 254688 239690 254690
rect 123477 254632 123482 254688
rect 123538 254632 239690 254688
rect 123477 254630 239690 254632
rect 123477 254627 123543 254630
rect 239630 254622 239690 254630
rect 239630 254562 240212 254622
rect 279926 254524 279986 255038
rect 283005 255035 283071 255038
rect -960 254146 480 254236
rect 48630 254146 48636 254148
rect -960 254086 48636 254146
rect -960 253996 480 254086
rect 48630 254084 48636 254086
rect 48700 254084 48706 254148
rect 287094 253874 287100 253876
rect 279926 253814 287100 253874
rect 227110 253738 227116 253740
rect 110462 253678 227116 253738
rect 110462 253670 110522 253678
rect 227110 253676 227116 253678
rect 227180 253676 227186 253740
rect 279926 253708 279986 253814
rect 287094 253812 287100 253814
rect 287164 253812 287170 253876
rect 109940 253610 110522 253670
rect 197997 253602 198063 253605
rect 197997 253600 239690 253602
rect 197997 253544 198002 253600
rect 198058 253544 239690 253600
rect 197997 253542 239690 253544
rect 197997 253539 198063 253542
rect 239630 253534 239690 253542
rect 239630 253474 240212 253534
rect 282821 253466 282887 253469
rect 279926 253464 282887 253466
rect 279926 253408 282826 253464
rect 282882 253408 282887 253464
rect 279926 253406 282887 253408
rect 279926 252892 279986 253406
rect 282821 253403 282887 253406
rect 451917 253194 451983 253197
rect 454677 253194 454743 253197
rect 451917 253192 454743 253194
rect 451917 253136 451922 253192
rect 451978 253136 454682 253192
rect 454738 253136 454743 253192
rect 451917 253134 454743 253136
rect 451917 253131 451983 253134
rect 454677 253131 454743 253134
rect 116393 252514 116459 252517
rect 116393 252512 239690 252514
rect 116393 252456 116398 252512
rect 116454 252456 239690 252512
rect 116393 252454 239690 252456
rect 116393 252451 116459 252454
rect 239630 252446 239690 252454
rect 239630 252386 240212 252446
rect 226190 252106 226196 252108
rect 110462 252046 226196 252106
rect 110462 252038 110522 252046
rect 226190 252044 226196 252046
rect 226260 252044 226266 252108
rect 292614 252106 292620 252108
rect 109940 251978 110522 252038
rect 279926 251970 279986 252076
rect 282870 252046 292620 252106
rect 282870 251970 282930 252046
rect 292614 252044 292620 252046
rect 292684 252044 292690 252108
rect 279926 251910 282930 251970
rect 228909 251426 228975 251429
rect 228909 251424 239690 251426
rect 228909 251368 228914 251424
rect 228970 251368 239690 251424
rect 228909 251366 239690 251368
rect 228909 251363 228975 251366
rect 239630 251358 239690 251366
rect 279926 251366 282930 251426
rect 239630 251298 240212 251358
rect 279926 251260 279986 251366
rect 282870 251290 282930 251366
rect 292665 251290 292731 251293
rect 282870 251288 292731 251290
rect 282870 251232 292670 251288
rect 292726 251232 292731 251288
rect 282870 251230 292731 251232
rect 292665 251227 292731 251230
rect 230054 250474 230060 250476
rect 110462 250414 230060 250474
rect 110462 250406 110522 250414
rect 230054 250412 230060 250414
rect 230124 250412 230130 250476
rect 109940 250346 110522 250406
rect 163497 250338 163563 250341
rect 279926 250338 279986 250444
rect 290089 250338 290155 250341
rect 163497 250336 239690 250338
rect 163497 250280 163502 250336
rect 163558 250280 239690 250336
rect 163497 250278 239690 250280
rect 279926 250336 290155 250338
rect 279926 250280 290094 250336
rect 290150 250280 290155 250336
rect 279926 250278 290155 250280
rect 163497 250275 163563 250278
rect 239630 250270 239690 250278
rect 290089 250275 290155 250278
rect 239630 250210 240212 250270
rect 279926 249522 279986 249628
rect 290181 249522 290247 249525
rect 279926 249520 290247 249522
rect 279926 249464 290186 249520
rect 290242 249464 290247 249520
rect 279926 249462 290247 249464
rect 290181 249459 290247 249462
rect 202137 249250 202203 249253
rect 202137 249248 239690 249250
rect 202137 249192 202142 249248
rect 202198 249192 239690 249248
rect 202137 249190 239690 249192
rect 202137 249187 202203 249190
rect 239630 249182 239690 249190
rect 239630 249122 240212 249182
rect 229870 248842 229876 248844
rect 110462 248782 229876 248842
rect 110462 248774 110522 248782
rect 229870 248780 229876 248782
rect 229940 248780 229946 248844
rect 109940 248714 110522 248774
rect 279926 248706 279986 248812
rect 285806 248706 285812 248708
rect 279926 248646 285812 248706
rect 285806 248644 285812 248646
rect 285876 248644 285882 248708
rect 209037 248162 209103 248165
rect 209037 248160 239690 248162
rect 209037 248104 209042 248160
rect 209098 248104 239690 248160
rect 209037 248102 239690 248104
rect 209037 248099 209103 248102
rect 239630 248094 239690 248102
rect 239630 248034 240212 248094
rect 279926 247890 279986 247996
rect 290273 247890 290339 247893
rect 279926 247888 290339 247890
rect 279926 247832 290278 247888
rect 290334 247832 290339 247888
rect 279926 247830 290339 247832
rect 290273 247827 290339 247830
rect 228214 247210 228220 247212
rect 110462 247150 228220 247210
rect 110462 247142 110522 247150
rect 228214 247148 228220 247150
rect 228284 247148 228290 247212
rect 109940 247082 110522 247142
rect 279926 247074 279986 247180
rect 291653 247074 291719 247077
rect 279926 247072 291719 247074
rect 279926 247016 291658 247072
rect 291714 247016 291719 247072
rect 279926 247014 291719 247016
rect 291653 247011 291719 247014
rect 239630 246946 240212 247006
rect 226977 246938 227043 246941
rect 239630 246938 239690 246946
rect 226977 246936 239690 246938
rect 226977 246880 226982 246936
rect 227038 246880 239690 246936
rect 226977 246878 239690 246880
rect 226977 246875 227043 246878
rect 279926 246258 279986 246364
rect 288382 246258 288388 246260
rect 279926 246198 288388 246258
rect 288382 246196 288388 246198
rect 288452 246196 288458 246260
rect 216029 245986 216095 245989
rect 216029 245984 239690 245986
rect 216029 245928 216034 245984
rect 216090 245928 239690 245984
rect 216029 245926 239690 245928
rect 216029 245923 216095 245926
rect 239630 245918 239690 245926
rect 239630 245858 240212 245918
rect 113817 245714 113883 245717
rect 114645 245714 114711 245717
rect 113817 245712 114711 245714
rect 113817 245656 113822 245712
rect 113878 245656 114650 245712
rect 114706 245656 114711 245712
rect 113817 245654 114711 245656
rect 113817 245651 113883 245654
rect 114645 245651 114711 245654
rect 231158 245578 231164 245580
rect 110462 245518 231164 245578
rect 110462 245510 110522 245518
rect 231158 245516 231164 245518
rect 231228 245516 231234 245580
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 109940 245450 110522 245510
rect 279926 245442 279986 245548
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 291326 245442 291332 245444
rect 279926 245382 291332 245442
rect 291326 245380 291332 245382
rect 291396 245380 291402 245444
rect 583520 245428 584960 245518
rect 48078 244972 48084 245036
rect 48148 245034 48154 245036
rect 48148 244974 50140 245034
rect 48148 244972 48154 244974
rect 211797 244898 211863 244901
rect 211797 244896 239690 244898
rect 211797 244840 211802 244896
rect 211858 244840 239690 244896
rect 211797 244838 239690 244840
rect 211797 244835 211863 244838
rect 239630 244830 239690 244838
rect 239630 244770 240212 244830
rect 279926 244626 279986 244732
rect 291142 244626 291148 244628
rect 279926 244566 291148 244626
rect 291142 244564 291148 244566
rect 291212 244564 291218 244628
rect 224534 243946 224540 243948
rect 110462 243886 224540 243946
rect 110462 243878 110522 243886
rect 224534 243884 224540 243886
rect 224604 243884 224610 243948
rect 291510 243946 291516 243948
rect 109940 243818 110522 243878
rect 126237 243810 126303 243813
rect 279926 243810 279986 243916
rect 287010 243886 291516 243946
rect 287010 243810 287070 243886
rect 291510 243884 291516 243886
rect 291580 243884 291586 243948
rect 126237 243808 239690 243810
rect 126237 243752 126242 243808
rect 126298 243752 239690 243808
rect 126237 243750 239690 243752
rect 279926 243750 287070 243810
rect 126237 243747 126303 243750
rect 239630 243742 239690 243750
rect 239630 243682 240212 243742
rect 279926 242994 279986 243100
rect 282821 242994 282887 242997
rect 279926 242992 282887 242994
rect 279926 242936 282826 242992
rect 282882 242936 282887 242992
rect 279926 242934 282887 242936
rect 282821 242931 282887 242934
rect 188337 242722 188403 242725
rect 188337 242720 239690 242722
rect 188337 242664 188342 242720
rect 188398 242664 239690 242720
rect 188337 242662 239690 242664
rect 188337 242659 188403 242662
rect 239630 242654 239690 242662
rect 239630 242594 240212 242654
rect 233734 242314 233740 242316
rect 110462 242254 233740 242314
rect 110462 242246 110522 242254
rect 233734 242252 233740 242254
rect 233804 242252 233810 242316
rect 288566 242314 288572 242316
rect 109940 242186 110522 242246
rect 279926 242178 279986 242284
rect 287010 242254 288572 242314
rect 287010 242178 287070 242254
rect 288566 242252 288572 242254
rect 288636 242252 288642 242316
rect 279926 242118 287070 242178
rect 239814 241506 240212 241566
rect 210417 241498 210483 241501
rect 239814 241498 239874 241506
rect 290774 241498 290780 241500
rect 210417 241496 239874 241498
rect 210417 241440 210422 241496
rect 210478 241440 239874 241496
rect 210417 241438 239874 241440
rect 210417 241435 210483 241438
rect 279926 241362 279986 241468
rect 287010 241438 290780 241498
rect 287010 241362 287070 241438
rect 290774 241436 290780 241438
rect 290844 241436 290850 241500
rect 279926 241302 287070 241362
rect -960 241090 480 241180
rect 3366 241090 3372 241092
rect -960 241030 3372 241090
rect -960 240940 480 241030
rect 3366 241028 3372 241030
rect 3436 241028 3442 241092
rect 223246 240682 223252 240684
rect 110462 240622 223252 240682
rect 110462 240614 110522 240622
rect 223246 240620 223252 240622
rect 223316 240620 223322 240684
rect 290365 240682 290431 240685
rect 287010 240680 290431 240682
rect 109940 240554 110522 240614
rect 142797 240546 142863 240549
rect 279926 240546 279986 240652
rect 287010 240624 290370 240680
rect 290426 240624 290431 240680
rect 287010 240622 290431 240624
rect 287010 240546 287070 240622
rect 290365 240619 290431 240622
rect 142797 240544 239690 240546
rect 142797 240488 142802 240544
rect 142858 240488 239690 240544
rect 142797 240486 239690 240488
rect 279926 240486 287070 240546
rect 142797 240483 142863 240486
rect 239630 240478 239690 240486
rect 239630 240418 240212 240478
rect 114645 240138 114711 240141
rect 116577 240138 116643 240141
rect 114645 240136 116643 240138
rect 114645 240080 114650 240136
rect 114706 240080 116582 240136
rect 116638 240080 116643 240136
rect 114645 240078 116643 240080
rect 114645 240075 114711 240078
rect 116577 240075 116643 240078
rect 151077 239458 151143 239461
rect 151077 239456 239690 239458
rect 151077 239400 151082 239456
rect 151138 239400 239690 239456
rect 151077 239398 239690 239400
rect 151077 239395 151143 239398
rect 239630 239390 239690 239398
rect 239630 239330 240212 239390
rect 279926 239322 279986 239836
rect 281533 239322 281599 239325
rect 279926 239320 281599 239322
rect 279926 239264 281538 239320
rect 281594 239264 281599 239320
rect 279926 239262 281599 239264
rect 281533 239259 281599 239262
rect 223062 239050 223068 239052
rect 110462 238990 223068 239050
rect 110462 238982 110522 238990
rect 223062 238988 223068 238990
rect 223132 238988 223138 239052
rect 109940 238922 110522 238982
rect 279926 238914 279986 239020
rect 285857 238914 285923 238917
rect 279926 238912 285923 238914
rect 279926 238856 285862 238912
rect 285918 238856 285923 238912
rect 279926 238854 285923 238856
rect 285857 238851 285923 238854
rect 440877 238778 440943 238781
rect 442257 238778 442323 238781
rect 440877 238776 442323 238778
rect 440877 238720 440882 238776
rect 440938 238720 442262 238776
rect 442318 238720 442323 238776
rect 440877 238718 442323 238720
rect 440877 238715 440943 238718
rect 442257 238715 442323 238718
rect 214557 238370 214623 238373
rect 214557 238368 239690 238370
rect 214557 238312 214562 238368
rect 214618 238312 239690 238368
rect 214557 238310 239690 238312
rect 214557 238307 214623 238310
rect 239630 238302 239690 238310
rect 239630 238242 240212 238302
rect 279926 237690 279986 238204
rect 281809 237690 281875 237693
rect 279926 237688 281875 237690
rect 279926 237632 281814 237688
rect 281870 237632 281875 237688
rect 279926 237630 281875 237632
rect 281809 237627 281875 237630
rect 279926 237494 280170 237554
rect 222878 237418 222884 237420
rect 110094 237358 222884 237418
rect 110094 237350 110154 237358
rect 222878 237356 222884 237358
rect 222948 237356 222954 237420
rect 279926 237388 279986 237494
rect 280110 237421 280170 237494
rect 280110 237416 280219 237421
rect 280110 237360 280158 237416
rect 280214 237360 280219 237416
rect 280110 237358 280219 237360
rect 280153 237355 280219 237358
rect 109940 237290 110154 237350
rect 140037 237282 140103 237285
rect 140037 237280 239690 237282
rect 140037 237224 140042 237280
rect 140098 237224 239690 237280
rect 140037 237222 239690 237224
rect 140037 237219 140103 237222
rect 239630 237214 239690 237222
rect 239630 237154 240212 237214
rect 231117 236194 231183 236197
rect 231117 236192 239690 236194
rect 231117 236136 231122 236192
rect 231178 236136 239690 236192
rect 231117 236134 239690 236136
rect 231117 236131 231183 236134
rect 239630 236126 239690 236134
rect 239630 236066 240212 236126
rect 279926 236058 279986 236572
rect 280337 236058 280403 236061
rect 279926 236056 280403 236058
rect 279926 236000 280342 236056
rect 280398 236000 280403 236056
rect 279926 235998 280403 236000
rect 280337 235995 280403 235998
rect 222694 235786 222700 235788
rect 110462 235726 222700 235786
rect 110462 235718 110522 235726
rect 222694 235724 222700 235726
rect 222764 235724 222770 235788
rect 109940 235658 110522 235718
rect 279926 235242 279986 235756
rect 281717 235242 281783 235245
rect 279926 235240 281783 235242
rect 279926 235184 281722 235240
rect 281778 235184 281783 235240
rect 279926 235182 281783 235184
rect 281717 235179 281783 235182
rect 199377 235106 199443 235109
rect 199377 235104 239690 235106
rect 199377 235048 199382 235104
rect 199438 235048 239690 235104
rect 199377 235046 239690 235048
rect 199377 235043 199443 235046
rect 239630 235038 239690 235046
rect 239630 234978 240212 235038
rect 279926 234698 279986 234940
rect 280245 234698 280311 234701
rect 279926 234696 280311 234698
rect 279926 234640 280250 234696
rect 280306 234640 280311 234696
rect 279926 234638 280311 234640
rect 280245 234635 280311 234638
rect 226926 234154 226932 234156
rect 110462 234094 226932 234154
rect 110462 234086 110522 234094
rect 226926 234092 226932 234094
rect 226996 234092 227002 234156
rect 109940 234026 110522 234086
rect 146937 234018 147003 234021
rect 146937 234016 239690 234018
rect 146937 233960 146942 234016
rect 146998 233960 239690 234016
rect 146937 233958 239690 233960
rect 146937 233955 147003 233958
rect 239630 233950 239690 233958
rect 239630 233890 240212 233950
rect 279926 233610 279986 234124
rect 281625 233610 281691 233613
rect 279926 233608 281691 233610
rect 279926 233552 281630 233608
rect 281686 233552 281691 233608
rect 279926 233550 281691 233552
rect 281625 233547 281691 233550
rect 279926 233414 280170 233474
rect 279926 233308 279986 233414
rect 280110 233338 280170 233414
rect 281993 233338 282059 233341
rect 280110 233336 282059 233338
rect 280110 233280 281998 233336
rect 282054 233280 282059 233336
rect 280110 233278 282059 233280
rect 281993 233275 282059 233278
rect 174537 232930 174603 232933
rect 174537 232928 239690 232930
rect 174537 232872 174542 232928
rect 174598 232872 239690 232928
rect 174537 232870 239690 232872
rect 174537 232867 174603 232870
rect 239630 232862 239690 232870
rect 239630 232802 240212 232862
rect 224350 232522 224356 232524
rect 110462 232462 224356 232522
rect 110462 232454 110522 232462
rect 224350 232460 224356 232462
rect 224420 232460 224426 232524
rect 109940 232394 110522 232454
rect 279926 231978 279986 232492
rect 580349 232386 580415 232389
rect 583520 232386 584960 232476
rect 580349 232384 584960 232386
rect 580349 232328 580354 232384
rect 580410 232328 584960 232384
rect 580349 232326 584960 232328
rect 580349 232323 580415 232326
rect 583520 232236 584960 232326
rect 285949 231978 286015 231981
rect 279926 231976 286015 231978
rect 279926 231920 285954 231976
rect 286010 231920 286015 231976
rect 279926 231918 286015 231920
rect 285949 231915 286015 231918
rect 138657 231842 138723 231845
rect 439497 231842 439563 231845
rect 440877 231842 440943 231845
rect 138657 231840 239690 231842
rect 138657 231784 138662 231840
rect 138718 231784 239690 231840
rect 138657 231782 239690 231784
rect 138657 231779 138723 231782
rect 239630 231774 239690 231782
rect 439497 231840 440943 231842
rect 439497 231784 439502 231840
rect 439558 231784 440882 231840
rect 440938 231784 440943 231840
rect 439497 231782 440943 231784
rect 439497 231779 439563 231782
rect 440877 231779 440943 231782
rect 239630 231714 240212 231774
rect 279926 231162 279986 231676
rect 281901 231162 281967 231165
rect 279926 231160 281967 231162
rect 279926 231104 281906 231160
rect 281962 231104 281967 231160
rect 279926 231102 281967 231104
rect 281901 231099 281967 231102
rect 226558 230890 226564 230892
rect 110462 230830 226564 230890
rect 110462 230822 110522 230830
rect 226558 230828 226564 230830
rect 226628 230828 226634 230892
rect 109940 230762 110522 230822
rect 191097 230754 191163 230757
rect 191097 230752 239690 230754
rect 191097 230696 191102 230752
rect 191158 230696 239690 230752
rect 191097 230694 239690 230696
rect 191097 230691 191163 230694
rect 239630 230686 239690 230694
rect 239630 230626 240212 230686
rect 279926 230618 279986 230860
rect 283097 230618 283163 230621
rect 279926 230616 283163 230618
rect 279926 230560 283102 230616
rect 283158 230560 283163 230616
rect 279926 230558 283163 230560
rect 283097 230555 283163 230558
rect 152457 229666 152523 229669
rect 152457 229664 239690 229666
rect 152457 229608 152462 229664
rect 152518 229608 239690 229664
rect 152457 229606 239690 229608
rect 152457 229603 152523 229606
rect 239630 229598 239690 229606
rect 239630 229538 240212 229598
rect 279926 229530 279986 230044
rect 284477 229530 284543 229533
rect 279926 229528 284543 229530
rect 279926 229472 284482 229528
rect 284538 229472 284543 229528
rect 279926 229470 284543 229472
rect 284477 229467 284543 229470
rect 226374 229258 226380 229260
rect 110462 229198 226380 229258
rect 110462 229190 110522 229198
rect 226374 229196 226380 229198
rect 226444 229196 226450 229260
rect 282177 229258 282243 229261
rect 280110 229256 282243 229258
rect 109940 229130 110522 229190
rect 279926 229122 279986 229228
rect 280110 229200 282182 229256
rect 282238 229200 282243 229256
rect 280110 229198 282243 229200
rect 280110 229122 280170 229198
rect 282177 229195 282243 229198
rect 279926 229062 280170 229122
rect 144177 228578 144243 228581
rect 144177 228576 239690 228578
rect 144177 228520 144182 228576
rect 144238 228520 239690 228576
rect 144177 228518 239690 228520
rect 144177 228515 144243 228518
rect 239630 228510 239690 228518
rect 239630 228450 240212 228510
rect -960 227884 480 228124
rect 279926 227898 279986 228412
rect 282269 227898 282335 227901
rect 279926 227896 282335 227898
rect 279926 227840 282274 227896
rect 282330 227840 282335 227896
rect 279926 227838 282335 227840
rect 282269 227835 282335 227838
rect 232262 227626 232268 227628
rect 110462 227566 232268 227626
rect 110462 227558 110522 227566
rect 232262 227564 232268 227566
rect 232332 227564 232338 227628
rect 109940 227498 110522 227558
rect 155217 227490 155283 227493
rect 155217 227488 239690 227490
rect 155217 227432 155222 227488
rect 155278 227432 239690 227488
rect 155217 227430 239690 227432
rect 155217 227427 155283 227430
rect 239630 227422 239690 227430
rect 239630 227362 240212 227422
rect 279926 227082 279986 227596
rect 284661 227082 284727 227085
rect 279926 227080 284727 227082
rect 279926 227024 284666 227080
rect 284722 227024 284727 227080
rect 279926 227022 284727 227024
rect 284661 227019 284727 227022
rect 279926 226402 279986 226780
rect 284753 226402 284819 226405
rect 279926 226400 284819 226402
rect 279926 226344 284758 226400
rect 284814 226344 284819 226400
rect 279926 226342 284819 226344
rect 284753 226339 284819 226342
rect 239630 226274 240212 226334
rect 223297 226266 223363 226269
rect 239630 226266 239690 226274
rect 223297 226264 239690 226266
rect 223297 226208 223302 226264
rect 223358 226208 239690 226264
rect 223297 226206 239690 226208
rect 223297 226203 223363 226206
rect 224166 225994 224172 225996
rect 110462 225934 224172 225994
rect 110462 225926 110522 225934
rect 224166 225932 224172 225934
rect 224236 225932 224242 225996
rect 109940 225866 110522 225926
rect 279926 225450 279986 225964
rect 279926 225390 280170 225450
rect 280110 225314 280170 225390
rect 282085 225314 282151 225317
rect 280110 225312 282151 225314
rect 280110 225256 282090 225312
rect 282146 225256 282151 225312
rect 280110 225254 282151 225256
rect 282085 225251 282151 225254
rect 239630 225186 240212 225246
rect 238017 225178 238083 225181
rect 239630 225178 239690 225186
rect 238017 225176 239690 225178
rect 238017 225120 238022 225176
rect 238078 225120 239690 225176
rect 238017 225118 239690 225120
rect 238017 225115 238083 225118
rect 279926 225042 279986 225148
rect 280521 225042 280587 225045
rect 279926 225040 280587 225042
rect 279926 224984 280526 225040
rect 280582 224984 280587 225040
rect 279926 224982 280587 224984
rect 280521 224979 280587 224982
rect 450537 224906 450603 224909
rect 451917 224906 451983 224909
rect 450537 224904 451983 224906
rect 450537 224848 450542 224904
rect 450598 224848 451922 224904
rect 451978 224848 451983 224904
rect 450537 224846 451983 224848
rect 450537 224843 450603 224846
rect 451917 224843 451983 224846
rect 232078 224362 232084 224364
rect 110462 224302 232084 224362
rect 110462 224294 110522 224302
rect 232078 224300 232084 224302
rect 232148 224300 232154 224364
rect 109940 224234 110522 224294
rect 116577 224226 116643 224229
rect 120717 224226 120783 224229
rect 116577 224224 120783 224226
rect 116577 224168 116582 224224
rect 116638 224168 120722 224224
rect 120778 224168 120783 224224
rect 116577 224166 120783 224168
rect 116577 224163 116643 224166
rect 120717 224163 120783 224166
rect 206277 224226 206343 224229
rect 206277 224224 239690 224226
rect 206277 224168 206282 224224
rect 206338 224168 239690 224224
rect 206277 224166 239690 224168
rect 206277 224163 206343 224166
rect 239630 224158 239690 224166
rect 239630 224098 240212 224158
rect 279926 223818 279986 224332
rect 279926 223758 280170 223818
rect 280110 223682 280170 223758
rect 284845 223682 284911 223685
rect 280110 223680 284911 223682
rect 280110 223624 284850 223680
rect 284906 223624 284911 223680
rect 280110 223622 284911 223624
rect 284845 223619 284911 223622
rect 215937 223138 216003 223141
rect 215937 223136 239690 223138
rect 215937 223080 215942 223136
rect 215998 223080 239690 223136
rect 215937 223078 239690 223080
rect 215937 223075 216003 223078
rect 239630 223070 239690 223078
rect 239630 223010 240212 223070
rect 279926 223002 279986 223516
rect 279926 222942 280170 223002
rect 280110 222866 280170 222942
rect 280429 222866 280495 222869
rect 280110 222864 280495 222866
rect 280110 222808 280434 222864
rect 280490 222808 280495 222864
rect 280110 222806 280495 222808
rect 280429 222803 280495 222806
rect 232589 222730 232655 222733
rect 110462 222728 232655 222730
rect 110462 222672 232594 222728
rect 232650 222672 232655 222728
rect 110462 222670 232655 222672
rect 110462 222662 110522 222670
rect 232589 222667 232655 222670
rect 109940 222602 110522 222662
rect 279926 222322 279986 222700
rect 283281 222322 283347 222325
rect 279926 222320 283347 222322
rect 279926 222264 283286 222320
rect 283342 222264 283347 222320
rect 279926 222262 283347 222264
rect 283281 222259 283347 222262
rect 203517 222050 203583 222053
rect 203517 222048 239690 222050
rect 203517 221992 203522 222048
rect 203578 221992 239690 222048
rect 203517 221990 239690 221992
rect 203517 221987 203583 221990
rect 239630 221982 239690 221990
rect 239630 221922 240212 221982
rect 279926 221370 279986 221884
rect 283373 221370 283439 221373
rect 279926 221368 283439 221370
rect 279926 221312 283378 221368
rect 283434 221312 283439 221368
rect 279926 221310 283439 221312
rect 283373 221307 283439 221310
rect 232497 221098 232563 221101
rect 110462 221096 232563 221098
rect 110462 221040 232502 221096
rect 232558 221040 232563 221096
rect 110462 221038 232563 221040
rect 110462 221030 110522 221038
rect 232497 221035 232563 221038
rect 109940 220970 110522 221030
rect 279926 220962 279986 221068
rect 282177 220962 282243 220965
rect 279926 220960 282243 220962
rect 279926 220904 282182 220960
rect 282238 220904 282243 220960
rect 279926 220902 282243 220904
rect 282177 220899 282243 220902
rect 239814 220834 240212 220894
rect 195237 220826 195303 220829
rect 239814 220826 239874 220834
rect 195237 220824 239874 220826
rect 195237 220768 195242 220824
rect 195298 220768 239874 220824
rect 195237 220766 239874 220768
rect 195237 220763 195303 220766
rect 213177 219874 213243 219877
rect 279926 219874 279986 220252
rect 282453 219874 282519 219877
rect 213177 219872 239690 219874
rect 213177 219816 213182 219872
rect 213238 219816 239690 219872
rect 213177 219814 239690 219816
rect 279926 219872 282519 219874
rect 279926 219816 282458 219872
rect 282514 219816 282519 219872
rect 279926 219814 282519 219816
rect 213177 219811 213243 219814
rect 239630 219806 239690 219814
rect 282453 219811 282519 219814
rect 239630 219746 240212 219806
rect 232681 219466 232747 219469
rect 282821 219466 282887 219469
rect 110094 219464 232747 219466
rect 110094 219408 232686 219464
rect 232742 219408 232747 219464
rect 280110 219464 282887 219466
rect 280110 219450 282826 219464
rect 110094 219406 232747 219408
rect 110094 219398 110154 219406
rect 232681 219403 232747 219406
rect 279926 219408 282826 219450
rect 282882 219408 282887 219464
rect 279926 219406 282887 219408
rect 109940 219338 110154 219398
rect 279926 219390 280170 219406
rect 282821 219403 282887 219406
rect 580206 218996 580212 219060
rect 580276 219058 580282 219060
rect 583520 219058 584960 219148
rect 580276 218998 584960 219058
rect 580276 218996 580282 218998
rect 583520 218908 584960 218998
rect 158713 218786 158779 218789
rect 158713 218784 239690 218786
rect 158713 218728 158718 218784
rect 158774 218728 239690 218784
rect 158713 218726 239690 218728
rect 158713 218723 158779 218726
rect 239630 218718 239690 218726
rect 239806 218718 239812 218720
rect 239630 218658 239812 218718
rect 239806 218656 239812 218658
rect 239876 218718 239882 218720
rect 239876 218658 240212 218718
rect 239876 218656 239882 218658
rect 279926 218106 279986 218620
rect 282361 218106 282427 218109
rect 279926 218104 282427 218106
rect 279926 218048 282366 218104
rect 282422 218048 282427 218104
rect 279926 218046 282427 218048
rect 282361 218043 282427 218046
rect 238334 217834 238340 217836
rect 110462 217774 238340 217834
rect 110462 217766 110522 217774
rect 238334 217772 238340 217774
rect 238404 217772 238410 217836
rect 288433 217834 288499 217837
rect 287010 217832 288499 217834
rect 109940 217706 110522 217766
rect 224166 217636 224172 217700
rect 224236 217698 224242 217700
rect 279926 217698 279986 217804
rect 287010 217776 288438 217832
rect 288494 217776 288499 217832
rect 287010 217774 288499 217776
rect 287010 217698 287070 217774
rect 288433 217771 288499 217774
rect 224236 217638 239690 217698
rect 279926 217638 287070 217698
rect 224236 217636 224242 217638
rect 239630 217630 239690 217638
rect 239630 217570 240212 217630
rect 279926 216882 279986 216988
rect 279926 216822 282194 216882
rect 237414 216684 237420 216748
rect 237484 216746 237490 216748
rect 238661 216746 238727 216749
rect 237484 216744 238727 216746
rect 237484 216688 238666 216744
rect 238722 216688 238727 216744
rect 237484 216686 238727 216688
rect 237484 216684 237490 216686
rect 238661 216683 238727 216686
rect 280797 216746 280863 216749
rect 281901 216746 281967 216749
rect 280797 216744 281967 216746
rect 280797 216688 280802 216744
rect 280858 216688 281906 216744
rect 281962 216688 281967 216744
rect 280797 216686 281967 216688
rect 282134 216746 282194 216822
rect 283465 216746 283531 216749
rect 282134 216744 283531 216746
rect 282134 216688 283470 216744
rect 283526 216688 283531 216744
rect 282134 216686 283531 216688
rect 280797 216683 280863 216686
rect 281901 216683 281967 216686
rect 283465 216683 283531 216686
rect 219934 216548 219940 216612
rect 220004 216610 220010 216612
rect 220004 216550 239690 216610
rect 220004 216548 220010 216550
rect 239630 216542 239690 216550
rect 239630 216482 240212 216542
rect 232773 216202 232839 216205
rect 110462 216200 232839 216202
rect 110462 216144 232778 216200
rect 232834 216144 232839 216200
rect 110462 216142 232839 216144
rect 110462 216134 110522 216142
rect 232773 216139 232839 216142
rect 109940 216074 110522 216134
rect 279926 215658 279986 216172
rect 283557 215658 283623 215661
rect 279926 215656 283623 215658
rect 279926 215600 283562 215656
rect 283618 215600 283623 215656
rect 279926 215598 283623 215600
rect 283557 215595 283623 215598
rect 228214 215460 228220 215524
rect 228284 215522 228290 215524
rect 228284 215462 239690 215522
rect 228284 215460 228290 215462
rect 239630 215454 239690 215462
rect 279926 215462 280170 215522
rect 239630 215394 240212 215454
rect 279926 215356 279986 215462
rect 280110 215386 280170 215462
rect 284385 215386 284451 215389
rect 280110 215384 284451 215386
rect 280110 215328 284390 215384
rect 284446 215328 284451 215384
rect 280110 215326 284451 215328
rect 284385 215323 284451 215326
rect 48221 215114 48287 215117
rect 48221 215112 50140 215114
rect -960 214978 480 215068
rect 48221 215056 48226 215112
rect 48282 215056 50140 215112
rect 48221 215054 50140 215056
rect 48221 215051 48287 215054
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 232957 214570 233023 214573
rect 110462 214568 233023 214570
rect 110462 214512 232962 214568
rect 233018 214512 233023 214568
rect 110462 214510 233023 214512
rect 110462 214502 110522 214510
rect 232957 214507 233023 214510
rect 109940 214442 110522 214502
rect 239630 214306 240212 214366
rect 237373 214298 237439 214301
rect 239630 214298 239690 214306
rect 237373 214296 239690 214298
rect 237373 214240 237378 214296
rect 237434 214240 239690 214296
rect 237373 214238 239690 214240
rect 237373 214235 237439 214238
rect 279926 214026 279986 214540
rect 283189 214026 283255 214029
rect 279926 214024 283255 214026
rect 279926 213968 283194 214024
rect 283250 213968 283255 214024
rect 279926 213966 283255 213968
rect 283189 213963 283255 213966
rect 231158 213284 231164 213348
rect 231228 213346 231234 213348
rect 231228 213286 239690 213346
rect 231228 213284 231234 213286
rect 239630 213278 239690 213286
rect 239630 213218 240212 213278
rect 279926 213210 279986 213724
rect 280613 213210 280679 213213
rect 279926 213208 280679 213210
rect 279926 213152 280618 213208
rect 280674 213152 280679 213208
rect 279926 213150 280679 213152
rect 280613 213147 280679 213150
rect 235206 212938 235212 212940
rect 110462 212878 235212 212938
rect 110462 212870 110522 212878
rect 235206 212876 235212 212878
rect 235276 212876 235282 212940
rect 109940 212810 110522 212870
rect 279926 212666 279986 212908
rect 281901 212666 281967 212669
rect 279926 212664 281967 212666
rect 279926 212608 281906 212664
rect 281962 212608 281967 212664
rect 279926 212606 281967 212608
rect 281901 212603 281967 212606
rect 116526 212196 116532 212260
rect 116596 212258 116602 212260
rect 116596 212198 239690 212258
rect 116596 212196 116602 212198
rect 239630 212190 239690 212198
rect 239630 212130 240212 212190
rect 279926 211714 279986 212092
rect 282821 211714 282887 211717
rect 279926 211712 282887 211714
rect 279926 211656 282826 211712
rect 282882 211656 282887 211712
rect 279926 211654 282887 211656
rect 282821 211651 282887 211654
rect 235390 211306 235396 211308
rect 110462 211246 235396 211306
rect 110462 211238 110522 211246
rect 235390 211244 235396 211246
rect 235460 211244 235466 211308
rect 109940 211178 110522 211238
rect 121453 211170 121519 211173
rect 123569 211170 123635 211173
rect 121453 211168 123635 211170
rect 121453 211112 121458 211168
rect 121514 211112 123574 211168
rect 123630 211112 123635 211168
rect 121453 211110 123635 211112
rect 279926 211170 279986 211276
rect 280838 211244 280844 211308
rect 280908 211244 280914 211308
rect 280846 211170 280906 211244
rect 279926 211110 280906 211170
rect 121453 211107 121519 211110
rect 123569 211107 123635 211110
rect 239630 211042 240212 211102
rect 122046 210972 122052 211036
rect 122116 211034 122122 211036
rect 239630 211034 239690 211042
rect 122116 210974 239690 211034
rect 122116 210972 122122 210974
rect 279926 210354 279986 210460
rect 281758 210428 281764 210492
rect 281828 210428 281834 210492
rect 281766 210354 281826 210428
rect 279926 210294 281826 210354
rect 230974 210020 230980 210084
rect 231044 210082 231050 210084
rect 231044 210022 239690 210082
rect 231044 210020 231050 210022
rect 239630 210014 239690 210022
rect 239630 209954 240212 210014
rect 235574 209674 235580 209676
rect 110462 209614 235580 209674
rect 110462 209606 110522 209614
rect 235574 209612 235580 209614
rect 235644 209612 235650 209676
rect 109940 209546 110522 209606
rect 279926 209130 279986 209644
rect 279926 209070 280170 209130
rect 206134 208932 206140 208996
rect 206204 208994 206210 208996
rect 280110 208994 280170 209070
rect 285029 208994 285095 208997
rect 206204 208934 239690 208994
rect 280110 208992 285095 208994
rect 280110 208936 285034 208992
rect 285090 208936 285095 208992
rect 280110 208934 285095 208936
rect 206204 208932 206210 208934
rect 239630 208926 239690 208934
rect 285029 208931 285095 208934
rect 239630 208866 240212 208926
rect 279926 208722 279986 208828
rect 281942 208796 281948 208860
rect 282012 208796 282018 208860
rect 281950 208722 282010 208796
rect 279926 208662 282010 208722
rect 235022 208042 235028 208044
rect 110462 207982 235028 208042
rect 110462 207974 110522 207982
rect 235022 207980 235028 207982
rect 235092 207980 235098 208044
rect 109940 207914 110522 207974
rect 210366 207844 210372 207908
rect 210436 207906 210442 207908
rect 210436 207846 239690 207906
rect 210436 207844 210442 207846
rect 239630 207838 239690 207846
rect 239630 207778 240212 207838
rect 279926 207498 279986 208012
rect 283649 207498 283715 207501
rect 279926 207496 283715 207498
rect 279926 207440 283654 207496
rect 283710 207440 283715 207496
rect 279926 207438 283715 207440
rect 283649 207435 283715 207438
rect 287513 207226 287579 207229
rect 287010 207224 287579 207226
rect 235533 207090 235599 207093
rect 235758 207090 235764 207092
rect 235533 207088 235764 207090
rect 235533 207032 235538 207088
rect 235594 207032 235764 207088
rect 235533 207030 235764 207032
rect 235533 207027 235599 207030
rect 235758 207028 235764 207030
rect 235828 207028 235834 207092
rect 279926 207090 279986 207196
rect 287010 207168 287518 207224
rect 287574 207168 287579 207224
rect 287010 207166 287579 207168
rect 287010 207090 287070 207166
rect 287513 207163 287579 207166
rect 279926 207030 287070 207090
rect 238518 206756 238524 206820
rect 238588 206818 238594 206820
rect 238588 206758 239690 206818
rect 238588 206756 238594 206758
rect 239630 206750 239690 206758
rect 239630 206690 240212 206750
rect 234889 206410 234955 206413
rect 287421 206410 287487 206413
rect 110462 206408 234955 206410
rect 110462 206352 234894 206408
rect 234950 206352 234955 206408
rect 287010 206408 287487 206410
rect 110462 206350 234955 206352
rect 110462 206342 110522 206350
rect 234889 206347 234955 206350
rect 109940 206282 110522 206342
rect 279926 206274 279986 206380
rect 287010 206352 287426 206408
rect 287482 206352 287487 206408
rect 287010 206350 287487 206352
rect 287010 206274 287070 206350
rect 287421 206347 287487 206350
rect 279926 206214 287070 206274
rect 280981 205730 281047 205733
rect 281993 205730 282059 205733
rect 280981 205728 282059 205730
rect 280981 205672 280986 205728
rect 281042 205672 281998 205728
rect 282054 205672 282059 205728
rect 280981 205670 282059 205672
rect 280981 205667 281047 205670
rect 281993 205667 282059 205670
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 239814 205602 240212 205662
rect 214649 205594 214715 205597
rect 239814 205594 239874 205602
rect 214649 205592 239874 205594
rect 214649 205536 214654 205592
rect 214710 205536 239874 205592
rect 583520 205580 584960 205670
rect 214649 205534 239874 205536
rect 214649 205531 214715 205534
rect 279926 205050 279986 205564
rect 279926 204990 280170 205050
rect 235625 204914 235691 204917
rect 238385 204914 238451 204917
rect 235625 204912 238451 204914
rect 235625 204856 235630 204912
rect 235686 204856 238390 204912
rect 238446 204856 238451 204912
rect 235625 204854 238451 204856
rect 280110 204914 280170 204990
rect 282821 204914 282887 204917
rect 280110 204912 282887 204914
rect 280110 204856 282826 204912
rect 282882 204856 282887 204912
rect 280110 204854 282887 204856
rect 235625 204851 235691 204854
rect 238385 204851 238451 204854
rect 282821 204851 282887 204854
rect 239254 204778 239260 204780
rect 110462 204718 239260 204778
rect 110462 204710 110522 204718
rect 239254 204716 239260 204718
rect 239324 204716 239330 204780
rect 109940 204650 110522 204710
rect 238150 204580 238156 204644
rect 238220 204642 238226 204644
rect 238220 204582 239690 204642
rect 238220 204580 238226 204582
rect 239630 204574 239690 204582
rect 239630 204514 240212 204574
rect 279926 204370 279986 204748
rect 286041 204370 286107 204373
rect 279926 204368 286107 204370
rect 279926 204312 286046 204368
rect 286102 204312 286107 204368
rect 279926 204310 286107 204312
rect 286041 204307 286107 204310
rect 281165 204234 281231 204237
rect 282453 204234 282519 204237
rect 281165 204232 282519 204234
rect 281165 204176 281170 204232
rect 281226 204176 282458 204232
rect 282514 204176 282519 204232
rect 281165 204174 282519 204176
rect 281165 204171 281231 204174
rect 282453 204171 282519 204174
rect 449157 204234 449223 204237
rect 450537 204234 450603 204237
rect 449157 204232 450603 204234
rect 449157 204176 449162 204232
rect 449218 204176 450542 204232
rect 450598 204176 450603 204232
rect 449157 204174 450603 204176
rect 449157 204171 449223 204174
rect 450537 204171 450603 204174
rect 238661 203554 238727 203557
rect 238661 203552 239690 203554
rect 238661 203496 238666 203552
rect 238722 203496 239690 203552
rect 238661 203494 239690 203496
rect 238661 203491 238727 203494
rect 239630 203486 239690 203494
rect 239630 203426 240212 203486
rect 279926 203418 279986 203932
rect 279926 203358 280170 203418
rect 280110 203282 280170 203358
rect 281993 203282 282059 203285
rect 280110 203280 282059 203282
rect 280110 203224 281998 203280
rect 282054 203224 282059 203280
rect 280110 203222 282059 203224
rect 281993 203219 282059 203222
rect 238150 203146 238156 203148
rect 110462 203086 238156 203146
rect 110462 203078 110522 203086
rect 238150 203084 238156 203086
rect 238220 203084 238226 203148
rect 109940 203018 110522 203078
rect 279926 203010 279986 203116
rect 284569 203010 284635 203013
rect 279926 203008 284635 203010
rect 279926 202952 284574 203008
rect 284630 202952 284635 203008
rect 279926 202950 284635 202952
rect 284569 202947 284635 202950
rect 228725 202466 228791 202469
rect 228725 202464 239690 202466
rect 228725 202408 228730 202464
rect 228786 202408 239690 202464
rect 228725 202406 239690 202408
rect 228725 202403 228791 202406
rect 239630 202398 239690 202406
rect 239630 202338 240212 202398
rect -960 201922 480 202012
rect 48446 201922 48452 201924
rect -960 201862 48452 201922
rect -960 201772 480 201862
rect 48446 201860 48452 201862
rect 48516 201860 48522 201924
rect 279926 201786 279986 202300
rect 286317 201786 286383 201789
rect 279926 201784 286383 201786
rect 279926 201728 286322 201784
rect 286378 201728 286383 201784
rect 279926 201726 286383 201728
rect 286317 201723 286383 201726
rect 279926 201590 280170 201650
rect 235257 201514 235323 201517
rect 110094 201512 235323 201514
rect 110094 201456 235262 201512
rect 235318 201456 235323 201512
rect 279926 201484 279986 201590
rect 280110 201517 280170 201590
rect 280061 201512 280170 201517
rect 110094 201454 235323 201456
rect 110094 201446 110154 201454
rect 235257 201451 235323 201454
rect 280061 201456 280066 201512
rect 280122 201456 280170 201512
rect 280061 201454 280170 201456
rect 280061 201451 280127 201454
rect 109940 201386 110154 201446
rect 237373 201378 237439 201381
rect 237373 201376 239690 201378
rect 237373 201320 237378 201376
rect 237434 201320 239690 201376
rect 237373 201318 239690 201320
rect 237373 201315 237439 201318
rect 239630 201310 239690 201318
rect 239630 201250 240212 201310
rect 123569 200698 123635 200701
rect 219433 200698 219499 200701
rect 123569 200696 219499 200698
rect 123569 200640 123574 200696
rect 123630 200640 219438 200696
rect 219494 200640 219499 200696
rect 123569 200638 219499 200640
rect 123569 200635 123635 200638
rect 219433 200635 219499 200638
rect 279926 200426 279986 200668
rect 286133 200426 286199 200429
rect 279926 200424 286199 200426
rect 279926 200368 286138 200424
rect 286194 200368 286199 200424
rect 279926 200366 286199 200368
rect 286133 200363 286199 200366
rect 238201 200290 238267 200293
rect 238201 200288 239690 200290
rect 238201 200232 238206 200288
rect 238262 200232 239690 200288
rect 238201 200230 239690 200232
rect 238201 200227 238267 200230
rect 239630 200222 239690 200230
rect 239630 200162 240212 200222
rect 75913 200018 75979 200021
rect 94497 200018 94563 200021
rect 75913 200016 94563 200018
rect 75913 199960 75918 200016
rect 75974 199960 94502 200016
rect 94558 199960 94563 200016
rect 75913 199958 94563 199960
rect 75913 199955 75979 199958
rect 94497 199955 94563 199958
rect 95969 200018 96035 200021
rect 107653 200018 107719 200021
rect 95969 200016 107719 200018
rect 95969 199960 95974 200016
rect 96030 199960 107658 200016
rect 107714 199960 107719 200016
rect 95969 199958 107719 199960
rect 95969 199955 96035 199958
rect 107653 199955 107719 199958
rect 100615 199882 100681 199885
rect 228265 199882 228331 199885
rect 100615 199880 228331 199882
rect 100615 199824 100620 199880
rect 100676 199824 228270 199880
rect 228326 199824 228331 199880
rect 100615 199822 228331 199824
rect 100615 199819 100681 199822
rect 228265 199819 228331 199822
rect 82721 199746 82787 199749
rect 100661 199746 100727 199749
rect 82721 199744 100727 199746
rect 82721 199688 82726 199744
rect 82782 199688 100666 199744
rect 100722 199688 100727 199744
rect 82721 199686 100727 199688
rect 82721 199683 82787 199686
rect 100661 199683 100727 199686
rect 102593 199746 102659 199749
rect 228173 199746 228239 199749
rect 102593 199744 228239 199746
rect 102593 199688 102598 199744
rect 102654 199688 228178 199744
rect 228234 199688 228239 199744
rect 102593 199686 228239 199688
rect 102593 199683 102659 199686
rect 228173 199683 228239 199686
rect 105905 199610 105971 199613
rect 225413 199610 225479 199613
rect 105905 199608 225479 199610
rect 105905 199552 105910 199608
rect 105966 199552 225418 199608
rect 225474 199552 225479 199608
rect 105905 199550 225479 199552
rect 105905 199547 105971 199550
rect 225413 199547 225479 199550
rect 92381 199474 92447 199477
rect 104893 199474 104959 199477
rect 92381 199472 104959 199474
rect 92381 199416 92386 199472
rect 92442 199416 104898 199472
rect 104954 199416 104959 199472
rect 92381 199414 104959 199416
rect 92381 199411 92447 199414
rect 104893 199411 104959 199414
rect 107561 199474 107627 199477
rect 225965 199474 226031 199477
rect 107561 199472 226031 199474
rect 107561 199416 107566 199472
rect 107622 199416 225970 199472
rect 226026 199416 226031 199472
rect 107561 199414 226031 199416
rect 107561 199411 107627 199414
rect 225965 199411 226031 199414
rect 84101 199338 84167 199341
rect 95233 199338 95299 199341
rect 84101 199336 95299 199338
rect 84101 199280 84106 199336
rect 84162 199280 95238 199336
rect 95294 199280 95299 199336
rect 84101 199278 95299 199280
rect 84101 199275 84167 199278
rect 95233 199275 95299 199278
rect 108941 199338 109007 199341
rect 226149 199338 226215 199341
rect 108941 199336 226215 199338
rect 108941 199280 108946 199336
rect 109002 199280 226154 199336
rect 226210 199280 226215 199336
rect 108941 199278 226215 199280
rect 279926 199338 279986 199852
rect 286225 199338 286291 199341
rect 279926 199336 286291 199338
rect 279926 199280 286230 199336
rect 286286 199280 286291 199336
rect 279926 199278 286291 199280
rect 108941 199275 109007 199278
rect 226149 199275 226215 199278
rect 286225 199275 286291 199278
rect 3366 199140 3372 199204
rect 3436 199202 3442 199204
rect 116526 199202 116532 199204
rect 3436 199142 116532 199202
rect 3436 199140 3442 199142
rect 116526 199140 116532 199142
rect 116596 199140 116602 199204
rect 219433 199202 219499 199205
rect 226333 199202 226399 199205
rect 219433 199200 226399 199202
rect 219433 199144 219438 199200
rect 219494 199144 226338 199200
rect 226394 199144 226399 199200
rect 219433 199142 226399 199144
rect 219433 199139 219499 199142
rect 226333 199139 226399 199142
rect 237373 199202 237439 199205
rect 237373 199200 239690 199202
rect 237373 199144 237378 199200
rect 237434 199144 239690 199200
rect 237373 199142 239690 199144
rect 237373 199139 237439 199142
rect 239630 199134 239690 199142
rect 239630 199074 240212 199134
rect 94313 199066 94379 199069
rect 230933 199066 230999 199069
rect 94313 199064 230999 199066
rect 94313 199008 94318 199064
rect 94374 199008 230938 199064
rect 230994 199008 230999 199064
rect 94313 199006 230999 199008
rect 94313 199003 94379 199006
rect 230933 199003 230999 199006
rect 81065 198930 81131 198933
rect 103421 198930 103487 198933
rect 81065 198928 103487 198930
rect 81065 198872 81070 198928
rect 81126 198872 103426 198928
rect 103482 198872 103487 198928
rect 81065 198870 103487 198872
rect 81065 198867 81131 198870
rect 103421 198867 103487 198870
rect 91001 198794 91067 198797
rect 106273 198794 106339 198797
rect 91001 198792 106339 198794
rect 91001 198736 91006 198792
rect 91062 198736 106278 198792
rect 106334 198736 106339 198792
rect 91001 198734 106339 198736
rect 279926 198794 279986 199036
rect 286409 198794 286475 198797
rect 279926 198792 286475 198794
rect 279926 198736 286414 198792
rect 286470 198736 286475 198792
rect 279926 198734 286475 198736
rect 91001 198731 91067 198734
rect 106273 198731 106339 198734
rect 286409 198731 286475 198734
rect 445385 198794 445451 198797
rect 449157 198794 449223 198797
rect 445385 198792 449223 198794
rect 445385 198736 445390 198792
rect 445446 198736 449162 198792
rect 449218 198736 449223 198792
rect 445385 198734 449223 198736
rect 445385 198731 445451 198734
rect 449157 198731 449223 198734
rect 77753 198658 77819 198661
rect 223205 198658 223271 198661
rect 77753 198656 223271 198658
rect 77753 198600 77758 198656
rect 77814 198600 223210 198656
rect 223266 198600 223271 198656
rect 77753 198598 223271 198600
rect 77753 198595 77819 198598
rect 223205 198595 223271 198598
rect 50981 198522 51047 198525
rect 70393 198522 70459 198525
rect 50981 198520 70459 198522
rect 50981 198464 50986 198520
rect 51042 198464 70398 198520
rect 70454 198464 70459 198520
rect 50981 198462 70459 198464
rect 50981 198459 51047 198462
rect 70393 198459 70459 198462
rect 87689 198522 87755 198525
rect 231209 198522 231275 198525
rect 87689 198520 231275 198522
rect 87689 198464 87694 198520
rect 87750 198464 231214 198520
rect 231270 198464 231275 198520
rect 87689 198462 231275 198464
rect 87689 198459 87755 198462
rect 231209 198459 231275 198462
rect 64505 198386 64571 198389
rect 85573 198386 85639 198389
rect 64505 198384 85639 198386
rect 64505 198328 64510 198384
rect 64566 198328 85578 198384
rect 85634 198328 85639 198384
rect 64505 198326 85639 198328
rect 64505 198323 64571 198326
rect 85573 198323 85639 198326
rect 89345 198386 89411 198389
rect 231393 198386 231459 198389
rect 89345 198384 231459 198386
rect 89345 198328 89350 198384
rect 89406 198328 231398 198384
rect 231454 198328 231459 198384
rect 89345 198326 231459 198328
rect 89345 198323 89411 198326
rect 231393 198323 231459 198326
rect 57881 198250 57947 198253
rect 79317 198250 79383 198253
rect 57881 198248 79383 198250
rect 57881 198192 57886 198248
rect 57942 198192 79322 198248
rect 79378 198192 79383 198248
rect 57881 198190 79383 198192
rect 57881 198187 57947 198190
rect 79317 198187 79383 198190
rect 86033 198250 86099 198253
rect 222929 198250 222995 198253
rect 86033 198248 222995 198250
rect 86033 198192 86038 198248
rect 86094 198192 222934 198248
rect 222990 198192 222995 198248
rect 86033 198190 222995 198192
rect 86033 198187 86099 198190
rect 222929 198187 222995 198190
rect 72785 198114 72851 198117
rect 97993 198114 98059 198117
rect 72785 198112 98059 198114
rect 72785 198056 72790 198112
rect 72846 198056 97998 198112
rect 98054 198056 98059 198112
rect 72785 198054 98059 198056
rect 72785 198051 72851 198054
rect 97993 198051 98059 198054
rect 226333 198114 226399 198117
rect 226333 198112 239690 198114
rect 226333 198056 226338 198112
rect 226394 198056 239690 198112
rect 226333 198054 239690 198056
rect 226333 198051 226399 198054
rect 239630 198046 239690 198054
rect 239630 197986 240212 198046
rect 69473 197978 69539 197981
rect 88333 197978 88399 197981
rect 69473 197976 88399 197978
rect 69473 197920 69478 197976
rect 69534 197920 88338 197976
rect 88394 197920 88399 197976
rect 69473 197918 88399 197920
rect 69473 197915 69539 197918
rect 88333 197915 88399 197918
rect 99189 197978 99255 197981
rect 228357 197978 228423 197981
rect 99189 197976 228423 197978
rect 99189 197920 99194 197976
rect 99250 197920 228362 197976
rect 228418 197920 228423 197976
rect 99189 197918 228423 197920
rect 99189 197915 99255 197918
rect 228357 197915 228423 197918
rect 56225 197842 56291 197845
rect 71773 197842 71839 197845
rect 56225 197840 71839 197842
rect 56225 197784 56230 197840
rect 56286 197784 71778 197840
rect 71834 197784 71839 197840
rect 56225 197782 71839 197784
rect 56225 197779 56291 197782
rect 71773 197779 71839 197782
rect 104249 197842 104315 197845
rect 225781 197842 225847 197845
rect 104249 197840 225847 197842
rect 104249 197784 104254 197840
rect 104310 197784 225786 197840
rect 225842 197784 225847 197840
rect 104249 197782 225847 197784
rect 104249 197779 104315 197782
rect 225781 197779 225847 197782
rect 54569 197706 54635 197709
rect 73153 197706 73219 197709
rect 54569 197704 73219 197706
rect 54569 197648 54574 197704
rect 54630 197648 73158 197704
rect 73214 197648 73219 197704
rect 54569 197646 73219 197648
rect 54569 197643 54635 197646
rect 73153 197643 73219 197646
rect 74441 197706 74507 197709
rect 96613 197706 96679 197709
rect 74441 197704 96679 197706
rect 74441 197648 74446 197704
rect 74502 197648 96618 197704
rect 96674 197648 96679 197704
rect 74441 197646 96679 197648
rect 279926 197706 279986 198220
rect 286501 197706 286567 197709
rect 279926 197704 286567 197706
rect 279926 197648 286506 197704
rect 286562 197648 286567 197704
rect 279926 197646 286567 197648
rect 74441 197643 74507 197646
rect 96613 197643 96679 197646
rect 286501 197643 286567 197646
rect 71129 197570 71195 197573
rect 86953 197570 87019 197573
rect 71129 197568 87019 197570
rect 71129 197512 71134 197568
rect 71190 197512 86958 197568
rect 87014 197512 87019 197568
rect 71129 197510 87019 197512
rect 71129 197507 71195 197510
rect 86953 197507 87019 197510
rect 97625 197570 97691 197573
rect 228541 197570 228607 197573
rect 97625 197568 228607 197570
rect 97625 197512 97630 197568
rect 97686 197512 228546 197568
rect 228602 197512 228607 197568
rect 97625 197510 228607 197512
rect 97625 197507 97691 197510
rect 228541 197507 228607 197510
rect 279926 197510 280170 197570
rect 52913 197434 52979 197437
rect 78581 197434 78647 197437
rect 52913 197432 78647 197434
rect 52913 197376 52918 197432
rect 52974 197376 78586 197432
rect 78642 197376 78647 197432
rect 52913 197374 78647 197376
rect 52913 197371 52979 197374
rect 78581 197371 78647 197374
rect 79409 197434 79475 197437
rect 104157 197434 104223 197437
rect 79409 197432 104223 197434
rect 79409 197376 79414 197432
rect 79470 197376 104162 197432
rect 104218 197376 104223 197432
rect 279926 197404 279986 197510
rect 280110 197434 280170 197510
rect 285765 197434 285831 197437
rect 280110 197432 285831 197434
rect 79409 197374 104223 197376
rect 280110 197376 285770 197432
rect 285826 197376 285831 197432
rect 280110 197374 285831 197376
rect 79409 197371 79475 197374
rect 104157 197371 104223 197374
rect 285765 197371 285831 197374
rect 67541 197298 67607 197301
rect 225597 197298 225663 197301
rect 67541 197296 225663 197298
rect 67541 197240 67546 197296
rect 67602 197240 225602 197296
rect 225658 197240 225663 197296
rect 67541 197238 225663 197240
rect 67541 197235 67607 197238
rect 225597 197235 225663 197238
rect 238385 197026 238451 197029
rect 238385 197024 239690 197026
rect 238385 196968 238390 197024
rect 238446 196968 239690 197024
rect 238385 196966 239690 196968
rect 238385 196963 238451 196966
rect 239630 196958 239690 196966
rect 239630 196898 240212 196958
rect 279926 196210 279986 196588
rect 279926 196150 282562 196210
rect 281349 196074 281415 196077
rect 282361 196074 282427 196077
rect 281349 196072 282427 196074
rect 281349 196016 281354 196072
rect 281410 196016 282366 196072
rect 282422 196016 282427 196072
rect 281349 196014 282427 196016
rect 282502 196074 282562 196150
rect 285673 196074 285739 196077
rect 282502 196072 285739 196074
rect 282502 196016 285678 196072
rect 285734 196016 285739 196072
rect 282502 196014 285739 196016
rect 281349 196011 281415 196014
rect 282361 196011 282427 196014
rect 285673 196011 285739 196014
rect 234521 195938 234587 195941
rect 234521 195936 239690 195938
rect 234521 195880 234526 195936
rect 234582 195880 239690 195936
rect 234521 195878 239690 195880
rect 234521 195875 234587 195878
rect 239630 195870 239690 195878
rect 239630 195810 240212 195870
rect 279926 195666 279986 195772
rect 285622 195740 285628 195804
rect 285692 195740 285698 195804
rect 285630 195666 285690 195740
rect 279926 195606 285690 195666
rect 95141 195258 95207 195261
rect 216029 195258 216095 195261
rect 95141 195256 216095 195258
rect 95141 195200 95146 195256
rect 95202 195200 216034 195256
rect 216090 195200 216095 195256
rect 95141 195198 216095 195200
rect 95141 195195 95207 195198
rect 216029 195195 216095 195198
rect 342846 195196 342852 195260
rect 342916 195258 342922 195260
rect 580206 195258 580212 195260
rect 342916 195198 580212 195258
rect 342916 195196 342922 195198
rect 580206 195196 580212 195198
rect 580276 195196 580282 195260
rect 233141 194850 233207 194853
rect 279926 194850 279986 194956
rect 280654 194924 280660 194988
rect 280724 194924 280730 194988
rect 280662 194850 280722 194924
rect 233141 194848 239690 194850
rect 233141 194792 233146 194848
rect 233202 194792 239690 194848
rect 233141 194790 239690 194792
rect 279926 194790 280722 194850
rect 442901 194850 442967 194853
rect 445385 194850 445451 194853
rect 442901 194848 445451 194850
rect 442901 194792 442906 194848
rect 442962 194792 445390 194848
rect 445446 194792 445451 194848
rect 442901 194790 445451 194792
rect 233141 194787 233207 194790
rect 239630 194782 239690 194790
rect 442901 194787 442967 194790
rect 445385 194787 445451 194790
rect 239630 194722 240212 194782
rect 15837 193898 15903 193901
rect 238109 193898 238175 193901
rect 15837 193896 238175 193898
rect 15837 193840 15842 193896
rect 15898 193840 238114 193896
rect 238170 193840 238175 193896
rect 15837 193838 238175 193840
rect 15837 193835 15903 193838
rect 238109 193835 238175 193838
rect 231761 193762 231827 193765
rect 231761 193760 239690 193762
rect 231761 193704 231766 193760
rect 231822 193704 239690 193760
rect 231761 193702 239690 193704
rect 231761 193699 231827 193702
rect 239630 193694 239690 193702
rect 239630 193634 240212 193694
rect 279926 193626 279986 194140
rect 284293 193626 284359 193629
rect 279926 193624 284359 193626
rect 279926 193568 284298 193624
rect 284354 193568 284359 193624
rect 279926 193566 284359 193568
rect 284293 193563 284359 193566
rect 279926 193430 280170 193490
rect 279926 193324 279986 193430
rect 280110 193354 280170 193430
rect 282269 193354 282335 193357
rect 280110 193352 282335 193354
rect 280110 193296 282274 193352
rect 282330 193296 282335 193352
rect 280110 193294 282335 193296
rect 282269 193291 282335 193294
rect 235533 192674 235599 192677
rect 235533 192672 239690 192674
rect 235533 192616 235538 192672
rect 235594 192616 239690 192672
rect 235533 192614 239690 192616
rect 235533 192611 235599 192614
rect 239630 192606 239690 192614
rect 239630 192546 240212 192606
rect 112805 192538 112871 192541
rect 228909 192538 228975 192541
rect 112805 192536 228975 192538
rect 112805 192480 112810 192536
rect 112866 192480 228914 192536
rect 228970 192480 228975 192536
rect 112805 192478 228975 192480
rect 112805 192475 112871 192478
rect 228909 192475 228975 192478
rect 279926 192402 279986 192508
rect 284518 192476 284524 192540
rect 284588 192476 284594 192540
rect 580441 192538 580507 192541
rect 583520 192538 584960 192628
rect 580441 192536 584960 192538
rect 580441 192480 580446 192536
rect 580502 192480 584960 192536
rect 580441 192478 584960 192480
rect 284526 192402 284586 192476
rect 580441 192475 580507 192478
rect 279926 192342 284586 192402
rect 583520 192388 584960 192478
rect 436001 191722 436067 191725
rect 439497 191722 439563 191725
rect 436001 191720 439563 191722
rect 237097 191586 237163 191589
rect 237097 191584 239690 191586
rect 237097 191528 237102 191584
rect 237158 191528 239690 191584
rect 237097 191526 239690 191528
rect 237097 191523 237163 191526
rect 239630 191518 239690 191526
rect 239630 191458 240212 191518
rect 279926 191178 279986 191692
rect 436001 191664 436006 191720
rect 436062 191664 439502 191720
rect 439558 191664 439563 191720
rect 436001 191662 439563 191664
rect 436001 191659 436067 191662
rect 439497 191659 439563 191662
rect 279926 191118 280170 191178
rect 280110 191042 280170 191118
rect 283005 191042 283071 191045
rect 280110 191040 283071 191042
rect 280110 190984 283010 191040
rect 283066 190984 283071 191040
rect 280110 190982 283071 190984
rect 283005 190979 283071 190982
rect 279926 190634 279986 190876
rect 282361 190634 282427 190637
rect 279926 190632 282427 190634
rect 279926 190576 282366 190632
rect 282422 190576 282427 190632
rect 279926 190574 282427 190576
rect 282361 190571 282427 190574
rect 442901 190498 442967 190501
rect 440190 190496 442967 190498
rect 440190 190440 442906 190496
rect 442962 190440 442967 190496
rect 440190 190438 442967 190440
rect 239630 190370 240212 190430
rect 237189 190362 237255 190365
rect 239630 190362 239690 190370
rect 237189 190360 239690 190362
rect 237189 190304 237194 190360
rect 237250 190304 239690 190360
rect 237189 190302 239690 190304
rect 436093 190362 436159 190365
rect 440190 190362 440250 190438
rect 442901 190435 442967 190438
rect 436093 190360 440250 190362
rect 436093 190304 436098 190360
rect 436154 190304 440250 190360
rect 436093 190302 440250 190304
rect 237189 190299 237255 190302
rect 436093 190299 436159 190302
rect 279926 190166 287070 190226
rect 279926 190060 279986 190166
rect 287010 190090 287070 190166
rect 289813 190090 289879 190093
rect 287010 190088 289879 190090
rect 287010 190032 289818 190088
rect 289874 190032 289879 190088
rect 287010 190030 289879 190032
rect 289813 190027 289879 190030
rect 235942 189348 235948 189412
rect 236012 189410 236018 189412
rect 236012 189350 239690 189410
rect 236012 189348 236018 189350
rect 239630 189342 239690 189350
rect 239630 189282 240212 189342
rect 279926 189138 279986 189244
rect 281574 189212 281580 189276
rect 281644 189212 281650 189276
rect 281582 189138 281642 189212
rect 279926 189078 281642 189138
rect -960 188866 480 188956
rect 231158 188866 231164 188868
rect -960 188806 231164 188866
rect -960 188716 480 188806
rect 231158 188804 231164 188806
rect 231228 188804 231234 188868
rect 279926 188534 287070 188594
rect 279926 188428 279986 188534
rect 287010 188458 287070 188534
rect 287789 188458 287855 188461
rect 287010 188456 287855 188458
rect 287010 188400 287794 188456
rect 287850 188400 287855 188456
rect 287010 188398 287855 188400
rect 287789 188395 287855 188398
rect 237230 188260 237236 188324
rect 237300 188322 237306 188324
rect 237300 188262 239690 188322
rect 237300 188260 237306 188262
rect 239630 188254 239690 188262
rect 239630 188194 240212 188254
rect 434621 187778 434687 187781
rect 436093 187778 436159 187781
rect 434621 187776 436159 187778
rect 434621 187720 434626 187776
rect 434682 187720 436098 187776
rect 436154 187720 436159 187776
rect 434621 187718 436159 187720
rect 434621 187715 434687 187718
rect 436093 187715 436159 187718
rect 287605 187642 287671 187645
rect 287010 187640 287671 187642
rect 279926 187506 279986 187612
rect 287010 187584 287610 187640
rect 287666 187584 287671 187640
rect 287010 187582 287671 187584
rect 287010 187506 287070 187582
rect 287605 187579 287671 187582
rect 279926 187446 287070 187506
rect 235809 187234 235875 187237
rect 235809 187232 239690 187234
rect 235809 187176 235814 187232
rect 235870 187176 239690 187232
rect 235809 187174 239690 187176
rect 235809 187171 235875 187174
rect 239630 187166 239690 187174
rect 239630 187106 240212 187166
rect 279926 186902 287070 186962
rect 279926 186796 279986 186902
rect 287010 186826 287070 186902
rect 287697 186826 287763 186829
rect 287010 186824 287763 186826
rect 287010 186768 287702 186824
rect 287758 186768 287763 186824
rect 287010 186766 287763 186768
rect 287697 186763 287763 186766
rect 237966 186084 237972 186148
rect 238036 186146 238042 186148
rect 238036 186086 239690 186146
rect 238036 186084 238042 186086
rect 239630 186078 239690 186086
rect 279926 186086 287070 186146
rect 239630 186018 240212 186078
rect 279926 185980 279986 186086
rect 287010 186010 287070 186086
rect 287881 186010 287947 186013
rect 287010 186008 287947 186010
rect 287010 185952 287886 186008
rect 287942 185952 287947 186008
rect 287010 185950 287947 185952
rect 287881 185947 287947 185950
rect 429193 185602 429259 185605
rect 436001 185602 436067 185605
rect 429193 185600 436067 185602
rect 429193 185544 429198 185600
rect 429254 185544 436006 185600
rect 436062 185544 436067 185600
rect 429193 185542 436067 185544
rect 429193 185539 429259 185542
rect 436001 185539 436067 185542
rect 279926 185058 279986 185164
rect 284702 185132 284708 185196
rect 284772 185132 284778 185196
rect 284710 185058 284770 185132
rect 279926 184998 284770 185058
rect 239814 184930 240212 184990
rect 235717 184922 235783 184925
rect 239814 184922 239874 184930
rect 235717 184920 239874 184922
rect 235717 184864 235722 184920
rect 235778 184864 239874 184920
rect 235717 184862 239874 184864
rect 428457 184922 428523 184925
rect 434621 184922 434687 184925
rect 428457 184920 434687 184922
rect 428457 184864 428462 184920
rect 428518 184864 434626 184920
rect 434682 184864 434687 184920
rect 428457 184862 434687 184864
rect 235717 184859 235783 184862
rect 428457 184859 428523 184862
rect 434621 184859 434687 184862
rect 279926 184242 279986 184348
rect 283414 184316 283420 184380
rect 283484 184316 283490 184380
rect 283422 184242 283482 184316
rect 279926 184182 283482 184242
rect 239630 183842 240212 183902
rect 238569 183834 238635 183837
rect 239630 183834 239690 183842
rect 238569 183832 239690 183834
rect 238569 183776 238574 183832
rect 238630 183776 239690 183832
rect 238569 183774 239690 183776
rect 238569 183771 238635 183774
rect 279366 183500 279372 183564
rect 279436 183500 279442 183564
rect 426433 183154 426499 183157
rect 429193 183154 429259 183157
rect 426433 183152 429259 183154
rect 426433 183096 426438 183152
rect 426494 183096 429198 183152
rect 429254 183096 429259 183152
rect 426433 183094 429259 183096
rect 426433 183091 426499 183094
rect 429193 183091 429259 183094
rect 239630 182754 240212 182814
rect 237782 182684 237788 182748
rect 237852 182746 237858 182748
rect 239630 182746 239690 182754
rect 237852 182686 239690 182746
rect 237852 182684 237858 182686
rect 279926 182610 279986 182716
rect 281022 182684 281028 182748
rect 281092 182684 281098 182748
rect 281030 182610 281090 182684
rect 279926 182550 281090 182610
rect 279926 181794 279986 181900
rect 282126 181868 282132 181932
rect 282196 181868 282202 181932
rect 282134 181794 282194 181868
rect 279926 181734 282194 181794
rect 239630 181666 240212 181726
rect 237966 181596 237972 181660
rect 238036 181658 238042 181660
rect 239630 181658 239690 181666
rect 238036 181598 239690 181658
rect 238036 181596 238042 181598
rect 31293 181386 31359 181389
rect 223297 181386 223363 181389
rect 31293 181384 223363 181386
rect 31293 181328 31298 181384
rect 31354 181328 223302 181384
rect 223358 181328 223363 181384
rect 31293 181326 223363 181328
rect 31293 181323 31359 181326
rect 223297 181323 223363 181326
rect 279926 181190 287070 181250
rect 279926 181084 279986 181190
rect 287010 181114 287070 181190
rect 289077 181114 289143 181117
rect 287010 181112 289143 181114
rect 287010 181056 289082 181112
rect 289138 181056 289143 181112
rect 287010 181054 289143 181056
rect 289077 181051 289143 181054
rect 239622 180576 239628 180640
rect 239692 180638 239698 180640
rect 239692 180578 240212 180638
rect 239692 180576 239698 180578
rect 279926 180162 279986 180268
rect 283046 180236 283052 180300
rect 283116 180236 283122 180300
rect 283054 180162 283114 180236
rect 279926 180102 283114 180162
rect 279926 179558 283298 179618
rect 239806 179488 239812 179552
rect 239876 179550 239882 179552
rect 239876 179490 240212 179550
rect 239876 179488 239882 179490
rect 279926 179452 279986 179558
rect 283238 179484 283298 179558
rect 283230 179420 283236 179484
rect 283300 179420 283306 179484
rect 427077 179482 427143 179485
rect 428457 179482 428523 179485
rect 427077 179480 428523 179482
rect 427077 179424 427082 179480
rect 427138 179424 428462 179480
rect 428518 179424 428523 179480
rect 427077 179422 428523 179424
rect 427077 179419 427143 179422
rect 428457 179419 428523 179422
rect 288934 179148 288940 179212
rect 289004 179210 289010 179212
rect 583520 179210 584960 179300
rect 289004 179150 584960 179210
rect 289004 179148 289010 179150
rect 583520 179060 584960 179150
rect 239765 178462 239831 178465
rect 239765 178460 240212 178462
rect 239765 178404 239770 178460
rect 239826 178404 240212 178460
rect 239765 178402 240212 178404
rect 239765 178399 239831 178402
rect 279926 178122 279986 178636
rect 282453 178122 282519 178125
rect 279926 178120 282519 178122
rect 279926 178064 282458 178120
rect 282514 178064 282519 178120
rect 279926 178062 282519 178064
rect 282453 178059 282519 178062
rect 288750 177850 288756 177852
rect 279926 177714 279986 177820
rect 287010 177790 288756 177850
rect 287010 177714 287070 177790
rect 288750 177788 288756 177790
rect 288820 177788 288826 177852
rect 279926 177654 287070 177714
rect 239857 177374 239923 177377
rect 239857 177372 240212 177374
rect 239857 177316 239862 177372
rect 239918 177316 240212 177372
rect 239857 177314 240212 177316
rect 239857 177311 239923 177314
rect 279926 176898 279986 177004
rect 282821 176898 282887 176901
rect 279926 176896 282887 176898
rect 279926 176840 282826 176896
rect 282882 176840 282887 176896
rect 279926 176838 282887 176840
rect 282821 176835 282887 176838
rect 290590 176218 290596 176220
rect 279926 176082 279986 176188
rect 287010 176158 290596 176218
rect 287010 176082 287070 176158
rect 290590 176156 290596 176158
rect 290660 176156 290666 176220
rect -960 175796 480 176036
rect 279926 176022 287070 176082
rect 425697 176082 425763 176085
rect 427077 176082 427143 176085
rect 425697 176080 427143 176082
rect 425697 176024 425702 176080
rect 425758 176024 427082 176080
rect 427138 176024 427143 176080
rect 425697 176022 427143 176024
rect 425697 176019 425763 176022
rect 427077 176019 427143 176022
rect 421557 175946 421623 175949
rect 426341 175946 426407 175949
rect 421557 175944 426407 175946
rect 421557 175888 421562 175944
rect 421618 175888 426346 175944
rect 426402 175888 426407 175944
rect 421557 175886 426407 175888
rect 421557 175883 421623 175886
rect 426341 175883 426407 175886
rect 279926 175478 287070 175538
rect 279926 175372 279986 175478
rect 287010 175402 287070 175478
rect 294454 175402 294460 175404
rect 287010 175342 294460 175402
rect 294454 175340 294460 175342
rect 294524 175340 294530 175404
rect 279926 174662 284402 174722
rect 279926 174556 279986 174662
rect 284342 174588 284402 174662
rect 284334 174524 284340 174588
rect 284404 174524 284410 174588
rect 279926 173846 282930 173906
rect 279926 173740 279986 173846
rect 282870 173772 282930 173846
rect 282862 173708 282868 173772
rect 282932 173708 282938 173772
rect 282913 173634 282979 173637
rect 279926 173632 282979 173634
rect 279926 173576 282918 173632
rect 282974 173576 282979 173632
rect 279926 173574 282979 173576
rect 279926 172924 279986 173574
rect 282913 173571 282979 173574
rect 282821 172274 282887 172277
rect 279926 172272 282887 172274
rect 279926 172216 282826 172272
rect 282882 172216 282887 172272
rect 279926 172214 282887 172216
rect 279926 172108 279986 172214
rect 282821 172211 282887 172214
rect 282729 171866 282795 171869
rect 279926 171864 282795 171866
rect 279926 171808 282734 171864
rect 282790 171808 282795 171864
rect 279926 171806 282795 171808
rect 279926 171292 279986 171806
rect 282729 171803 282795 171806
rect 282821 170778 282887 170781
rect 279926 170776 282887 170778
rect 279926 170720 282826 170776
rect 282882 170720 282887 170776
rect 279926 170718 282887 170720
rect 279926 170476 279986 170718
rect 282821 170715 282887 170718
rect 282821 169690 282887 169693
rect 280110 169688 282887 169690
rect 279926 169554 279986 169660
rect 280110 169632 282826 169688
rect 282882 169632 282887 169688
rect 280110 169630 282887 169632
rect 280110 169554 280170 169630
rect 282821 169627 282887 169630
rect 279926 169494 280170 169554
rect 282821 169282 282887 169285
rect 279926 169280 282887 169282
rect 279926 169224 282826 169280
rect 282882 169224 282887 169280
rect 279926 169222 282887 169224
rect 279926 168844 279986 169222
rect 282821 169219 282887 169222
rect 282821 168194 282887 168197
rect 279926 168192 282887 168194
rect 279926 168136 282826 168192
rect 282882 168136 282887 168192
rect 279926 168134 282887 168136
rect 279926 168028 279986 168134
rect 282821 168131 282887 168134
rect 282729 167786 282795 167789
rect 279926 167784 282795 167786
rect 279926 167728 282734 167784
rect 282790 167728 282795 167784
rect 279926 167726 282795 167728
rect 279926 167212 279986 167726
rect 282729 167723 282795 167726
rect 421557 166426 421623 166429
rect 287010 166424 421623 166426
rect 279926 166290 279986 166396
rect 287010 166368 421562 166424
rect 421618 166368 421623 166424
rect 287010 166366 421623 166368
rect 287010 166290 287070 166366
rect 421557 166363 421623 166366
rect 279926 166230 287070 166290
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 425697 165610 425763 165613
rect 287010 165608 425763 165610
rect 279926 165474 279986 165580
rect 287010 165552 425702 165608
rect 425758 165552 425763 165608
rect 287010 165550 425763 165552
rect 287010 165474 287070 165550
rect 425697 165547 425763 165550
rect 279926 165414 287070 165474
rect 482369 164794 482435 164797
rect 287010 164792 482435 164794
rect 279926 164658 279986 164764
rect 287010 164736 482374 164792
rect 482430 164736 482435 164792
rect 287010 164734 482435 164736
rect 287010 164658 287070 164734
rect 482369 164731 482435 164734
rect 279926 164598 287070 164658
rect 499573 163978 499639 163981
rect 287010 163976 499639 163978
rect 279926 163842 279986 163948
rect 287010 163920 499578 163976
rect 499634 163920 499639 163976
rect 287010 163918 499639 163920
rect 287010 163842 287070 163918
rect 499573 163915 499639 163918
rect 279926 163782 287070 163842
rect 540237 163162 540303 163165
rect 287010 163160 540303 163162
rect 279926 163026 279986 163132
rect 287010 163104 540242 163160
rect 540298 163104 540303 163160
rect 287010 163102 540303 163104
rect 287010 163026 287070 163102
rect 540237 163099 540303 163102
rect -960 162890 480 162980
rect 279926 162966 287070 163026
rect 40677 162890 40743 162893
rect -960 162888 40743 162890
rect -960 162832 40682 162888
rect 40738 162832 40743 162888
rect -960 162830 40743 162832
rect -960 162740 480 162830
rect 40677 162827 40743 162830
rect 555366 162346 555372 162348
rect 279926 162210 279986 162316
rect 287010 162286 555372 162346
rect 287010 162210 287070 162286
rect 555366 162284 555372 162286
rect 555436 162284 555442 162348
rect 279926 162150 287070 162210
rect 279742 161606 287070 161666
rect 279742 161500 279802 161606
rect 287010 161530 287070 161606
rect 551134 161530 551140 161532
rect 287010 161470 551140 161530
rect 551134 161468 551140 161470
rect 551204 161468 551210 161532
rect 548374 160714 548380 160716
rect 279926 160578 279986 160684
rect 287010 160654 548380 160714
rect 287010 160578 287070 160654
rect 548374 160652 548380 160654
rect 548444 160652 548450 160716
rect 279926 160518 287070 160578
rect 547086 159898 547092 159900
rect 279926 159762 279986 159868
rect 287010 159838 547092 159898
rect 287010 159762 287070 159838
rect 547086 159836 547092 159838
rect 547156 159836 547162 159900
rect 279926 159702 287070 159762
rect 544326 159082 544332 159084
rect 279926 158946 279986 159052
rect 287010 159022 544332 159082
rect 287010 158946 287070 159022
rect 544326 159020 544332 159022
rect 544396 159020 544402 159084
rect 279926 158886 287070 158946
rect 558126 158266 558132 158268
rect 279926 158130 279986 158236
rect 287010 158206 558132 158266
rect 287010 158130 287070 158206
rect 558126 158204 558132 158206
rect 558196 158204 558202 158268
rect 279926 158070 287070 158130
rect 279926 157526 287070 157586
rect 279926 157420 279986 157526
rect 287010 157450 287070 157526
rect 295926 157450 295932 157452
rect 287010 157390 295932 157450
rect 295926 157388 295932 157390
rect 295996 157388 296002 157452
rect 345606 156634 345612 156636
rect 279926 156498 279986 156604
rect 287010 156574 345612 156634
rect 287010 156498 287070 156574
rect 345606 156572 345612 156574
rect 345676 156572 345682 156636
rect 279926 156438 287070 156498
rect 287646 155818 287652 155820
rect 279926 155682 279986 155788
rect 287010 155758 287652 155818
rect 287010 155682 287070 155758
rect 287646 155756 287652 155758
rect 287716 155756 287722 155820
rect 279926 155622 287070 155682
rect 342846 155002 342852 155004
rect 279926 154866 279986 154972
rect 287010 154942 342852 155002
rect 287010 154866 287070 154942
rect 342846 154940 342852 154942
rect 342916 154940 342922 155004
rect 279926 154806 287070 154866
rect 288934 154186 288940 154188
rect 279926 154050 279986 154156
rect 287010 154126 288940 154186
rect 287010 154050 287070 154126
rect 288934 154124 288940 154126
rect 289004 154124 289010 154188
rect 279926 153990 287070 154050
rect 351126 153370 351132 153372
rect 279926 153234 279986 153340
rect 287010 153310 351132 153370
rect 287010 153234 287070 153310
rect 351126 153308 351132 153310
rect 351196 153308 351202 153372
rect 279926 153174 287070 153234
rect 580533 152690 580599 152693
rect 583520 152690 584960 152780
rect 580533 152688 584960 152690
rect 580533 152632 580538 152688
rect 580594 152632 584960 152688
rect 580533 152630 584960 152632
rect 580533 152627 580599 152630
rect 306966 152554 306972 152556
rect 279926 152418 279986 152524
rect 287010 152494 306972 152554
rect 287010 152418 287070 152494
rect 306966 152492 306972 152494
rect 307036 152492 307042 152556
rect 583520 152540 584960 152630
rect 279926 152358 287070 152418
rect 288934 151738 288940 151740
rect 279926 151602 279986 151708
rect 287010 151678 288940 151738
rect 287010 151602 287070 151678
rect 288934 151676 288940 151678
rect 289004 151676 289010 151740
rect 279926 151542 287070 151602
rect 551134 150922 551140 150924
rect 279926 150786 279986 150892
rect 287010 150862 551140 150922
rect 287010 150786 287070 150862
rect 551134 150860 551140 150862
rect 551204 150860 551210 150924
rect 279926 150726 287070 150786
rect -960 149834 480 149924
rect 3366 149834 3372 149836
rect -960 149774 3372 149834
rect -960 149684 480 149774
rect 3366 149772 3372 149774
rect 3436 149772 3442 149836
rect 237281 146978 237347 146981
rect 237281 146976 239690 146978
rect 237281 146920 237286 146976
rect 237342 146920 239690 146976
rect 237281 146918 239690 146920
rect 237281 146915 237347 146918
rect 239630 146910 239690 146918
rect 239630 146850 240212 146910
rect 239630 145762 240212 145822
rect 238201 145754 238267 145757
rect 239630 145754 239690 145762
rect 238201 145752 239690 145754
rect 238201 145696 238206 145752
rect 238262 145696 239690 145752
rect 238201 145694 239690 145696
rect 238201 145691 238267 145694
rect 240358 144672 240364 144736
rect 240428 144672 240434 144736
rect 23013 144122 23079 144125
rect 206277 144122 206343 144125
rect 23013 144120 206343 144122
rect 23013 144064 23018 144120
rect 23074 144064 206282 144120
rect 206338 144064 206343 144120
rect 23013 144062 206343 144064
rect 23013 144059 23079 144062
rect 206277 144059 206343 144062
rect 235901 143714 235967 143717
rect 235901 143712 239690 143714
rect 235901 143656 235906 143712
rect 235962 143656 239690 143712
rect 235901 143654 239690 143656
rect 235901 143651 235967 143654
rect 239630 143646 239690 143654
rect 239630 143586 240212 143646
rect 240174 142496 240180 142560
rect 240244 142496 240250 142560
rect 232078 142020 232084 142084
rect 232148 142082 232154 142084
rect 292614 142082 292620 142084
rect 232148 142022 292620 142082
rect 232148 142020 232154 142022
rect 292614 142020 292620 142022
rect 292684 142020 292690 142084
rect 232589 141946 232655 141949
rect 292665 141946 292731 141949
rect 232589 141944 292731 141946
rect 232589 141888 232594 141944
rect 232650 141888 292670 141944
rect 292726 141888 292731 141944
rect 232589 141886 292731 141888
rect 232589 141883 232655 141886
rect 292665 141883 292731 141886
rect 238385 141810 238451 141813
rect 289997 141810 290063 141813
rect 238385 141808 290063 141810
rect 238385 141752 238390 141808
rect 238446 141752 290002 141808
rect 290058 141752 290063 141808
rect 238385 141750 290063 141752
rect 238385 141747 238451 141750
rect 289997 141747 290063 141750
rect 238569 141674 238635 141677
rect 289905 141674 289971 141677
rect 238569 141672 289971 141674
rect 238569 141616 238574 141672
rect 238630 141616 289910 141672
rect 289966 141616 289971 141672
rect 238569 141614 289971 141616
rect 238569 141611 238635 141614
rect 289905 141611 289971 141614
rect 238334 141476 238340 141540
rect 238404 141538 238410 141540
rect 285806 141538 285812 141540
rect 238404 141478 285812 141538
rect 238404 141476 238410 141478
rect 285806 141476 285812 141478
rect 285876 141476 285882 141540
rect 105721 141402 105787 141405
rect 202137 141402 202203 141405
rect 105721 141400 202203 141402
rect 105721 141344 105726 141400
rect 105782 141344 202142 141400
rect 202198 141344 202203 141400
rect 105721 141342 202203 141344
rect 105721 141339 105787 141342
rect 202137 141339 202203 141342
rect 239581 141402 239647 141405
rect 240174 141402 240180 141404
rect 239581 141400 240180 141402
rect 239581 141344 239586 141400
rect 239642 141344 240180 141400
rect 239581 141342 240180 141344
rect 239581 141339 239647 141342
rect 240174 141340 240180 141342
rect 240244 141340 240250 141404
rect 273294 141340 273300 141404
rect 273364 141402 273370 141404
rect 290273 141402 290339 141405
rect 273364 141400 290339 141402
rect 273364 141344 290278 141400
rect 290334 141344 290339 141400
rect 273364 141342 290339 141344
rect 273364 141340 273370 141342
rect 290273 141339 290339 141342
rect 48630 140660 48636 140724
rect 48700 140722 48706 140724
rect 235901 140722 235967 140725
rect 48700 140720 235967 140722
rect 48700 140664 235906 140720
rect 235962 140664 235967 140720
rect 48700 140662 235967 140664
rect 48700 140660 48706 140662
rect 235901 140659 235967 140662
rect 237741 140724 237807 140725
rect 237741 140720 237788 140724
rect 237852 140722 237858 140724
rect 237741 140664 237746 140720
rect 237741 140660 237788 140664
rect 237852 140662 237898 140722
rect 237852 140660 237858 140662
rect 237966 140660 237972 140724
rect 238036 140722 238042 140724
rect 238477 140722 238543 140725
rect 239673 140724 239739 140725
rect 239622 140722 239628 140724
rect 238036 140720 238543 140722
rect 238036 140664 238482 140720
rect 238538 140664 238543 140720
rect 238036 140662 238543 140664
rect 239582 140662 239628 140722
rect 239692 140720 239739 140724
rect 239734 140664 239739 140720
rect 238036 140660 238042 140662
rect 237741 140659 237807 140660
rect 238477 140659 238543 140662
rect 239622 140660 239628 140662
rect 239692 140660 239739 140664
rect 239673 140659 239739 140660
rect 3366 140524 3372 140588
rect 3436 140586 3442 140588
rect 266905 140586 266971 140589
rect 3436 140584 266971 140586
rect 3436 140528 266910 140584
rect 266966 140528 266971 140584
rect 3436 140526 266971 140528
rect 3436 140524 3442 140526
rect 266905 140523 266971 140526
rect 275277 140586 275343 140589
rect 281533 140586 281599 140589
rect 275277 140584 281599 140586
rect 275277 140528 275282 140584
rect 275338 140528 281538 140584
rect 281594 140528 281599 140584
rect 275277 140526 281599 140528
rect 275277 140523 275343 140526
rect 281533 140523 281599 140526
rect 48446 140388 48452 140452
rect 48516 140450 48522 140452
rect 288750 140450 288756 140452
rect 48516 140390 288756 140450
rect 48516 140388 48522 140390
rect 288750 140388 288756 140390
rect 288820 140388 288826 140452
rect 59261 140314 59327 140317
rect 288801 140314 288867 140317
rect 59261 140312 288867 140314
rect 59261 140256 59266 140312
rect 59322 140256 288806 140312
rect 288862 140256 288867 140312
rect 59261 140254 288867 140256
rect 59261 140251 59327 140254
rect 288801 140251 288867 140254
rect 232957 140178 233023 140181
rect 291653 140178 291719 140181
rect 232957 140176 291719 140178
rect 232957 140120 232962 140176
rect 233018 140120 291658 140176
rect 291714 140120 291719 140176
rect 232957 140118 291719 140120
rect 232957 140115 233023 140118
rect 291653 140115 291719 140118
rect 201493 140042 201559 140045
rect 280521 140042 280587 140045
rect 201493 140040 280587 140042
rect 201493 139984 201498 140040
rect 201554 139984 280526 140040
rect 280582 139984 280587 140040
rect 201493 139982 280587 139984
rect 201493 139979 201559 139982
rect 280521 139979 280587 139982
rect 235257 139906 235323 139909
rect 290365 139906 290431 139909
rect 235257 139904 290431 139906
rect 235257 139848 235262 139904
rect 235318 139848 290370 139904
rect 290426 139848 290431 139904
rect 235257 139846 290431 139848
rect 235257 139843 235323 139846
rect 290365 139843 290431 139846
rect 232773 139770 232839 139773
rect 273294 139770 273300 139772
rect 232773 139768 273300 139770
rect 232773 139712 232778 139768
rect 232834 139712 273300 139768
rect 232773 139710 273300 139712
rect 232773 139707 232839 139710
rect 273294 139708 273300 139710
rect 273364 139708 273370 139772
rect 240777 139634 240843 139637
rect 240910 139634 240916 139636
rect 240777 139632 240916 139634
rect 240777 139576 240782 139632
rect 240838 139576 240916 139632
rect 240777 139574 240916 139576
rect 240777 139571 240843 139574
rect 240910 139572 240916 139574
rect 240980 139572 240986 139636
rect 266997 139634 267063 139637
rect 281809 139634 281875 139637
rect 266997 139632 281875 139634
rect 266997 139576 267002 139632
rect 267058 139576 281814 139632
rect 281870 139576 281875 139632
rect 266997 139574 281875 139576
rect 266997 139571 267063 139574
rect 281809 139571 281875 139574
rect 288750 139436 288756 139500
rect 288820 139498 288826 139500
rect 289077 139498 289143 139501
rect 288820 139496 289143 139498
rect 288820 139440 289082 139496
rect 289138 139440 289143 139496
rect 288820 139438 289143 139440
rect 288820 139436 288826 139438
rect 289077 139435 289143 139438
rect 206277 139362 206343 139365
rect 235717 139362 235783 139365
rect 206277 139360 235783 139362
rect 206277 139304 206282 139360
rect 206338 139304 235722 139360
rect 235778 139304 235783 139360
rect 206277 139302 235783 139304
rect 206277 139299 206343 139302
rect 235717 139299 235783 139302
rect 351126 139300 351132 139364
rect 351196 139362 351202 139364
rect 583520 139362 584960 139452
rect 351196 139302 584960 139362
rect 351196 139300 351202 139302
rect 235022 139164 235028 139228
rect 235092 139226 235098 139228
rect 236821 139226 236887 139229
rect 290181 139226 290247 139229
rect 235092 139166 236378 139226
rect 235092 139164 235098 139166
rect 187325 139090 187391 139093
rect 233141 139090 233207 139093
rect 187325 139088 233207 139090
rect 187325 139032 187330 139088
rect 187386 139032 233146 139088
rect 233202 139032 233207 139088
rect 187325 139030 233207 139032
rect 187325 139027 187391 139030
rect 233141 139027 233207 139030
rect 235758 139028 235764 139092
rect 235828 139090 235834 139092
rect 236318 139090 236378 139166
rect 236821 139224 290247 139226
rect 236821 139168 236826 139224
rect 236882 139168 290186 139224
rect 290242 139168 290247 139224
rect 583520 139212 584960 139302
rect 236821 139166 290247 139168
rect 236821 139163 236887 139166
rect 290181 139163 290247 139166
rect 291510 139090 291516 139092
rect 235828 139030 236194 139090
rect 236318 139030 291516 139090
rect 235828 139028 235834 139030
rect 62573 138954 62639 138957
rect 235901 138954 235967 138957
rect 62573 138952 235967 138954
rect 62573 138896 62578 138952
rect 62634 138896 235906 138952
rect 235962 138896 235967 138952
rect 62573 138894 235967 138896
rect 236134 138954 236194 139030
rect 291510 139028 291516 139030
rect 291580 139028 291586 139092
rect 291326 138954 291332 138956
rect 236134 138894 291332 138954
rect 62573 138891 62639 138894
rect 235901 138891 235967 138894
rect 291326 138892 291332 138894
rect 291396 138892 291402 138956
rect 60917 138818 60983 138821
rect 235625 138818 235691 138821
rect 60917 138816 235691 138818
rect 60917 138760 60922 138816
rect 60978 138760 235630 138816
rect 235686 138760 235691 138816
rect 60917 138758 235691 138760
rect 60917 138755 60983 138758
rect 235625 138755 235691 138758
rect 235942 138756 235948 138820
rect 236012 138818 236018 138820
rect 291142 138818 291148 138820
rect 236012 138758 291148 138818
rect 236012 138756 236018 138758
rect 291142 138756 291148 138758
rect 291212 138756 291218 138820
rect 183737 138682 183803 138685
rect 218053 138682 218119 138685
rect 183737 138680 218119 138682
rect 183737 138624 183742 138680
rect 183798 138624 218058 138680
rect 218114 138624 218119 138680
rect 183737 138622 218119 138624
rect 183737 138619 183803 138622
rect 218053 138619 218119 138622
rect 219249 138682 219315 138685
rect 235901 138682 235967 138685
rect 219249 138680 235967 138682
rect 219249 138624 219254 138680
rect 219310 138624 235906 138680
rect 235962 138624 235967 138680
rect 219249 138622 235967 138624
rect 219249 138619 219315 138622
rect 235901 138619 235967 138622
rect 215661 138546 215727 138549
rect 235809 138546 235875 138549
rect 215661 138544 235875 138546
rect 215661 138488 215666 138544
rect 215722 138488 235814 138544
rect 235870 138488 235875 138544
rect 215661 138486 235875 138488
rect 215661 138483 215727 138486
rect 235809 138483 235875 138486
rect 239254 138484 239260 138548
rect 239324 138546 239330 138548
rect 288566 138546 288572 138548
rect 239324 138486 288572 138546
rect 239324 138484 239330 138486
rect 288566 138484 288572 138486
rect 288636 138484 288642 138548
rect 176653 138410 176719 138413
rect 215293 138410 215359 138413
rect 290089 138410 290155 138413
rect 176653 138408 215359 138410
rect 176653 138352 176658 138408
rect 176714 138352 215298 138408
rect 215354 138352 215359 138408
rect 176653 138350 215359 138352
rect 176653 138347 176719 138350
rect 215293 138347 215359 138350
rect 234570 138408 290155 138410
rect 234570 138352 290094 138408
rect 290150 138352 290155 138408
rect 234570 138350 290155 138352
rect 144729 138274 144795 138277
rect 205633 138274 205699 138277
rect 144729 138272 205699 138274
rect 144729 138216 144734 138272
rect 144790 138216 205638 138272
rect 205694 138216 205699 138272
rect 144729 138214 205699 138216
rect 144729 138211 144795 138214
rect 205633 138211 205699 138214
rect 232497 138274 232563 138277
rect 232497 138272 234170 138274
rect 232497 138216 232502 138272
rect 232558 138216 234170 138272
rect 232497 138214 234170 138216
rect 232497 138211 232563 138214
rect 3366 138076 3372 138140
rect 3436 138138 3442 138140
rect 233877 138138 233943 138141
rect 3436 138136 233943 138138
rect 3436 138080 233882 138136
rect 233938 138080 233943 138136
rect 3436 138078 233943 138080
rect 234110 138138 234170 138214
rect 234570 138138 234630 138350
rect 290089 138347 290155 138350
rect 235073 138274 235139 138277
rect 238753 138274 238819 138277
rect 288382 138274 288388 138276
rect 235073 138272 238819 138274
rect 235073 138216 235078 138272
rect 235134 138216 238758 138272
rect 238814 138216 238819 138272
rect 235073 138214 238819 138216
rect 235073 138211 235139 138214
rect 238753 138211 238819 138214
rect 244230 138214 288388 138274
rect 234110 138078 234630 138138
rect 3436 138076 3442 138078
rect 233877 138075 233943 138078
rect 235390 138076 235396 138140
rect 235460 138138 235466 138140
rect 244230 138138 244290 138214
rect 288382 138212 288388 138214
rect 288452 138212 288458 138276
rect 235460 138078 244290 138138
rect 235460 138076 235466 138078
rect 65885 138002 65951 138005
rect 262121 138002 262187 138005
rect 65885 138000 262187 138002
rect 65885 137944 65890 138000
rect 65946 137944 262126 138000
rect 262182 137944 262187 138000
rect 65885 137942 262187 137944
rect 65885 137939 65951 137942
rect 262121 137939 262187 137942
rect 262305 138002 262371 138005
rect 285857 138002 285923 138005
rect 262305 138000 285923 138002
rect 262305 137944 262310 138000
rect 262366 137944 285862 138000
rect 285918 137944 285923 138000
rect 262305 137942 285923 137944
rect 262305 137939 262371 137942
rect 285857 137939 285923 137942
rect 26509 137866 26575 137869
rect 115841 137866 115907 137869
rect 26509 137864 115907 137866
rect 26509 137808 26514 137864
rect 26570 137808 115846 137864
rect 115902 137808 115907 137864
rect 26509 137806 115907 137808
rect 26509 137803 26575 137806
rect 115841 137803 115907 137806
rect 232262 137804 232268 137868
rect 232332 137866 232338 137868
rect 287094 137866 287100 137868
rect 232332 137806 287100 137866
rect 232332 137804 232338 137806
rect 287094 137804 287100 137806
rect 287164 137804 287170 137868
rect 17033 137730 17099 137733
rect 44173 137730 44239 137733
rect 17033 137728 44239 137730
rect 17033 137672 17038 137728
rect 17094 137672 44178 137728
rect 44234 137672 44239 137728
rect 17033 137670 44239 137672
rect 17033 137667 17099 137670
rect 44173 137667 44239 137670
rect 238150 137668 238156 137732
rect 238220 137730 238226 137732
rect 290774 137730 290780 137732
rect 238220 137670 290780 137730
rect 238220 137668 238226 137670
rect 290774 137668 290780 137670
rect 290844 137668 290850 137732
rect 21817 137594 21883 137597
rect 66161 137594 66227 137597
rect 21817 137592 66227 137594
rect 21817 137536 21822 137592
rect 21878 137536 66166 137592
rect 66222 137536 66227 137592
rect 21817 137534 66227 137536
rect 21817 137531 21883 137534
rect 66161 137531 66227 137534
rect 118785 137594 118851 137597
rect 277301 137594 277367 137597
rect 118785 137592 277367 137594
rect 118785 137536 118790 137592
rect 118846 137536 277306 137592
rect 277362 137536 277367 137592
rect 118785 137534 277367 137536
rect 118785 137531 118851 137534
rect 277301 137531 277367 137534
rect 115197 137458 115263 137461
rect 276105 137458 276171 137461
rect 115197 137456 276171 137458
rect 115197 137400 115202 137456
rect 115258 137400 276110 137456
rect 276166 137400 276171 137456
rect 115197 137398 276171 137400
rect 115197 137395 115263 137398
rect 276105 137395 276171 137398
rect 44265 137322 44331 137325
rect 252185 137322 252251 137325
rect 44265 137320 252251 137322
rect 44265 137264 44270 137320
rect 44326 137264 252190 137320
rect 252246 137264 252251 137320
rect 44265 137262 252251 137264
rect 44265 137259 44331 137262
rect 252185 137259 252251 137262
rect 254669 137322 254735 137325
rect 280153 137322 280219 137325
rect 254669 137320 280219 137322
rect 254669 137264 254674 137320
rect 254730 137264 280158 137320
rect 280214 137264 280219 137320
rect 254669 137262 280219 137264
rect 254669 137259 254735 137262
rect 280153 137259 280219 137262
rect 30097 137186 30163 137189
rect 118693 137186 118759 137189
rect 30097 137184 118759 137186
rect 30097 137128 30102 137184
rect 30158 137128 118698 137184
rect 118754 137128 118759 137184
rect 30097 137126 118759 137128
rect 30097 137123 30163 137126
rect 118693 137123 118759 137126
rect 247585 137186 247651 137189
rect 281717 137186 281783 137189
rect 247585 137184 281783 137186
rect 247585 137128 247590 137184
rect 247646 137128 281722 137184
rect 281778 137128 281783 137184
rect 247585 137126 281783 137128
rect 247585 137123 247651 137126
rect 281717 137123 281783 137126
rect 33593 137050 33659 137053
rect 233141 137050 233207 137053
rect 33593 137048 233207 137050
rect 33593 136992 33598 137048
rect 33654 136992 233146 137048
rect 233202 136992 233207 137048
rect 33593 136990 233207 136992
rect 33593 136987 33659 136990
rect 233141 136987 233207 136990
rect 37181 136914 37247 136917
rect 237373 136914 237439 136917
rect 37181 136912 237439 136914
rect -960 136778 480 136868
rect 37181 136856 37186 136912
rect 37242 136856 237378 136912
rect 237434 136856 237439 136912
rect 37181 136854 237439 136856
rect 37181 136851 37247 136854
rect 237373 136851 237439 136854
rect 3366 136778 3372 136780
rect -960 136718 3372 136778
rect -960 136628 480 136718
rect 3366 136716 3372 136718
rect 3436 136716 3442 136780
rect 40677 136778 40743 136781
rect 247033 136778 247099 136781
rect 40677 136776 247099 136778
rect 40677 136720 40682 136776
rect 40738 136720 247038 136776
rect 247094 136720 247099 136776
rect 40677 136718 247099 136720
rect 40677 136715 40743 136718
rect 247033 136715 247099 136718
rect 244089 136370 244155 136373
rect 280245 136370 280311 136373
rect 244089 136368 280311 136370
rect 244089 136312 244094 136368
rect 244150 136312 280250 136368
rect 280306 136312 280311 136368
rect 244089 136310 280311 136312
rect 244089 136307 244155 136310
rect 280245 136307 280311 136310
rect 166073 136234 166139 136237
rect 283465 136234 283531 136237
rect 166073 136232 283531 136234
rect 166073 136176 166078 136232
rect 166134 136176 283470 136232
rect 283526 136176 283531 136232
rect 166073 136174 283531 136176
rect 166073 136171 166139 136174
rect 283465 136171 283531 136174
rect 162485 136098 162551 136101
rect 283557 136098 283623 136101
rect 162485 136096 283623 136098
rect 162485 136040 162490 136096
rect 162546 136040 283562 136096
rect 283618 136040 283623 136096
rect 162485 136038 283623 136040
rect 162485 136035 162551 136038
rect 283557 136035 283623 136038
rect 239673 135962 239739 135965
rect 580257 135962 580323 135965
rect 239673 135960 580323 135962
rect 239673 135904 239678 135960
rect 239734 135904 580262 135960
rect 580318 135904 580323 135960
rect 239673 135902 580323 135904
rect 239673 135899 239739 135902
rect 580257 135899 580323 135902
rect 246297 134874 246363 134877
rect 281625 134874 281691 134877
rect 246297 134872 281691 134874
rect 246297 134816 246302 134872
rect 246358 134816 281630 134872
rect 281686 134816 281691 134872
rect 246297 134814 281691 134816
rect 246297 134811 246363 134814
rect 281625 134811 281691 134814
rect 194409 134738 194475 134741
rect 280429 134738 280495 134741
rect 194409 134736 280495 134738
rect 194409 134680 194414 134736
rect 194470 134680 280434 134736
rect 280490 134680 280495 134736
rect 194409 134678 280495 134680
rect 194409 134675 194475 134678
rect 280429 134675 280495 134678
rect 126973 134602 127039 134605
rect 283649 134602 283715 134605
rect 126973 134600 283715 134602
rect 126973 134544 126978 134600
rect 127034 134544 283654 134600
rect 283710 134544 283715 134600
rect 126973 134542 283715 134544
rect 126973 134539 127039 134542
rect 283649 134539 283715 134542
rect 28901 134466 28967 134469
rect 284702 134466 284708 134468
rect 28901 134464 284708 134466
rect 28901 134408 28906 134464
rect 28962 134408 284708 134464
rect 28901 134406 284708 134408
rect 28901 134403 28967 134406
rect 284702 134404 284708 134406
rect 284772 134404 284778 134468
rect 233417 133378 233483 133381
rect 285949 133378 286015 133381
rect 233417 133376 286015 133378
rect 233417 133320 233422 133376
rect 233478 133320 285954 133376
rect 286010 133320 286015 133376
rect 233417 133318 286015 133320
rect 233417 133315 233483 133318
rect 285949 133315 286015 133318
rect 101397 133242 101463 133245
rect 282269 133242 282335 133245
rect 101397 133240 282335 133242
rect 101397 133184 101402 133240
rect 101458 133184 282274 133240
rect 282330 133184 282335 133240
rect 101397 133182 282335 133184
rect 101397 133179 101463 133182
rect 282269 133179 282335 133182
rect 3366 133044 3372 133108
rect 3436 133106 3442 133108
rect 283230 133106 283236 133108
rect 3436 133046 283236 133106
rect 3436 133044 3442 133046
rect 283230 133044 283236 133046
rect 283300 133044 283306 133108
rect 208577 132018 208643 132021
rect 284753 132018 284819 132021
rect 208577 132016 284819 132018
rect 208577 131960 208582 132016
rect 208638 131960 284758 132016
rect 284814 131960 284819 132016
rect 208577 131958 284819 131960
rect 208577 131955 208643 131958
rect 284753 131955 284819 131958
rect 197905 131882 197971 131885
rect 284845 131882 284911 131885
rect 197905 131880 284911 131882
rect 197905 131824 197910 131880
rect 197966 131824 284850 131880
rect 284906 131824 284911 131880
rect 197905 131822 284911 131824
rect 197905 131819 197971 131822
rect 284845 131819 284911 131822
rect 103329 131746 103395 131749
rect 286317 131746 286383 131749
rect 103329 131744 286383 131746
rect 103329 131688 103334 131744
rect 103390 131688 286322 131744
rect 286378 131688 286383 131744
rect 103329 131686 286383 131688
rect 103329 131683 103395 131686
rect 286317 131683 286383 131686
rect 141233 130522 141299 130525
rect 280838 130522 280844 130524
rect 141233 130520 280844 130522
rect 141233 130464 141238 130520
rect 141294 130464 280844 130520
rect 141233 130462 280844 130464
rect 141233 130459 141299 130462
rect 280838 130460 280844 130462
rect 280908 130460 280914 130524
rect 89161 130386 89227 130389
rect 286409 130386 286475 130389
rect 89161 130384 286475 130386
rect 89161 130328 89166 130384
rect 89222 130328 286414 130384
rect 286470 130328 286475 130384
rect 89161 130326 286475 130328
rect 89161 130323 89227 130326
rect 286409 130323 286475 130326
rect 190821 129298 190887 129301
rect 283281 129298 283347 129301
rect 190821 129296 283347 129298
rect 190821 129240 190826 129296
rect 190882 129240 283286 129296
rect 283342 129240 283347 129296
rect 190821 129238 283347 129240
rect 190821 129235 190887 129238
rect 283281 129235 283347 129238
rect 151813 129162 151879 129165
rect 280613 129162 280679 129165
rect 151813 129160 280679 129162
rect 151813 129104 151818 129160
rect 151874 129104 280618 129160
rect 280674 129104 280679 129160
rect 151813 129102 280679 129104
rect 151813 129099 151879 129102
rect 280613 129099 280679 129102
rect 85665 129026 85731 129029
rect 286501 129026 286567 129029
rect 85665 129024 286567 129026
rect 85665 128968 85670 129024
rect 85726 128968 286506 129024
rect 286562 128968 286567 129024
rect 85665 128966 286567 128968
rect 85665 128963 85731 128966
rect 286501 128963 286567 128966
rect 130561 127802 130627 127805
rect 281942 127802 281948 127804
rect 130561 127800 281948 127802
rect 130561 127744 130566 127800
rect 130622 127744 281948 127800
rect 130561 127742 281948 127744
rect 130561 127739 130627 127742
rect 281942 127740 281948 127742
rect 282012 127740 282018 127804
rect 14733 127666 14799 127669
rect 281022 127666 281028 127668
rect 14733 127664 281028 127666
rect 14733 127608 14738 127664
rect 14794 127608 281028 127664
rect 14733 127606 281028 127608
rect 14733 127603 14799 127606
rect 281022 127604 281028 127606
rect 281092 127604 281098 127668
rect 212165 126442 212231 126445
rect 284661 126442 284727 126445
rect 212165 126440 284727 126442
rect 212165 126384 212170 126440
rect 212226 126384 284666 126440
rect 284722 126384 284727 126440
rect 212165 126382 284727 126384
rect 212165 126379 212231 126382
rect 284661 126379 284727 126382
rect 11697 126306 11763 126309
rect 282126 126306 282132 126308
rect 11697 126304 282132 126306
rect 11697 126248 11702 126304
rect 11758 126248 282132 126304
rect 11697 126246 282132 126248
rect 11697 126243 11763 126246
rect 282126 126244 282132 126246
rect 282196 126244 282202 126308
rect 583520 125884 584960 126124
rect 45461 124946 45527 124949
rect 191097 124946 191163 124949
rect 45461 124944 191163 124946
rect 45461 124888 45466 124944
rect 45522 124888 191102 124944
rect 191158 124888 191163 124944
rect 45461 124886 191163 124888
rect 45461 124883 45527 124886
rect 191097 124883 191163 124886
rect 222745 124946 222811 124949
rect 284477 124946 284543 124949
rect 222745 124944 284543 124946
rect 222745 124888 222750 124944
rect 222806 124888 284482 124944
rect 284538 124888 284543 124944
rect 222745 124886 284543 124888
rect 222745 124883 222811 124886
rect 284477 124883 284543 124886
rect 92749 124810 92815 124813
rect 286225 124810 286291 124813
rect 92749 124808 286291 124810
rect 92749 124752 92754 124808
rect 92810 124752 286230 124808
rect 286286 124752 286291 124808
rect 92749 124750 286291 124752
rect 92749 124747 92815 124750
rect 286225 124747 286291 124750
rect -960 123572 480 123812
rect 91553 123586 91619 123589
rect 211797 123586 211863 123589
rect 91553 123584 211863 123586
rect 91553 123528 91558 123584
rect 91614 123528 211802 123584
rect 211858 123528 211863 123584
rect 91553 123526 211863 123528
rect 91553 123523 91619 123526
rect 211797 123523 211863 123526
rect 226333 123586 226399 123589
rect 283097 123586 283163 123589
rect 226333 123584 283163 123586
rect 226333 123528 226338 123584
rect 226394 123528 283102 123584
rect 283158 123528 283163 123584
rect 226333 123526 283163 123528
rect 226333 123523 226399 123526
rect 283097 123523 283163 123526
rect 114001 123450 114067 123453
rect 286041 123450 286107 123453
rect 114001 123448 286107 123450
rect 114001 123392 114006 123448
rect 114062 123392 286046 123448
rect 286102 123392 286107 123448
rect 114001 123390 286107 123392
rect 114001 123387 114067 123390
rect 286041 123387 286107 123390
rect 18229 122226 18295 122229
rect 215937 122226 216003 122229
rect 18229 122224 216003 122226
rect 18229 122168 18234 122224
rect 18290 122168 215942 122224
rect 215998 122168 216003 122224
rect 18229 122166 216003 122168
rect 18229 122163 18295 122166
rect 215937 122163 216003 122166
rect 43069 122090 43135 122093
rect 287789 122090 287855 122093
rect 43069 122088 287855 122090
rect 43069 122032 43074 122088
rect 43130 122032 287794 122088
rect 287850 122032 287855 122088
rect 43069 122030 287855 122032
rect 43069 122027 43135 122030
rect 287789 122027 287855 122030
rect 98637 120866 98703 120869
rect 226977 120866 227043 120869
rect 98637 120864 227043 120866
rect 98637 120808 98642 120864
rect 98698 120808 226982 120864
rect 227038 120808 227043 120864
rect 98637 120806 227043 120808
rect 98637 120803 98703 120806
rect 226977 120803 227043 120806
rect 35985 120730 36051 120733
rect 287697 120730 287763 120733
rect 35985 120728 287763 120730
rect 35985 120672 35990 120728
rect 36046 120672 287702 120728
rect 287758 120672 287763 120728
rect 35985 120670 287763 120672
rect 35985 120667 36051 120670
rect 287697 120667 287763 120670
rect 134149 119506 134215 119509
rect 285029 119506 285095 119509
rect 134149 119504 285095 119506
rect 134149 119448 134154 119504
rect 134210 119448 285034 119504
rect 285090 119448 285095 119504
rect 134149 119446 285095 119448
rect 134149 119443 134215 119446
rect 285029 119443 285095 119446
rect 96245 119370 96311 119373
rect 286133 119370 286199 119373
rect 96245 119368 286199 119370
rect 96245 119312 96250 119368
rect 96306 119312 286138 119368
rect 286194 119312 286199 119368
rect 96245 119310 286199 119312
rect 96245 119307 96311 119310
rect 286133 119307 286199 119310
rect 137645 118146 137711 118149
rect 281758 118146 281764 118148
rect 137645 118144 281764 118146
rect 137645 118088 137650 118144
rect 137706 118088 281764 118144
rect 137645 118086 281764 118088
rect 137645 118083 137711 118086
rect 281758 118084 281764 118086
rect 281828 118084 281834 118148
rect 93945 118010 94011 118013
rect 268929 118010 268995 118013
rect 93945 118008 268995 118010
rect 93945 117952 93950 118008
rect 94006 117952 268934 118008
rect 268990 117952 268995 118008
rect 93945 117950 268995 117952
rect 93945 117947 94011 117950
rect 268929 117947 268995 117950
rect 148317 116650 148383 116653
rect 281901 116650 281967 116653
rect 148317 116648 281967 116650
rect 148317 116592 148322 116648
rect 148378 116592 281906 116648
rect 281962 116592 281967 116648
rect 148317 116590 281967 116592
rect 148317 116587 148383 116590
rect 281901 116587 281967 116590
rect 19425 116514 19491 116517
rect 279366 116514 279372 116516
rect 19425 116512 279372 116514
rect 19425 116456 19430 116512
rect 19486 116456 279372 116512
rect 19425 116454 279372 116456
rect 19425 116451 19491 116454
rect 279366 116452 279372 116454
rect 279436 116452 279442 116516
rect 24209 115154 24275 115157
rect 283414 115154 283420 115156
rect 24209 115152 283420 115154
rect 24209 115096 24214 115152
rect 24270 115096 283420 115152
rect 24209 115094 283420 115096
rect 24209 115091 24275 115094
rect 283414 115092 283420 115094
rect 283484 115092 283490 115156
rect 38377 113794 38443 113797
rect 144177 113794 144243 113797
rect 38377 113792 144243 113794
rect 38377 113736 38382 113792
rect 38438 113736 144182 113792
rect 144238 113736 144243 113792
rect 38377 113734 144243 113736
rect 38377 113731 38443 113734
rect 144177 113731 144243 113734
rect 239806 112780 239812 112844
rect 239876 112842 239882 112844
rect 583520 112842 584960 112932
rect 239876 112782 584960 112842
rect 239876 112780 239882 112782
rect 583520 112692 584960 112782
rect 35249 112434 35315 112437
rect 238017 112434 238083 112437
rect 35249 112432 238083 112434
rect 35249 112376 35254 112432
rect 35310 112376 238022 112432
rect 238078 112376 238083 112432
rect 35249 112374 238083 112376
rect 35249 112371 35315 112374
rect 238017 112371 238083 112374
rect 41873 111074 41939 111077
rect 152457 111074 152523 111077
rect 41873 111072 152523 111074
rect 41873 111016 41878 111072
rect 41934 111016 152462 111072
rect 152518 111016 152523 111072
rect 41873 111014 152523 111016
rect 41873 111011 41939 111014
rect 152457 111011 152523 111014
rect 155401 111074 155467 111077
rect 283189 111074 283255 111077
rect 155401 111072 283255 111074
rect 155401 111016 155406 111072
rect 155462 111016 283194 111072
rect 283250 111016 283255 111072
rect 155401 111014 283255 111016
rect 155401 111011 155467 111014
rect 283189 111011 283255 111014
rect -960 110666 480 110756
rect 47577 110666 47643 110669
rect -960 110664 47643 110666
rect -960 110608 47582 110664
rect 47638 110608 47643 110664
rect -960 110606 47643 110608
rect -960 110516 480 110606
rect 47577 110603 47643 110606
rect 34789 109714 34855 109717
rect 155217 109714 155283 109717
rect 34789 109712 155283 109714
rect 34789 109656 34794 109712
rect 34850 109656 155222 109712
rect 155278 109656 155283 109712
rect 34789 109654 155283 109656
rect 34789 109651 34855 109654
rect 155217 109651 155283 109654
rect 158897 109714 158963 109717
rect 284385 109714 284451 109717
rect 158897 109712 284451 109714
rect 158897 109656 158902 109712
rect 158958 109656 284390 109712
rect 284446 109656 284451 109712
rect 158897 109654 284451 109656
rect 158897 109651 158963 109654
rect 284385 109651 284451 109654
rect 110505 108490 110571 108493
rect 281993 108490 282059 108493
rect 110505 108488 282059 108490
rect 110505 108432 110510 108488
rect 110566 108432 281998 108488
rect 282054 108432 282059 108488
rect 110505 108430 282059 108432
rect 110505 108427 110571 108430
rect 281993 108427 282059 108430
rect 90357 108354 90423 108357
rect 267733 108354 267799 108357
rect 90357 108352 267799 108354
rect 90357 108296 90362 108352
rect 90418 108296 267738 108352
rect 267794 108296 267799 108352
rect 90357 108294 267799 108296
rect 90357 108291 90423 108294
rect 267733 108291 267799 108294
rect 97441 106858 97507 106861
rect 270125 106858 270191 106861
rect 97441 106856 270191 106858
rect 97441 106800 97446 106856
rect 97502 106800 270130 106856
rect 270186 106800 270191 106856
rect 97441 106798 270191 106800
rect 97441 106795 97507 106798
rect 270125 106795 270191 106798
rect 104525 105498 104591 105501
rect 271137 105498 271203 105501
rect 104525 105496 271203 105498
rect 104525 105440 104530 105496
rect 104586 105440 271142 105496
rect 271198 105440 271203 105496
rect 104525 105438 271203 105440
rect 104525 105435 104591 105438
rect 271137 105435 271203 105438
rect 122281 104274 122347 104277
rect 278497 104274 278563 104277
rect 122281 104272 278563 104274
rect 122281 104216 122286 104272
rect 122342 104216 278502 104272
rect 278558 104216 278563 104272
rect 122281 104214 278563 104216
rect 122281 104211 122347 104214
rect 278497 104211 278563 104214
rect 39573 104138 39639 104141
rect 287605 104138 287671 104141
rect 39573 104136 287671 104138
rect 39573 104080 39578 104136
rect 39634 104080 287610 104136
rect 287666 104080 287671 104136
rect 39573 104078 287671 104080
rect 39573 104075 39639 104078
rect 287605 104075 287671 104078
rect 119889 102914 119955 102917
rect 197997 102914 198063 102917
rect 119889 102912 198063 102914
rect 119889 102856 119894 102912
rect 119950 102856 198002 102912
rect 198058 102856 198063 102912
rect 119889 102854 198063 102856
rect 119889 102851 119955 102854
rect 197997 102851 198063 102854
rect 99833 102778 99899 102781
rect 280061 102778 280127 102781
rect 99833 102776 280127 102778
rect 99833 102720 99838 102776
rect 99894 102720 280066 102776
rect 280122 102720 280127 102776
rect 99833 102718 280127 102720
rect 99833 102715 99899 102718
rect 280061 102715 280127 102718
rect 102225 101554 102291 101557
rect 209037 101554 209103 101557
rect 102225 101552 209103 101554
rect 102225 101496 102230 101552
rect 102286 101496 209042 101552
rect 209098 101496 209103 101552
rect 102225 101494 209103 101496
rect 102225 101491 102291 101494
rect 209037 101491 209103 101494
rect 32397 101418 32463 101421
rect 287881 101418 287947 101421
rect 32397 101416 287947 101418
rect 32397 101360 32402 101416
rect 32458 101360 287886 101416
rect 287942 101360 287947 101416
rect 32397 101358 287947 101360
rect 32397 101355 32463 101358
rect 287881 101355 287947 101358
rect 124673 100194 124739 100197
rect 287513 100194 287579 100197
rect 124673 100192 287579 100194
rect 124673 100136 124678 100192
rect 124734 100136 287518 100192
rect 287574 100136 287579 100192
rect 124673 100134 287579 100136
rect 124673 100131 124739 100134
rect 287513 100131 287579 100134
rect 13537 100058 13603 100061
rect 203517 100058 203583 100061
rect 13537 100056 203583 100058
rect 13537 100000 13542 100056
rect 13598 100000 203522 100056
rect 203578 100000 203583 100056
rect 13537 99998 203583 100000
rect 13537 99995 13603 99998
rect 203517 99995 203583 99998
rect 306966 99452 306972 99516
rect 307036 99514 307042 99516
rect 583520 99514 584960 99604
rect 307036 99454 584960 99514
rect 307036 99452 307042 99454
rect 583520 99364 584960 99454
rect 106917 98834 106983 98837
rect 284569 98834 284635 98837
rect 106917 98832 284635 98834
rect 106917 98776 106922 98832
rect 106978 98776 284574 98832
rect 284630 98776 284635 98832
rect 106917 98774 284635 98776
rect 106917 98771 106983 98774
rect 284569 98771 284635 98774
rect 8753 98698 8819 98701
rect 195237 98698 195303 98701
rect 8753 98696 195303 98698
rect 8753 98640 8758 98696
rect 8814 98640 195242 98696
rect 195298 98640 195303 98696
rect 8753 98638 195303 98640
rect 8753 98635 8819 98638
rect 195237 98635 195303 98638
rect -960 97610 480 97700
rect 3366 97610 3372 97612
rect -960 97550 3372 97610
rect -960 97460 480 97550
rect 3366 97548 3372 97550
rect 3436 97548 3442 97612
rect 111609 97338 111675 97341
rect 274909 97338 274975 97341
rect 111609 97336 274975 97338
rect 111609 97280 111614 97336
rect 111670 97280 274914 97336
rect 274970 97280 274975 97336
rect 111609 97278 274975 97280
rect 111609 97275 111675 97278
rect 274909 97275 274975 97278
rect 46657 97202 46723 97205
rect 281574 97202 281580 97204
rect 46657 97200 281580 97202
rect 46657 97144 46662 97200
rect 46718 97144 281580 97200
rect 46657 97142 281580 97144
rect 46657 97139 46723 97142
rect 281574 97140 281580 97142
rect 281644 97140 281650 97204
rect 108113 95842 108179 95845
rect 273713 95842 273779 95845
rect 108113 95840 273779 95842
rect 108113 95784 108118 95840
rect 108174 95784 273718 95840
rect 273774 95784 273779 95840
rect 108113 95782 273779 95784
rect 108113 95779 108179 95782
rect 273713 95779 273779 95782
rect 101029 94482 101095 94485
rect 271321 94482 271387 94485
rect 101029 94480 271387 94482
rect 101029 94424 101034 94480
rect 101090 94424 271326 94480
rect 271382 94424 271387 94480
rect 101029 94422 271387 94424
rect 101029 94419 101095 94422
rect 271321 94419 271387 94422
rect 86861 93122 86927 93125
rect 266537 93122 266603 93125
rect 86861 93120 266603 93122
rect 86861 93064 86866 93120
rect 86922 93064 266542 93120
rect 266598 93064 266603 93120
rect 86861 93062 266603 93064
rect 86861 93059 86927 93062
rect 266537 93059 266603 93062
rect 2865 91762 2931 91765
rect 222837 91762 222903 91765
rect 2865 91760 222903 91762
rect 2865 91704 2870 91760
rect 2926 91704 222842 91760
rect 222898 91704 222903 91760
rect 2865 91702 222903 91704
rect 2865 91699 2931 91702
rect 222837 91699 222903 91702
rect 87689 90538 87755 90541
rect 213177 90538 213243 90541
rect 87689 90536 213243 90538
rect 87689 90480 87694 90536
rect 87750 90480 213182 90536
rect 213238 90480 213243 90536
rect 87689 90478 213243 90480
rect 87689 90475 87755 90478
rect 213177 90475 213243 90478
rect 121085 90402 121151 90405
rect 287421 90402 287487 90405
rect 121085 90400 287487 90402
rect 121085 90344 121090 90400
rect 121146 90344 287426 90400
rect 287482 90344 287487 90400
rect 121085 90342 287487 90344
rect 121085 90339 121151 90342
rect 287421 90339 287487 90342
rect 3734 88980 3740 89044
rect 3804 89042 3810 89044
rect 283046 89042 283052 89044
rect 3804 88982 283052 89042
rect 3804 88980 3810 88982
rect 283046 88980 283052 88982
rect 283116 88980 283122 89044
rect 288934 88980 288940 89044
rect 289004 89042 289010 89044
rect 580206 89042 580212 89044
rect 289004 88982 580212 89042
rect 289004 88980 289010 88982
rect 580206 88980 580212 88982
rect 580276 88980 580282 89044
rect 65609 87954 65675 87957
rect 91737 87954 91803 87957
rect 65609 87952 91803 87954
rect 65609 87896 65614 87952
rect 65670 87896 91742 87952
rect 91798 87896 91803 87952
rect 65609 87894 91803 87896
rect 65609 87891 65675 87894
rect 91737 87891 91803 87894
rect 52913 87818 52979 87821
rect 86217 87818 86283 87821
rect 52913 87816 86283 87818
rect 52913 87760 52918 87816
rect 52974 87760 86222 87816
rect 86278 87760 86283 87816
rect 52913 87758 86283 87760
rect 52913 87755 52979 87758
rect 86217 87755 86283 87758
rect 60641 87682 60707 87685
rect 84837 87682 84903 87685
rect 60641 87680 84903 87682
rect 60641 87624 60646 87680
rect 60702 87624 84842 87680
rect 84898 87624 84903 87680
rect 60641 87622 84903 87624
rect 60641 87619 60707 87622
rect 84837 87619 84903 87622
rect 62021 87546 62087 87549
rect 87781 87546 87847 87549
rect 62021 87544 87847 87546
rect 62021 87488 62026 87544
rect 62082 87488 87786 87544
rect 87842 87488 87847 87544
rect 62021 87486 87847 87488
rect 62021 87483 62087 87486
rect 87781 87483 87847 87486
rect 57605 87410 57671 87413
rect 85021 87410 85087 87413
rect 57605 87408 85087 87410
rect 57605 87352 57610 87408
rect 57666 87352 85026 87408
rect 85082 87352 85087 87408
rect 57605 87350 85087 87352
rect 57605 87347 57671 87350
rect 85021 87347 85087 87350
rect 59261 87274 59327 87277
rect 91921 87274 91987 87277
rect 59261 87272 91987 87274
rect 59261 87216 59266 87272
rect 59322 87216 91926 87272
rect 91982 87216 91987 87272
rect 59261 87214 91987 87216
rect 59261 87211 59327 87214
rect 91921 87211 91987 87214
rect 54661 87138 54727 87141
rect 87597 87138 87663 87141
rect 54661 87136 87663 87138
rect 54661 87080 54666 87136
rect 54722 87080 87602 87136
rect 87658 87080 87663 87136
rect 54661 87078 87663 87080
rect 54661 87075 54727 87078
rect 87597 87075 87663 87078
rect 3366 86260 3372 86324
rect 3436 86322 3442 86324
rect 228214 86322 228220 86324
rect 3436 86262 228220 86322
rect 3436 86260 3442 86262
rect 228214 86260 228220 86262
rect 228284 86260 228290 86324
rect 56501 86186 56567 86189
rect 311433 86186 311499 86189
rect 56501 86184 311499 86186
rect 56501 86128 56506 86184
rect 56562 86128 311438 86184
rect 311494 86128 311499 86184
rect 56501 86126 311499 86128
rect 56501 86123 56567 86126
rect 311433 86123 311499 86126
rect 492581 86186 492647 86189
rect 583520 86186 584960 86276
rect 492581 86184 584960 86186
rect 492581 86128 492586 86184
rect 492642 86128 584960 86184
rect 492581 86126 584960 86128
rect 492581 86123 492647 86126
rect 583520 86036 584960 86126
rect 68645 85914 68711 85917
rect 273897 85914 273963 85917
rect 68645 85912 273963 85914
rect 68645 85856 68650 85912
rect 68706 85856 273902 85912
rect 273958 85856 273963 85912
rect 68645 85854 273963 85856
rect 68645 85851 68711 85854
rect 273897 85851 273963 85854
rect 50981 85778 51047 85781
rect 271137 85778 271203 85781
rect 50981 85776 271203 85778
rect 50981 85720 50986 85776
rect 51042 85720 271142 85776
rect 271198 85720 271203 85776
rect 50981 85718 271203 85720
rect 50981 85715 51047 85718
rect 271137 85715 271203 85718
rect 63861 85642 63927 85645
rect 329189 85642 329255 85645
rect 63861 85640 329255 85642
rect 63861 85584 63866 85640
rect 63922 85584 329194 85640
rect 329250 85584 329255 85640
rect 63861 85582 329255 85584
rect 63861 85579 63927 85582
rect 329189 85579 329255 85582
rect 80743 84962 80809 84965
rect 364609 84962 364675 84965
rect 80743 84960 364675 84962
rect 80743 84904 80748 84960
rect 80804 84904 364614 84960
rect 364670 84904 364675 84960
rect 80743 84902 364675 84904
rect 80743 84899 80809 84902
rect 364609 84899 364675 84902
rect 77615 84826 77681 84829
rect 357525 84826 357591 84829
rect 77615 84824 357591 84826
rect -960 84690 480 84780
rect 77615 84768 77620 84824
rect 77676 84768 357530 84824
rect 357586 84768 357591 84824
rect 77615 84766 357591 84768
rect 77615 84763 77681 84766
rect 357525 84763 357591 84766
rect 3366 84690 3372 84692
rect -960 84630 3372 84690
rect -960 84540 480 84630
rect 3366 84628 3372 84630
rect 3436 84628 3442 84692
rect 71359 84690 71425 84693
rect 343357 84690 343423 84693
rect 71359 84688 343423 84690
rect 71359 84632 71364 84688
rect 71420 84632 343362 84688
rect 343418 84632 343423 84688
rect 71359 84630 343423 84632
rect 71359 84627 71425 84630
rect 343357 84627 343423 84630
rect 79179 84554 79245 84557
rect 361113 84554 361179 84557
rect 79179 84552 361179 84554
rect 79179 84496 79184 84552
rect 79240 84496 361118 84552
rect 361174 84496 361179 84552
rect 79179 84494 361179 84496
rect 79179 84491 79245 84494
rect 361113 84491 361179 84494
rect 432597 83058 432663 83061
rect 84916 83056 432663 83058
rect 84916 83000 432602 83056
rect 432658 83000 432663 83056
rect 84916 82998 432663 83000
rect 432597 82995 432663 82998
rect 48221 81698 48287 81701
rect 428549 81698 428615 81701
rect 48221 81696 50140 81698
rect 48221 81640 48226 81696
rect 48282 81640 50140 81696
rect 48221 81638 50140 81640
rect 84916 81696 428615 81698
rect 84916 81640 428554 81696
rect 428610 81640 428615 81696
rect 84916 81638 428615 81640
rect 48221 81635 48287 81638
rect 428549 81635 428615 81638
rect 85021 80746 85087 80749
rect 315021 80746 315087 80749
rect 85021 80744 315087 80746
rect 85021 80688 85026 80744
rect 85082 80688 315026 80744
rect 315082 80688 315087 80744
rect 85021 80686 315087 80688
rect 85021 80683 85087 80686
rect 315021 80683 315087 80686
rect 47853 80338 47919 80341
rect 105537 80338 105603 80341
rect 47853 80336 50140 80338
rect 47853 80280 47858 80336
rect 47914 80280 50140 80336
rect 47853 80278 50140 80280
rect 84916 80336 105603 80338
rect 84916 80280 105542 80336
rect 105598 80280 105603 80336
rect 84916 80278 105603 80280
rect 47853 80275 47919 80278
rect 105537 80275 105603 80278
rect 84837 79386 84903 79389
rect 322105 79386 322171 79389
rect 84837 79384 322171 79386
rect 84837 79328 84842 79384
rect 84898 79328 322110 79384
rect 322166 79328 322171 79384
rect 84837 79326 322171 79328
rect 84837 79323 84903 79326
rect 322105 79323 322171 79326
rect 49417 78978 49483 78981
rect 421557 78978 421623 78981
rect 49417 78976 50140 78978
rect 49417 78920 49422 78976
rect 49478 78920 50140 78976
rect 49417 78918 50140 78920
rect 84916 78976 421623 78978
rect 84916 78920 421562 78976
rect 421618 78920 421623 78976
rect 84916 78918 421623 78920
rect 49417 78915 49483 78918
rect 421557 78915 421623 78918
rect 49325 77618 49391 77621
rect 417417 77618 417483 77621
rect 49325 77616 50140 77618
rect 49325 77560 49330 77616
rect 49386 77560 50140 77616
rect 49325 77558 50140 77560
rect 84916 77616 417483 77618
rect 84916 77560 417422 77616
rect 417478 77560 417483 77616
rect 84916 77558 417483 77560
rect 49325 77555 49391 77558
rect 417417 77555 417483 77558
rect 414657 76258 414723 76261
rect 84916 76256 414723 76258
rect 50478 75989 50538 76228
rect 84916 76200 414662 76256
rect 414718 76200 414723 76256
rect 84916 76198 414723 76200
rect 414657 76195 414723 76198
rect 50429 75984 50538 75989
rect 50429 75928 50434 75984
rect 50490 75928 50538 75984
rect 50429 75926 50538 75928
rect 50429 75923 50495 75926
rect 49601 74898 49667 74901
rect 410517 74898 410583 74901
rect 49601 74896 50140 74898
rect 49601 74840 49606 74896
rect 49662 74840 50140 74896
rect 49601 74838 50140 74840
rect 84916 74896 410583 74898
rect 84916 74840 410522 74896
rect 410578 74840 410583 74896
rect 84916 74838 410583 74840
rect 49601 74835 49667 74838
rect 410517 74835 410583 74838
rect 450537 73538 450603 73541
rect 84916 73536 450603 73538
rect 50478 73269 50538 73508
rect 84916 73480 450542 73536
rect 450598 73480 450603 73536
rect 84916 73478 450603 73480
rect 450537 73475 450603 73478
rect 50478 73264 50587 73269
rect 50478 73208 50526 73264
rect 50582 73208 50587 73264
rect 50478 73206 50587 73208
rect 50521 73203 50587 73206
rect 580257 72994 580323 72997
rect 583520 72994 584960 73084
rect 580257 72992 584960 72994
rect 580257 72936 580262 72992
rect 580318 72936 584960 72992
rect 580257 72934 584960 72936
rect 580257 72931 580323 72934
rect 583520 72844 584960 72934
rect 49509 72178 49575 72181
rect 446397 72178 446463 72181
rect 49509 72176 50140 72178
rect 49509 72120 49514 72176
rect 49570 72120 50140 72176
rect 49509 72118 50140 72120
rect 84916 72176 446463 72178
rect 84916 72120 446402 72176
rect 446458 72120 446463 72176
rect 84916 72118 446463 72120
rect 49509 72115 49575 72118
rect 446397 72115 446463 72118
rect -960 71634 480 71724
rect 35157 71634 35223 71637
rect -960 71632 35223 71634
rect -960 71576 35162 71632
rect 35218 71576 35223 71632
rect -960 71574 35223 71576
rect -960 71484 480 71574
rect 35157 71571 35223 71574
rect 443637 70818 443703 70821
rect 84916 70816 443703 70818
rect 50110 70413 50170 70788
rect 84916 70760 443642 70816
rect 443698 70760 443703 70816
rect 84916 70758 443703 70760
rect 443637 70755 443703 70758
rect 50110 70408 50219 70413
rect 50110 70352 50158 70408
rect 50214 70352 50219 70408
rect 50110 70350 50219 70352
rect 50153 70347 50219 70350
rect 49233 69458 49299 69461
rect 258717 69458 258783 69461
rect 49233 69456 50140 69458
rect 49233 69400 49238 69456
rect 49294 69400 50140 69456
rect 49233 69398 50140 69400
rect 84916 69456 258783 69458
rect 84916 69400 258722 69456
rect 258778 69400 258783 69456
rect 84916 69398 258783 69400
rect 49233 69395 49299 69398
rect 258717 69395 258783 69398
rect 49141 68098 49207 68101
rect 425697 68098 425763 68101
rect 49141 68096 50140 68098
rect 49141 68040 49146 68096
rect 49202 68040 50140 68096
rect 49141 68038 50140 68040
rect 84916 68096 425763 68098
rect 84916 68040 425702 68096
rect 425758 68040 425763 68096
rect 84916 68038 425763 68040
rect 49141 68035 49207 68038
rect 425697 68035 425763 68038
rect 436737 66738 436803 66741
rect 84916 66736 436803 66738
rect 50294 66333 50354 66708
rect 84916 66680 436742 66736
rect 436798 66680 436803 66736
rect 84916 66678 436803 66680
rect 436737 66675 436803 66678
rect 50245 66328 50354 66333
rect 50245 66272 50250 66328
rect 50306 66272 50354 66328
rect 50245 66270 50354 66272
rect 50245 66267 50311 66270
rect 48129 65378 48195 65381
rect 431217 65378 431283 65381
rect 48129 65376 50140 65378
rect 48129 65320 48134 65376
rect 48190 65320 50140 65376
rect 48129 65318 50140 65320
rect 84916 65376 431283 65378
rect 84916 65320 431222 65376
rect 431278 65320 431283 65376
rect 84916 65318 431283 65320
rect 48129 65315 48195 65318
rect 431217 65315 431283 65318
rect 47485 64018 47551 64021
rect 429837 64018 429903 64021
rect 47485 64016 50140 64018
rect 47485 63960 47490 64016
rect 47546 63960 50140 64016
rect 47485 63958 50140 63960
rect 84916 64016 429903 64018
rect 84916 63960 429842 64016
rect 429898 63960 429903 64016
rect 84916 63958 429903 63960
rect 47485 63955 47551 63958
rect 429837 63955 429903 63958
rect 48037 62658 48103 62661
rect 427077 62658 427143 62661
rect 48037 62656 50140 62658
rect 48037 62600 48042 62656
rect 48098 62600 50140 62656
rect 48037 62598 50140 62600
rect 84916 62656 427143 62658
rect 84916 62600 427082 62656
rect 427138 62600 427143 62656
rect 84916 62598 427143 62600
rect 48037 62595 48103 62598
rect 427077 62595 427143 62598
rect 47577 61298 47643 61301
rect 422937 61298 423003 61301
rect 47577 61296 50140 61298
rect 47577 61240 47582 61296
rect 47638 61240 50140 61296
rect 47577 61238 50140 61240
rect 84916 61296 423003 61298
rect 84916 61240 422942 61296
rect 422998 61240 423003 61296
rect 84916 61238 423003 61240
rect 47577 61235 47643 61238
rect 422937 61235 423003 61238
rect 47945 59938 48011 59941
rect 418797 59938 418863 59941
rect 47945 59936 50140 59938
rect 47945 59880 47950 59936
rect 48006 59880 50140 59936
rect 47945 59878 50140 59880
rect 84916 59936 418863 59938
rect 84916 59880 418802 59936
rect 418858 59880 418863 59936
rect 84916 59878 418863 59880
rect 47945 59875 48011 59878
rect 418797 59875 418863 59878
rect 580206 59604 580212 59668
rect 580276 59666 580282 59668
rect 583520 59666 584960 59756
rect 580276 59606 584960 59666
rect 580276 59604 580282 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3366 58578 3372 58580
rect -960 58518 3372 58578
rect -960 58428 480 58518
rect 3366 58516 3372 58518
rect 3436 58516 3442 58580
rect 47761 58578 47827 58581
rect 334617 58578 334683 58581
rect 47761 58576 50140 58578
rect 47761 58520 47766 58576
rect 47822 58520 50140 58576
rect 47761 58518 50140 58520
rect 84916 58576 334683 58578
rect 84916 58520 334622 58576
rect 334678 58520 334683 58576
rect 84916 58518 334683 58520
rect 47761 58515 47827 58518
rect 334617 58515 334683 58518
rect 47669 57218 47735 57221
rect 411897 57218 411963 57221
rect 47669 57216 50140 57218
rect 47669 57160 47674 57216
rect 47730 57160 50140 57216
rect 47669 57158 50140 57160
rect 84916 57216 411963 57218
rect 84916 57160 411902 57216
rect 411958 57160 411963 57216
rect 84916 57158 411963 57160
rect 47669 57155 47735 57158
rect 411897 57155 411963 57158
rect 49049 55858 49115 55861
rect 355317 55858 355383 55861
rect 49049 55856 50140 55858
rect 49049 55800 49054 55856
rect 49110 55800 50140 55856
rect 49049 55798 50140 55800
rect 84916 55856 355383 55858
rect 84916 55800 355322 55856
rect 355378 55800 355383 55856
rect 84916 55798 355383 55800
rect 49049 55795 49115 55798
rect 355317 55795 355383 55798
rect 87781 54634 87847 54637
rect 325601 54634 325667 54637
rect 87781 54632 325667 54634
rect 87781 54576 87786 54632
rect 87842 54576 325606 54632
rect 325662 54576 325667 54632
rect 87781 54574 325667 54576
rect 87781 54571 87847 54574
rect 325601 54571 325667 54574
rect 260097 54498 260163 54501
rect 84916 54496 260163 54498
rect 50478 53954 50538 54468
rect 84916 54440 260102 54496
rect 260158 54440 260163 54496
rect 84916 54438 260163 54440
rect 260097 54435 260163 54438
rect 50613 53954 50679 53957
rect 50478 53952 50679 53954
rect 50478 53896 50618 53952
rect 50674 53896 50679 53952
rect 50478 53894 50679 53896
rect 50613 53891 50679 53894
rect 84653 53274 84719 53277
rect 188337 53274 188403 53277
rect 84653 53272 188403 53274
rect 84653 53216 84658 53272
rect 84714 53216 188342 53272
rect 188398 53216 188403 53272
rect 84653 53214 188403 53216
rect 84653 53211 84719 53214
rect 188337 53211 188403 53214
rect 91921 53138 91987 53141
rect 318517 53138 318583 53141
rect 91921 53136 318583 53138
rect 50110 52597 50170 53108
rect 91921 53080 91926 53136
rect 91982 53080 318522 53136
rect 318578 53080 318583 53136
rect 91921 53078 318583 53080
rect 91921 53075 91987 53078
rect 318517 53075 318583 53078
rect 50061 52592 50170 52597
rect 50061 52536 50066 52592
rect 50122 52536 50170 52592
rect 50061 52534 50170 52536
rect 84886 52594 84946 53040
rect 87045 52594 87111 52597
rect 87689 52594 87755 52597
rect 84886 52592 87755 52594
rect 84886 52536 87050 52592
rect 87106 52536 87694 52592
rect 87750 52536 87755 52592
rect 84886 52534 87755 52536
rect 50061 52531 50127 52534
rect 87045 52531 87111 52534
rect 87689 52531 87755 52534
rect 86217 51914 86283 51917
rect 304349 51914 304415 51917
rect 86217 51912 304415 51914
rect 86217 51856 86222 51912
rect 86278 51856 304354 51912
rect 304410 51856 304415 51912
rect 86217 51854 304415 51856
rect 86217 51851 86283 51854
rect 304349 51851 304415 51854
rect 86953 51778 87019 51781
rect 88241 51778 88307 51781
rect 84916 51776 88307 51778
rect 84916 51720 86958 51776
rect 87014 51720 88246 51776
rect 88302 51720 88307 51776
rect 84916 51718 88307 51720
rect 86953 51715 87019 51718
rect 88241 51715 88307 51718
rect 105537 51778 105603 51781
rect 471053 51778 471119 51781
rect 105537 51776 471119 51778
rect 105537 51720 105542 51776
rect 105598 51720 471058 51776
rect 471114 51720 471119 51776
rect 105537 51718 471119 51720
rect 105537 51715 105603 51718
rect 471053 51715 471119 51718
rect 67909 50282 67975 50285
rect 284293 50282 284359 50285
rect 67909 50280 284359 50282
rect 67909 50224 67914 50280
rect 67970 50224 284298 50280
rect 284354 50224 284359 50280
rect 67909 50222 284359 50224
rect 67909 50219 67975 50222
rect 284293 50219 284359 50222
rect 71497 49330 71563 49333
rect 280654 49330 280660 49332
rect 71497 49328 280660 49330
rect 71497 49272 71502 49328
rect 71558 49272 280660 49328
rect 71497 49270 280660 49272
rect 71497 49267 71563 49270
rect 280654 49268 280660 49270
rect 280724 49268 280730 49332
rect 50337 49194 50403 49197
rect 289813 49194 289879 49197
rect 50337 49192 289879 49194
rect 50337 49136 50342 49192
rect 50398 49136 289818 49192
rect 289874 49136 289879 49192
rect 50337 49134 289879 49136
rect 50337 49131 50403 49134
rect 289813 49131 289879 49134
rect 48221 49058 48287 49061
rect 289077 49058 289143 49061
rect 48221 49056 289143 49058
rect 48221 49000 48226 49056
rect 48282 49000 289082 49056
rect 289138 49000 289143 49056
rect 48221 48998 289143 49000
rect 48221 48995 48287 48998
rect 289077 48995 289143 48998
rect 49325 48922 49391 48925
rect 545481 48922 545547 48925
rect 49325 48920 545547 48922
rect 49325 48864 49330 48920
rect 49386 48864 545486 48920
rect 545542 48864 545547 48920
rect 49325 48862 545547 48864
rect 49325 48859 49391 48862
rect 545481 48859 545547 48862
rect 77201 48106 77267 48109
rect 79317 48106 79383 48109
rect 77201 48104 79383 48106
rect 77201 48048 77206 48104
rect 77262 48048 79322 48104
rect 79378 48048 79383 48104
rect 77201 48046 79383 48048
rect 77201 48043 77267 48046
rect 79317 48043 79383 48046
rect 60641 47970 60707 47973
rect 62757 47970 62823 47973
rect 60641 47968 62823 47970
rect 60641 47912 60646 47968
rect 60702 47912 62762 47968
rect 62818 47912 62823 47968
rect 60641 47910 62823 47912
rect 60641 47907 60707 47910
rect 62757 47907 62823 47910
rect 78581 47970 78647 47973
rect 79501 47970 79567 47973
rect 78581 47968 79567 47970
rect 78581 47912 78586 47968
rect 78642 47912 79506 47968
rect 79562 47912 79567 47968
rect 78581 47910 79567 47912
rect 78581 47907 78647 47910
rect 79501 47907 79567 47910
rect 84101 47970 84167 47973
rect 87689 47970 87755 47973
rect 84101 47968 87755 47970
rect 84101 47912 84106 47968
rect 84162 47912 87694 47968
rect 87750 47912 87755 47968
rect 84101 47910 87755 47912
rect 84101 47907 84167 47910
rect 87689 47907 87755 47910
rect 50981 47834 51047 47837
rect 435357 47834 435423 47837
rect 50981 47832 435423 47834
rect 50981 47776 50986 47832
rect 51042 47776 435362 47832
rect 435418 47776 435423 47832
rect 50981 47774 435423 47776
rect 50981 47771 51047 47774
rect 435357 47771 435423 47774
rect 52361 47698 52427 47701
rect 439497 47698 439563 47701
rect 52361 47696 439563 47698
rect 52361 47640 52366 47696
rect 52422 47640 439502 47696
rect 439558 47640 439563 47696
rect 52361 47638 439563 47640
rect 52361 47635 52427 47638
rect 439497 47635 439563 47638
rect 53741 47562 53807 47565
rect 442257 47562 442323 47565
rect 53741 47560 442323 47562
rect 53741 47504 53746 47560
rect 53802 47504 442262 47560
rect 442318 47504 442323 47560
rect 53741 47502 442323 47504
rect 53741 47499 53807 47502
rect 442257 47499 442323 47502
rect 64781 47018 64847 47021
rect 65609 47018 65675 47021
rect 64781 47016 65675 47018
rect 64781 46960 64786 47016
rect 64842 46960 65614 47016
rect 65670 46960 65675 47016
rect 64781 46958 65675 46960
rect 64781 46955 64847 46958
rect 65609 46955 65675 46958
rect 74441 47018 74507 47021
rect 75177 47018 75243 47021
rect 74441 47016 75243 47018
rect 74441 46960 74446 47016
rect 74502 46960 75182 47016
rect 75238 46960 75243 47016
rect 74441 46958 75243 46960
rect 74441 46955 74507 46958
rect 75177 46955 75243 46958
rect 47853 46338 47919 46341
rect 267181 46338 267247 46341
rect 47853 46336 267247 46338
rect 47853 46280 47858 46336
rect 47914 46280 267186 46336
rect 267242 46280 267247 46336
rect 47853 46278 267247 46280
rect 47853 46275 47919 46278
rect 267181 46275 267247 46278
rect 490414 46276 490420 46340
rect 490484 46338 490490 46340
rect 583520 46338 584960 46428
rect 490484 46278 584960 46338
rect 490484 46276 490490 46278
rect 56501 46202 56567 46205
rect 481725 46202 481791 46205
rect 56501 46200 481791 46202
rect 56501 46144 56506 46200
rect 56562 46144 481730 46200
rect 481786 46144 481791 46200
rect 583520 46188 584960 46278
rect 56501 46142 481791 46144
rect 56501 46139 56567 46142
rect 481725 46139 481791 46142
rect -960 45522 480 45612
rect 219934 45522 219940 45524
rect -960 45462 219940 45522
rect -960 45372 480 45462
rect 219934 45460 219940 45462
rect 220004 45460 220010 45524
rect 60825 44978 60891 44981
rect 284518 44978 284524 44980
rect 60825 44976 284524 44978
rect 60825 44920 60830 44976
rect 60886 44920 284524 44976
rect 60825 44918 284524 44920
rect 60825 44915 60891 44918
rect 284518 44916 284524 44918
rect 284588 44916 284594 44980
rect 49417 44842 49483 44845
rect 549069 44842 549135 44845
rect 49417 44840 549135 44842
rect 49417 44784 49422 44840
rect 49478 44784 549074 44840
rect 549130 44784 549135 44840
rect 49417 44782 549135 44784
rect 49417 44779 49483 44782
rect 549069 44779 549135 44782
rect 48129 43618 48195 43621
rect 282177 43618 282243 43621
rect 48129 43616 282243 43618
rect 48129 43560 48134 43616
rect 48190 43560 282182 43616
rect 282238 43560 282243 43616
rect 48129 43558 282243 43560
rect 48129 43555 48195 43558
rect 282177 43555 282243 43558
rect 63309 43482 63375 43485
rect 499389 43482 499455 43485
rect 63309 43480 499455 43482
rect 63309 43424 63314 43480
rect 63370 43424 499394 43480
rect 499450 43424 499455 43480
rect 63309 43422 499455 43424
rect 63309 43419 63375 43422
rect 499389 43419 499455 43422
rect 50061 42258 50127 42261
rect 297265 42258 297331 42261
rect 50061 42256 297331 42258
rect 50061 42200 50066 42256
rect 50122 42200 297270 42256
rect 297326 42200 297331 42256
rect 50061 42198 297331 42200
rect 50061 42195 50127 42198
rect 297265 42195 297331 42198
rect 66069 42122 66135 42125
rect 506473 42122 506539 42125
rect 66069 42120 506539 42122
rect 66069 42064 66074 42120
rect 66130 42064 506478 42120
rect 506534 42064 506539 42120
rect 66069 42062 506539 42064
rect 66069 42059 66135 42062
rect 506473 42059 506539 42062
rect 81249 40762 81315 40765
rect 400121 40762 400187 40765
rect 81249 40760 400187 40762
rect 81249 40704 81254 40760
rect 81310 40704 400126 40760
rect 400182 40704 400187 40760
rect 81249 40702 400187 40704
rect 81249 40699 81315 40702
rect 400121 40699 400187 40702
rect 68829 40626 68895 40629
rect 512637 40626 512703 40629
rect 68829 40624 512703 40626
rect 68829 40568 68834 40624
rect 68890 40568 512642 40624
rect 512698 40568 512703 40624
rect 68829 40566 512703 40568
rect 68829 40563 68895 40566
rect 512637 40563 512703 40566
rect 82997 39402 83063 39405
rect 403617 39402 403683 39405
rect 82997 39400 403683 39402
rect 82997 39344 83002 39400
rect 83058 39344 403622 39400
rect 403678 39344 403683 39400
rect 82997 39342 403683 39344
rect 82997 39339 83063 39342
rect 403617 39339 403683 39342
rect 49141 39266 49207 39269
rect 520733 39266 520799 39269
rect 49141 39264 520799 39266
rect 49141 39208 49146 39264
rect 49202 39208 520738 39264
rect 520794 39208 520799 39264
rect 49141 39206 520799 39208
rect 49141 39203 49207 39206
rect 520733 39203 520799 39206
rect 51349 38178 51415 38181
rect 254577 38178 254643 38181
rect 51349 38176 254643 38178
rect 51349 38120 51354 38176
rect 51410 38120 254582 38176
rect 254638 38120 254643 38176
rect 51349 38118 254643 38120
rect 51349 38115 51415 38118
rect 254577 38115 254643 38118
rect 74993 38042 75059 38045
rect 285622 38042 285628 38044
rect 74993 38040 285628 38042
rect 74993 37984 74998 38040
rect 75054 37984 285628 38040
rect 74993 37982 285628 37984
rect 74993 37979 75059 37982
rect 285622 37980 285628 37982
rect 285692 37980 285698 38044
rect 49233 37906 49299 37909
rect 524229 37906 524295 37909
rect 49233 37904 524295 37906
rect 49233 37848 49238 37904
rect 49294 37848 524234 37904
rect 524290 37848 524295 37904
rect 49233 37846 524295 37848
rect 49233 37843 49299 37846
rect 524229 37843 524295 37846
rect 65517 36682 65583 36685
rect 259361 36682 259427 36685
rect 65517 36680 259427 36682
rect 65517 36624 65522 36680
rect 65578 36624 259366 36680
rect 259422 36624 259427 36680
rect 65517 36622 259427 36624
rect 65517 36619 65583 36622
rect 259361 36619 259427 36622
rect 49509 36546 49575 36549
rect 531313 36546 531379 36549
rect 49509 36544 531379 36546
rect 49509 36488 49514 36544
rect 49570 36488 531318 36544
rect 531374 36488 531379 36544
rect 49509 36486 531379 36488
rect 49509 36483 49575 36486
rect 531313 36483 531379 36486
rect 83273 35322 83339 35325
rect 265341 35322 265407 35325
rect 83273 35320 265407 35322
rect 83273 35264 83278 35320
rect 83334 35264 265346 35320
rect 265402 35264 265407 35320
rect 83273 35262 265407 35264
rect 83273 35259 83339 35262
rect 265341 35259 265407 35262
rect 50521 35186 50587 35189
rect 534901 35186 534967 35189
rect 50521 35184 534967 35186
rect 50521 35128 50526 35184
rect 50582 35128 534906 35184
rect 534962 35128 534967 35184
rect 50521 35126 534967 35128
rect 50521 35123 50587 35126
rect 534901 35123 534967 35126
rect 69105 33962 69171 33965
rect 260557 33962 260623 33965
rect 69105 33960 260623 33962
rect 69105 33904 69110 33960
rect 69166 33904 260562 33960
rect 260618 33904 260623 33960
rect 69105 33902 260623 33904
rect 69105 33899 69171 33902
rect 260557 33899 260623 33902
rect 49601 33826 49667 33829
rect 538397 33826 538463 33829
rect 49601 33824 538463 33826
rect 49601 33768 49606 33824
rect 49662 33768 538402 33824
rect 538458 33768 538463 33824
rect 49601 33766 538463 33768
rect 49601 33763 49667 33766
rect 538397 33763 538463 33766
rect 239857 33146 239923 33149
rect 583520 33146 584960 33236
rect 239857 33144 584960 33146
rect 239857 33088 239862 33144
rect 239918 33088 584960 33144
rect 239857 33086 584960 33088
rect 239857 33083 239923 33086
rect 583520 32996 584960 33086
rect 4889 32874 4955 32877
rect 87045 32874 87111 32877
rect 4889 32872 87111 32874
rect 4889 32816 4894 32872
rect 4950 32816 87050 32872
rect 87106 32816 87111 32872
rect 4889 32814 87111 32816
rect 4889 32811 4955 32814
rect 87045 32811 87111 32814
rect 59629 32738 59695 32741
rect 199377 32738 199443 32741
rect 59629 32736 199443 32738
rect 59629 32680 59634 32736
rect 59690 32680 199382 32736
rect 199438 32680 199443 32736
rect 59629 32678 199443 32680
rect 59629 32675 59695 32678
rect 199377 32675 199443 32678
rect 82077 32602 82143 32605
rect 285765 32602 285831 32605
rect 82077 32600 285831 32602
rect -960 32466 480 32556
rect 82077 32544 82082 32600
rect 82138 32544 285770 32600
rect 285826 32544 285831 32600
rect 82077 32542 285831 32544
rect 82077 32539 82143 32542
rect 285765 32539 285831 32542
rect 4797 32466 4863 32469
rect -960 32464 4863 32466
rect -960 32408 4802 32464
rect 4858 32408 4863 32464
rect -960 32406 4863 32408
rect -960 32316 480 32406
rect 4797 32403 4863 32406
rect 70209 32466 70275 32469
rect 278037 32466 278103 32469
rect 70209 32464 278103 32466
rect 70209 32408 70214 32464
rect 70270 32408 278042 32464
rect 278098 32408 278103 32464
rect 70209 32406 278103 32408
rect 70209 32403 70275 32406
rect 278037 32403 278103 32406
rect 56041 31242 56107 31245
rect 146937 31242 147003 31245
rect 56041 31240 147003 31242
rect 56041 31184 56046 31240
rect 56102 31184 146942 31240
rect 146998 31184 147003 31240
rect 56041 31182 147003 31184
rect 56041 31179 56107 31182
rect 146937 31179 147003 31182
rect 70301 31106 70367 31109
rect 214557 31106 214623 31109
rect 70301 31104 214623 31106
rect 70301 31048 70306 31104
rect 70362 31048 214562 31104
rect 214618 31048 214623 31104
rect 70301 31046 214623 31048
rect 70301 31043 70367 31046
rect 214557 31043 214623 31046
rect 50429 30970 50495 30973
rect 541985 30970 542051 30973
rect 50429 30968 542051 30970
rect 50429 30912 50434 30968
rect 50490 30912 541990 30968
rect 542046 30912 542051 30968
rect 50429 30910 542051 30912
rect 50429 30907 50495 30910
rect 541985 30907 542051 30910
rect 52545 29882 52611 29885
rect 174537 29882 174603 29885
rect 52545 29880 174603 29882
rect 52545 29824 52550 29880
rect 52606 29824 174542 29880
rect 174598 29824 174603 29880
rect 52545 29822 174603 29824
rect 52545 29819 52611 29822
rect 174537 29819 174603 29822
rect 80881 29746 80947 29749
rect 210417 29746 210483 29749
rect 80881 29744 210483 29746
rect 80881 29688 80886 29744
rect 80942 29688 210422 29744
rect 210478 29688 210483 29744
rect 80881 29686 210483 29688
rect 80881 29683 80947 29686
rect 210417 29683 210483 29686
rect 50613 29610 50679 29613
rect 552657 29610 552723 29613
rect 50613 29608 552723 29610
rect 50613 29552 50618 29608
rect 50674 29552 552662 29608
rect 552718 29552 552723 29608
rect 50613 29550 552723 29552
rect 50613 29547 50679 29550
rect 552657 29547 552723 29550
rect 48957 28522 49023 28525
rect 138657 28522 138723 28525
rect 48957 28520 138723 28522
rect 48957 28464 48962 28520
rect 49018 28464 138662 28520
rect 138718 28464 138723 28520
rect 48957 28462 138723 28464
rect 48957 28459 49023 28462
rect 138657 28459 138723 28462
rect 63217 28386 63283 28389
rect 231117 28386 231183 28389
rect 63217 28384 231183 28386
rect 63217 28328 63222 28384
rect 63278 28328 231122 28384
rect 231178 28328 231183 28384
rect 63217 28326 231183 28328
rect 63217 28323 63283 28326
rect 231117 28323 231183 28326
rect 47669 28250 47735 28253
rect 559741 28250 559807 28253
rect 47669 28248 559807 28250
rect 47669 28192 47674 28248
rect 47730 28192 559746 28248
rect 559802 28192 559807 28248
rect 47669 28190 559807 28192
rect 47669 28187 47735 28190
rect 559741 28187 559807 28190
rect 4061 27026 4127 27029
rect 178677 27026 178743 27029
rect 4061 27024 178743 27026
rect 4061 26968 4066 27024
rect 4122 26968 178682 27024
rect 178738 26968 178743 27024
rect 4061 26966 178743 26968
rect 4061 26963 4127 26966
rect 178677 26963 178743 26966
rect 47761 26890 47827 26893
rect 562317 26890 562383 26893
rect 47761 26888 562383 26890
rect 47761 26832 47766 26888
rect 47822 26832 562322 26888
rect 562378 26832 562383 26888
rect 47761 26830 562383 26832
rect 47761 26827 47827 26830
rect 562317 26827 562383 26830
rect 58433 25666 58499 25669
rect 256969 25666 257035 25669
rect 58433 25664 257035 25666
rect 58433 25608 58438 25664
rect 58494 25608 256974 25664
rect 257030 25608 257035 25664
rect 58433 25606 257035 25608
rect 58433 25603 58499 25606
rect 256969 25603 257035 25606
rect 47945 25530 48011 25533
rect 566825 25530 566891 25533
rect 47945 25528 566891 25530
rect 47945 25472 47950 25528
rect 48006 25472 566830 25528
rect 566886 25472 566891 25528
rect 47945 25470 566891 25472
rect 47945 25467 48011 25470
rect 566825 25467 566891 25470
rect 79501 24306 79567 24309
rect 393037 24306 393103 24309
rect 79501 24304 393103 24306
rect 79501 24248 79506 24304
rect 79562 24248 393042 24304
rect 393098 24248 393103 24304
rect 79501 24246 393103 24248
rect 79501 24243 79567 24246
rect 393037 24243 393103 24246
rect 49049 24170 49115 24173
rect 556153 24170 556219 24173
rect 49049 24168 556219 24170
rect 49049 24112 49054 24168
rect 49110 24112 556158 24168
rect 556214 24112 556219 24168
rect 49049 24110 556219 24112
rect 49049 24107 49115 24110
rect 556153 24107 556219 24110
rect 62021 22810 62087 22813
rect 258165 22810 258231 22813
rect 62021 22808 258231 22810
rect 62021 22752 62026 22808
rect 62082 22752 258170 22808
rect 258226 22752 258231 22808
rect 62021 22750 258231 22752
rect 62021 22747 62087 22750
rect 258165 22747 258231 22750
rect 48037 22674 48103 22677
rect 573909 22674 573975 22677
rect 48037 22672 573975 22674
rect 48037 22616 48042 22672
rect 48098 22616 573914 22672
rect 573970 22616 573975 22672
rect 48037 22614 573975 22616
rect 48037 22611 48103 22614
rect 573909 22611 573975 22614
rect 54937 21586 55003 21589
rect 255773 21586 255839 21589
rect 54937 21584 255839 21586
rect 54937 21528 54942 21584
rect 54998 21528 255778 21584
rect 255834 21528 255839 21584
rect 54937 21526 255839 21528
rect 54937 21523 55003 21526
rect 255773 21523 255839 21526
rect 78581 21450 78647 21453
rect 285673 21450 285739 21453
rect 78581 21448 285739 21450
rect 78581 21392 78586 21448
rect 78642 21392 285678 21448
rect 285734 21392 285739 21448
rect 78581 21390 285739 21392
rect 78581 21387 78647 21390
rect 285673 21387 285739 21390
rect 47577 21314 47643 21317
rect 570321 21314 570387 21317
rect 47577 21312 570387 21314
rect 47577 21256 47582 21312
rect 47638 21256 570326 21312
rect 570382 21256 570387 21312
rect 47577 21254 570387 21256
rect 47577 21251 47643 21254
rect 570321 21251 570387 21254
rect 75177 20090 75243 20093
rect 382365 20090 382431 20093
rect 75177 20088 382431 20090
rect 75177 20032 75182 20088
rect 75238 20032 382370 20088
rect 382426 20032 382431 20088
rect 75177 20030 382431 20032
rect 75177 20027 75243 20030
rect 382365 20027 382431 20030
rect 65609 19954 65675 19957
rect 502977 19954 503043 19957
rect 65609 19952 503043 19954
rect 65609 19896 65614 19952
rect 65670 19896 502982 19952
rect 503038 19896 503043 19952
rect 65609 19894 503043 19896
rect 65609 19891 65675 19894
rect 502977 19891 503043 19894
rect 551134 19756 551140 19820
rect 551204 19818 551210 19820
rect 583520 19818 584960 19908
rect 551204 19758 584960 19818
rect 551204 19756 551210 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 288750 19410 288756 19412
rect -960 19350 288756 19410
rect -960 19260 480 19350
rect 288750 19348 288756 19350
rect 288820 19348 288826 19412
rect 87689 18730 87755 18733
rect 407205 18730 407271 18733
rect 87689 18728 407271 18730
rect 87689 18672 87694 18728
rect 87750 18672 407210 18728
rect 407266 18672 407271 18728
rect 87689 18670 407271 18672
rect 87689 18667 87755 18670
rect 407205 18667 407271 18670
rect 50153 18594 50219 18597
rect 527817 18594 527883 18597
rect 50153 18592 527883 18594
rect 50153 18536 50158 18592
rect 50214 18536 527822 18592
rect 527878 18536 527883 18592
rect 50153 18534 527883 18536
rect 50153 18531 50219 18534
rect 527817 18531 527883 18534
rect 80697 17370 80763 17373
rect 396533 17370 396599 17373
rect 80697 17368 396599 17370
rect 80697 17312 80702 17368
rect 80758 17312 396538 17368
rect 396594 17312 396599 17368
rect 80697 17310 396599 17312
rect 80697 17307 80763 17310
rect 396533 17307 396599 17310
rect 50245 17234 50311 17237
rect 517145 17234 517211 17237
rect 50245 17232 517211 17234
rect 50245 17176 50250 17232
rect 50306 17176 517150 17232
rect 517206 17176 517211 17232
rect 50245 17174 517211 17176
rect 50245 17171 50311 17174
rect 517145 17171 517211 17174
rect 79317 16010 79383 16013
rect 389449 16010 389515 16013
rect 79317 16008 389515 16010
rect 79317 15952 79322 16008
rect 79378 15952 389454 16008
rect 389510 15952 389515 16008
rect 79317 15950 389515 15952
rect 79317 15947 79383 15950
rect 389449 15947 389515 15950
rect 47485 15874 47551 15877
rect 576117 15874 576183 15877
rect 47485 15872 576183 15874
rect 47485 15816 47490 15872
rect 47546 15816 576122 15872
rect 576178 15816 576183 15872
rect 47485 15814 576183 15816
rect 47485 15811 47551 15814
rect 576117 15811 576183 15814
rect 57237 14786 57303 14789
rect 283005 14786 283071 14789
rect 57237 14784 283071 14786
rect 57237 14728 57242 14784
rect 57298 14728 283010 14784
rect 283066 14728 283071 14784
rect 57237 14726 283071 14728
rect 57237 14723 57303 14726
rect 283005 14723 283071 14726
rect 76557 14650 76623 14653
rect 385953 14650 386019 14653
rect 76557 14648 386019 14650
rect 76557 14592 76562 14648
rect 76618 14592 385958 14648
rect 386014 14592 386019 14648
rect 76557 14590 386019 14592
rect 76557 14587 76623 14590
rect 385953 14587 386019 14590
rect 67449 14514 67515 14517
rect 508497 14514 508563 14517
rect 67449 14512 508563 14514
rect 67449 14456 67454 14512
rect 67510 14456 508502 14512
rect 508558 14456 508563 14512
rect 67449 14454 508563 14456
rect 67449 14451 67515 14454
rect 508497 14451 508563 14454
rect 72969 13154 73035 13157
rect 378869 13154 378935 13157
rect 72969 13152 378935 13154
rect 72969 13096 72974 13152
rect 73030 13096 378874 13152
rect 378930 13096 378935 13152
rect 72969 13094 378935 13096
rect 72969 13091 73035 13094
rect 378869 13091 378935 13094
rect 61929 13018 61995 13021
rect 495893 13018 495959 13021
rect 61929 13016 495959 13018
rect 61929 12960 61934 13016
rect 61990 12960 495898 13016
rect 495954 12960 495959 13016
rect 61929 12958 495959 12960
rect 61929 12955 61995 12958
rect 495893 12955 495959 12958
rect 72417 11794 72483 11797
rect 375281 11794 375347 11797
rect 72417 11792 375347 11794
rect 72417 11736 72422 11792
rect 72478 11736 375286 11792
rect 375342 11736 375347 11792
rect 72417 11734 375347 11736
rect 72417 11731 72483 11734
rect 375281 11731 375347 11734
rect 62757 11658 62823 11661
rect 492305 11658 492371 11661
rect 62757 11656 492371 11658
rect 62757 11600 62762 11656
rect 62818 11600 492310 11656
rect 492366 11600 492371 11656
rect 62757 11598 492371 11600
rect 62757 11595 62823 11598
rect 492305 11595 492371 11598
rect 66713 10434 66779 10437
rect 140037 10434 140103 10437
rect 66713 10432 140103 10434
rect 66713 10376 66718 10432
rect 66774 10376 140042 10432
rect 140098 10376 140103 10432
rect 66713 10374 140103 10376
rect 66713 10371 66779 10374
rect 140037 10371 140103 10374
rect 59169 10298 59235 10301
rect 488809 10298 488875 10301
rect 59169 10296 488875 10298
rect 59169 10240 59174 10296
rect 59230 10240 488814 10296
rect 488870 10240 488875 10296
rect 59169 10238 488875 10240
rect 59169 10235 59235 10238
rect 488809 10235 488875 10238
rect 87965 9210 88031 9213
rect 126237 9210 126303 9213
rect 87965 9208 126303 9210
rect 87965 9152 87970 9208
rect 88026 9152 126242 9208
rect 126298 9152 126303 9208
rect 87965 9150 126303 9152
rect 87965 9147 88031 9150
rect 126237 9147 126303 9150
rect 55029 9074 55095 9077
rect 290181 9074 290247 9077
rect 55029 9072 290247 9074
rect 55029 9016 55034 9072
rect 55090 9016 290186 9072
rect 290242 9016 290247 9072
rect 55029 9014 290247 9016
rect 55029 9011 55095 9014
rect 290181 9011 290247 9014
rect 57789 8938 57855 8941
rect 485221 8938 485287 8941
rect 57789 8936 485287 8938
rect 57789 8880 57794 8936
rect 57850 8880 485226 8936
rect 485282 8880 485287 8936
rect 57789 8878 485287 8880
rect 57789 8875 57855 8878
rect 485221 8875 485287 8878
rect 73797 7850 73863 7853
rect 151077 7850 151143 7853
rect 73797 7848 151143 7850
rect 73797 7792 73802 7848
rect 73858 7792 151082 7848
rect 151138 7792 151143 7848
rect 73797 7790 151143 7792
rect 73797 7787 73863 7790
rect 151077 7787 151143 7790
rect 4102 7652 4108 7716
rect 4172 7714 4178 7716
rect 224166 7714 224172 7716
rect 4172 7654 224172 7714
rect 4172 7652 4178 7654
rect 224166 7652 224172 7654
rect 224236 7652 224242 7716
rect 91737 7578 91803 7581
rect 332685 7578 332751 7581
rect 91737 7576 332751 7578
rect 91737 7520 91742 7576
rect 91798 7520 332690 7576
rect 332746 7520 332751 7576
rect 91737 7518 332751 7520
rect 91737 7515 91803 7518
rect 332685 7515 332751 7518
rect 334617 7578 334683 7581
rect 417877 7578 417943 7581
rect 334617 7576 417943 7578
rect 334617 7520 334622 7576
rect 334678 7520 417882 7576
rect 417938 7520 417943 7576
rect 334617 7518 417943 7520
rect 334617 7515 334683 7518
rect 417877 7515 417943 7518
rect 425697 7578 425763 7581
rect 442625 7578 442691 7581
rect 425697 7576 442691 7578
rect 425697 7520 425702 7576
rect 425758 7520 442630 7576
rect 442686 7520 442691 7576
rect 425697 7518 442691 7520
rect 425697 7515 425763 7518
rect 442625 7515 442691 7518
rect 79685 6762 79751 6765
rect 264145 6762 264211 6765
rect 79685 6760 264211 6762
rect 79685 6704 79690 6760
rect 79746 6704 264150 6760
rect 264206 6704 264211 6760
rect 79685 6702 264211 6704
rect 79685 6699 79751 6702
rect 264145 6699 264211 6702
rect 76189 6626 76255 6629
rect 262949 6626 263015 6629
rect 76189 6624 263015 6626
rect -960 6490 480 6580
rect 76189 6568 76194 6624
rect 76250 6568 262954 6624
rect 263010 6568 263015 6624
rect 76189 6566 263015 6568
rect 76189 6563 76255 6566
rect 262949 6563 263015 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 4102 6490 4108 6492
rect -960 6430 4108 6490
rect -960 6340 480 6430
rect 4102 6428 4108 6430
rect 4172 6428 4178 6492
rect 72601 6490 72667 6493
rect 261661 6490 261727 6493
rect 72601 6488 261727 6490
rect 72601 6432 72606 6488
rect 72662 6432 261666 6488
rect 261722 6432 261727 6488
rect 583520 6476 584960 6566
rect 72601 6430 261727 6432
rect 72601 6427 72667 6430
rect 261661 6427 261727 6430
rect 47853 6354 47919 6357
rect 253381 6354 253447 6357
rect 47853 6352 253447 6354
rect 47853 6296 47858 6352
rect 47914 6296 253386 6352
rect 253442 6296 253447 6352
rect 47853 6294 253447 6296
rect 47853 6291 47919 6294
rect 253381 6291 253447 6294
rect 12341 6218 12407 6221
rect 242617 6218 242683 6221
rect 12341 6216 242683 6218
rect 12341 6160 12346 6216
rect 12402 6160 242622 6216
rect 242678 6160 242683 6216
rect 12341 6158 242683 6160
rect 12341 6155 12407 6158
rect 242617 6155 242683 6158
rect 258717 6218 258783 6221
rect 286593 6218 286659 6221
rect 258717 6216 286659 6218
rect 258717 6160 258722 6216
rect 258778 6160 286598 6216
rect 286654 6160 286659 6216
rect 258717 6158 286659 6160
rect 258717 6155 258783 6158
rect 286593 6155 286659 6158
rect 77385 5130 77451 5133
rect 142797 5130 142863 5133
rect 77385 5128 142863 5130
rect 77385 5072 77390 5128
rect 77446 5072 142802 5128
rect 142858 5072 142863 5128
rect 77385 5070 142863 5072
rect 77385 5067 77451 5070
rect 142797 5067 142863 5070
rect 87597 4994 87663 4997
rect 307937 4994 308003 4997
rect 87597 4992 308003 4994
rect 87597 4936 87602 4992
rect 87658 4936 307942 4992
rect 307998 4936 308003 4992
rect 87597 4934 308003 4936
rect 87597 4931 87663 4934
rect 307937 4931 308003 4934
rect 431217 4994 431283 4997
rect 435541 4994 435607 4997
rect 431217 4992 435607 4994
rect 431217 4936 431222 4992
rect 431278 4936 435546 4992
rect 435602 4936 435607 4992
rect 431217 4934 435607 4936
rect 431217 4931 431283 4934
rect 435541 4931 435607 4934
rect 7649 4858 7715 4861
rect 241421 4858 241487 4861
rect 7649 4856 241487 4858
rect 7649 4800 7654 4856
rect 7710 4800 241426 4856
rect 241482 4800 241487 4856
rect 7649 4798 241487 4800
rect 7649 4795 7715 4798
rect 241421 4795 241487 4798
rect 260097 4858 260163 4861
rect 283097 4858 283163 4861
rect 260097 4856 283163 4858
rect 260097 4800 260102 4856
rect 260158 4800 283102 4856
rect 283158 4800 283163 4856
rect 260097 4798 283163 4800
rect 260097 4795 260163 4798
rect 283097 4795 283163 4798
rect 355317 4858 355383 4861
rect 410793 4858 410859 4861
rect 355317 4856 410859 4858
rect 355317 4800 355322 4856
rect 355378 4800 410798 4856
rect 410854 4800 410859 4856
rect 355317 4798 410859 4800
rect 355317 4795 355383 4798
rect 410793 4795 410859 4798
rect 411897 4858 411963 4861
rect 414289 4858 414355 4861
rect 411897 4856 414355 4858
rect 411897 4800 411902 4856
rect 411958 4800 414294 4856
rect 414350 4800 414355 4856
rect 411897 4798 414355 4800
rect 411897 4795 411963 4798
rect 414289 4795 414355 4798
rect 429837 4858 429903 4861
rect 432045 4858 432111 4861
rect 429837 4856 432111 4858
rect 429837 4800 429842 4856
rect 429898 4800 432050 4856
rect 432106 4800 432111 4856
rect 429837 4798 432111 4800
rect 429837 4795 429903 4798
rect 432045 4795 432111 4798
rect 450537 4858 450603 4861
rect 453297 4858 453363 4861
rect 450537 4856 453363 4858
rect 450537 4800 450542 4856
rect 450598 4800 453302 4856
rect 453358 4800 453363 4856
rect 450537 4798 453363 4800
rect 450537 4795 450603 4798
rect 453297 4795 453363 4798
rect 418797 4178 418863 4181
rect 421373 4178 421439 4181
rect 418797 4176 421439 4178
rect 418797 4120 418802 4176
rect 418858 4120 421378 4176
rect 421434 4120 421439 4176
rect 418797 4118 421439 4120
rect 418797 4115 418863 4118
rect 421373 4115 421439 4118
rect 422937 4178 423003 4181
rect 424961 4178 425027 4181
rect 422937 4176 425027 4178
rect 422937 4120 422942 4176
rect 422998 4120 424966 4176
rect 425022 4120 425027 4176
rect 422937 4118 425027 4120
rect 422937 4115 423003 4118
rect 424961 4115 425027 4118
rect 427077 4178 427143 4181
rect 428457 4178 428523 4181
rect 427077 4176 428523 4178
rect 427077 4120 427082 4176
rect 427138 4120 428462 4176
rect 428518 4120 428523 4176
rect 427077 4118 428523 4120
rect 427077 4115 427143 4118
rect 428457 4115 428523 4118
rect 436737 4178 436803 4181
rect 439129 4178 439195 4181
rect 436737 4176 439195 4178
rect 436737 4120 436742 4176
rect 436798 4120 439134 4176
rect 439190 4120 439195 4176
rect 436737 4118 439195 4120
rect 436737 4115 436803 4118
rect 439129 4115 439195 4118
rect 443637 4178 443703 4181
rect 446213 4178 446279 4181
rect 443637 4176 446279 4178
rect 443637 4120 443642 4176
rect 443698 4120 446218 4176
rect 446274 4120 446279 4176
rect 443637 4118 446279 4120
rect 443637 4115 443703 4118
rect 446213 4115 446279 4118
rect 446397 4178 446463 4181
rect 449801 4178 449867 4181
rect 446397 4176 449867 4178
rect 446397 4120 446402 4176
rect 446458 4120 449806 4176
rect 449862 4120 449867 4176
rect 446397 4118 449867 4120
rect 446397 4115 446463 4118
rect 449801 4115 449867 4118
rect 267181 4042 267247 4045
rect 268837 4042 268903 4045
rect 267181 4040 268903 4042
rect 267181 3984 267186 4040
rect 267242 3984 268842 4040
rect 268898 3984 268903 4040
rect 267181 3982 268903 3984
rect 267181 3979 267247 3982
rect 268837 3979 268903 3982
rect 277853 4042 277919 4045
rect 281349 4042 281415 4045
rect 277853 4040 281415 4042
rect 277853 3984 277858 4040
rect 277914 3984 281354 4040
rect 281410 3984 281415 4040
rect 277853 3982 281415 3984
rect 277853 3979 277919 3982
rect 281349 3979 281415 3982
rect 435357 4042 435423 4045
rect 438853 4042 438919 4045
rect 435357 4040 438919 4042
rect 435357 3984 435362 4040
rect 435418 3984 438858 4040
rect 438914 3984 438919 4040
rect 435357 3982 438919 3984
rect 435357 3979 435423 3982
rect 438853 3979 438919 3982
rect 508497 4042 508563 4045
rect 510061 4042 510127 4045
rect 508497 4040 510127 4042
rect 508497 3984 508502 4040
rect 508558 3984 510066 4040
rect 510122 3984 510127 4040
rect 508497 3982 510127 3984
rect 508497 3979 508563 3982
rect 510061 3979 510127 3982
rect 576117 4042 576183 4045
rect 577405 4042 577471 4045
rect 576117 4040 577471 4042
rect 576117 3984 576122 4040
rect 576178 3984 577410 4040
rect 577466 3984 577471 4040
rect 576117 3982 577471 3984
rect 576117 3979 576183 3982
rect 577405 3979 577471 3982
rect 237005 3906 237071 3909
rect 280981 3906 281047 3909
rect 237005 3904 281047 3906
rect 237005 3848 237010 3904
rect 237066 3848 280986 3904
rect 281042 3848 281047 3904
rect 237005 3846 281047 3848
rect 237005 3843 237071 3846
rect 280981 3843 281047 3846
rect 421557 3906 421623 3909
rect 467465 3906 467531 3909
rect 421557 3904 467531 3906
rect 421557 3848 421562 3904
rect 421618 3848 467470 3904
rect 467526 3848 467531 3904
rect 421557 3846 467531 3848
rect 421557 3843 421623 3846
rect 467465 3843 467531 3846
rect 15837 3770 15903 3773
rect 6870 3768 15903 3770
rect 6870 3712 15842 3768
rect 15898 3712 15903 3768
rect 6870 3710 15903 3712
rect 1669 3498 1735 3501
rect 4889 3498 4955 3501
rect 1669 3496 4955 3498
rect 1669 3440 1674 3496
rect 1730 3440 4894 3496
rect 4950 3440 4955 3496
rect 1669 3438 4955 3440
rect 1669 3435 1735 3438
rect 4889 3435 4955 3438
rect 6453 3498 6519 3501
rect 6870 3498 6930 3710
rect 15837 3707 15903 3710
rect 205081 3770 205147 3773
rect 206277 3770 206343 3773
rect 205081 3768 206343 3770
rect 205081 3712 205086 3768
rect 205142 3712 206282 3768
rect 206338 3712 206343 3768
rect 205081 3710 206343 3712
rect 205081 3707 205147 3710
rect 206277 3707 206343 3710
rect 229829 3770 229895 3773
rect 280797 3770 280863 3773
rect 229829 3768 280863 3770
rect 229829 3712 229834 3768
rect 229890 3712 280802 3768
rect 280858 3712 280863 3768
rect 229829 3710 280863 3712
rect 229829 3707 229895 3710
rect 280797 3707 280863 3710
rect 428549 3770 428615 3773
rect 474549 3770 474615 3773
rect 428549 3768 474615 3770
rect 428549 3712 428554 3768
rect 428610 3712 474554 3768
rect 474610 3712 474615 3768
rect 428549 3710 474615 3712
rect 428549 3707 428615 3710
rect 474549 3707 474615 3710
rect 180241 3634 180307 3637
rect 281165 3634 281231 3637
rect 180241 3632 281231 3634
rect 180241 3576 180246 3632
rect 180302 3576 281170 3632
rect 281226 3576 281231 3632
rect 180241 3574 281231 3576
rect 180241 3571 180307 3574
rect 281165 3571 281231 3574
rect 410517 3634 410583 3637
rect 456885 3634 456951 3637
rect 410517 3632 456951 3634
rect 410517 3576 410522 3632
rect 410578 3576 456890 3632
rect 456946 3576 456951 3632
rect 410517 3574 456951 3576
rect 410517 3571 410583 3574
rect 456885 3571 456951 3574
rect 6453 3496 6930 3498
rect 6453 3440 6458 3496
rect 6514 3440 6930 3496
rect 6453 3438 6930 3440
rect 9949 3498 10015 3501
rect 11697 3498 11763 3501
rect 9949 3496 11763 3498
rect 9949 3440 9954 3496
rect 10010 3440 11702 3496
rect 11758 3440 11763 3496
rect 9949 3438 11763 3440
rect 6453 3435 6519 3438
rect 9949 3435 10015 3438
rect 11697 3435 11763 3438
rect 27705 3498 27771 3501
rect 35249 3498 35315 3501
rect 27705 3496 35315 3498
rect 27705 3440 27710 3496
rect 27766 3440 35254 3496
rect 35310 3440 35315 3496
rect 27705 3438 35315 3440
rect 27705 3435 27771 3438
rect 35249 3435 35315 3438
rect 64321 3498 64387 3501
rect 101397 3498 101463 3501
rect 64321 3496 101463 3498
rect 64321 3440 64326 3496
rect 64382 3440 101402 3496
rect 101458 3440 101463 3496
rect 64321 3438 101463 3440
rect 64321 3435 64387 3438
rect 101397 3435 101463 3438
rect 109309 3498 109375 3501
rect 163497 3498 163563 3501
rect 109309 3496 163563 3498
rect 109309 3440 109314 3496
rect 109370 3440 163502 3496
rect 163558 3440 163563 3496
rect 109309 3438 163563 3440
rect 109309 3435 109375 3438
rect 163497 3435 163563 3438
rect 173157 3498 173223 3501
rect 277853 3498 277919 3501
rect 173157 3496 277919 3498
rect 173157 3440 173162 3496
rect 173218 3440 277858 3496
rect 277914 3440 277919 3496
rect 173157 3438 277919 3440
rect 173157 3435 173223 3438
rect 277853 3435 277919 3438
rect 278037 3498 278103 3501
rect 279509 3498 279575 3501
rect 278037 3496 279575 3498
rect 278037 3440 278042 3496
rect 278098 3440 279514 3496
rect 279570 3440 279575 3496
rect 278037 3438 279575 3440
rect 278037 3435 278103 3438
rect 279509 3435 279575 3438
rect 282177 3498 282243 3501
rect 293677 3498 293743 3501
rect 282177 3496 293743 3498
rect 282177 3440 282182 3496
rect 282238 3440 293682 3496
rect 293738 3440 293743 3496
rect 282177 3438 293743 3440
rect 282177 3435 282243 3438
rect 293677 3435 293743 3438
rect 417417 3498 417483 3501
rect 463969 3498 464035 3501
rect 417417 3496 464035 3498
rect 417417 3440 417422 3496
rect 417478 3440 463974 3496
rect 464030 3440 464035 3496
rect 417417 3438 464035 3440
rect 417417 3435 417483 3438
rect 463969 3435 464035 3438
rect 512637 3498 512703 3501
rect 513557 3498 513623 3501
rect 512637 3496 513623 3498
rect 512637 3440 512642 3496
rect 512698 3440 513562 3496
rect 513618 3440 513623 3496
rect 512637 3438 513623 3440
rect 512637 3435 512703 3438
rect 513557 3435 513623 3438
rect 562317 3498 562383 3501
rect 563237 3498 563303 3501
rect 562317 3496 563303 3498
rect 562317 3440 562322 3496
rect 562378 3440 563242 3496
rect 563298 3440 563303 3496
rect 562317 3438 563303 3440
rect 562317 3435 562383 3438
rect 563237 3435 563303 3438
rect 5257 3362 5323 3365
rect 117957 3362 118023 3365
rect 5257 3360 118023 3362
rect 5257 3304 5262 3360
rect 5318 3304 117962 3360
rect 118018 3304 118023 3360
rect 5257 3302 118023 3304
rect 5257 3299 5323 3302
rect 117957 3299 118023 3302
rect 169569 3362 169635 3365
rect 288433 3362 288499 3365
rect 169569 3360 288499 3362
rect 169569 3304 169574 3360
rect 169630 3304 288438 3360
rect 288494 3304 288499 3360
rect 169569 3302 288499 3304
rect 169569 3299 169635 3302
rect 288433 3299 288499 3302
rect 289077 3362 289143 3365
rect 300761 3362 300827 3365
rect 289077 3360 300827 3362
rect 289077 3304 289082 3360
rect 289138 3304 300766 3360
rect 300822 3304 300827 3360
rect 289077 3302 300827 3304
rect 289077 3299 289143 3302
rect 300761 3299 300827 3302
rect 439497 3362 439563 3365
rect 582189 3362 582255 3365
rect 439497 3360 582255 3362
rect 439497 3304 439502 3360
rect 439558 3304 582194 3360
rect 582250 3304 582255 3360
rect 439497 3302 582255 3304
rect 439497 3299 439563 3302
rect 582189 3299 582255 3302
rect 240501 3226 240567 3229
rect 246297 3226 246363 3229
rect 240501 3224 246363 3226
rect 240501 3168 240506 3224
rect 240562 3168 246302 3224
rect 246358 3168 246363 3224
rect 240501 3166 246363 3168
rect 240501 3163 240567 3166
rect 246297 3163 246363 3166
rect 258257 3226 258323 3229
rect 266997 3226 267063 3229
rect 258257 3224 267063 3226
rect 258257 3168 258262 3224
rect 258318 3168 267002 3224
rect 267058 3168 267063 3224
rect 258257 3166 267063 3168
rect 258257 3163 258323 3166
rect 266997 3163 267063 3166
rect 271137 3226 271203 3229
rect 272425 3226 272491 3229
rect 271137 3224 272491 3226
rect 271137 3168 271142 3224
rect 271198 3168 272430 3224
rect 272486 3168 272491 3224
rect 271137 3166 272491 3168
rect 271137 3163 271203 3166
rect 272425 3163 272491 3166
rect 273897 3226 273963 3229
rect 276013 3226 276079 3229
rect 273897 3224 276079 3226
rect 273897 3168 273902 3224
rect 273958 3168 276018 3224
rect 276074 3168 276079 3224
rect 273897 3166 276079 3168
rect 273897 3163 273963 3166
rect 276013 3163 276079 3166
rect 432597 3226 432663 3229
rect 478137 3226 478203 3229
rect 432597 3224 478203 3226
rect 432597 3168 432602 3224
rect 432658 3168 478142 3224
rect 478198 3168 478203 3224
rect 432597 3166 478203 3168
rect 432597 3163 432663 3166
rect 478137 3163 478203 3166
rect 265341 3090 265407 3093
rect 275277 3090 275343 3093
rect 265341 3088 275343 3090
rect 265341 3032 265346 3088
rect 265402 3032 275282 3088
rect 275338 3032 275343 3088
rect 265341 3030 275343 3032
rect 265341 3027 265407 3030
rect 275277 3027 275343 3030
rect 414657 3090 414723 3093
rect 460381 3090 460447 3093
rect 414657 3088 460447 3090
rect 414657 3032 414662 3088
rect 414718 3032 460386 3088
rect 460442 3032 460447 3088
rect 414657 3030 460447 3032
rect 414657 3027 414723 3030
rect 460381 3027 460447 3030
rect 117589 2954 117655 2957
rect 264973 2954 265039 2957
rect 117589 2952 265039 2954
rect 117589 2896 117594 2952
rect 117650 2896 264978 2952
rect 265034 2896 265039 2952
rect 117589 2894 265039 2896
rect 117589 2891 117655 2894
rect 264973 2891 265039 2894
rect 53741 2818 53807 2821
rect 241421 2818 241487 2821
rect 53741 2816 241487 2818
rect 53741 2760 53746 2816
rect 53802 2760 241426 2816
rect 241482 2760 241487 2816
rect 53741 2758 241487 2760
rect 53741 2755 53807 2758
rect 241421 2755 241487 2758
<< via3 >>
rect 483060 700436 483124 700500
rect 55996 700300 56060 700364
rect 479564 700300 479628 700364
rect 59124 699756 59188 699820
rect 555372 683844 555436 683908
rect 31708 671196 31772 671260
rect 14412 658140 14476 658204
rect 55076 657596 55140 657660
rect 170996 657460 171060 657524
rect 489868 654196 489932 654260
rect 44772 644948 44836 645012
rect 52316 644676 52380 644740
rect 296484 644676 296548 644740
rect 46796 644540 46860 644604
rect 44036 644268 44100 644332
rect 375420 644268 375484 644332
rect 179276 643240 179340 643244
rect 179276 643184 179326 643240
rect 179326 643184 179340 643240
rect 179276 643180 179340 643184
rect 54708 642500 54772 642564
rect 48636 642228 48700 642292
rect 296852 642228 296916 642292
rect 177252 641684 177316 641748
rect 179092 641684 179156 641748
rect 489500 641684 489564 641748
rect 487660 641140 487724 641204
rect 50844 641004 50908 641068
rect 55812 640324 55876 640388
rect 41276 640052 41340 640116
rect 58940 639780 59004 639844
rect 486188 638964 486252 639028
rect 39804 638692 39868 638756
rect 487108 637664 487172 637668
rect 487108 637608 487158 637664
rect 487158 637608 487172 637664
rect 487108 637604 487172 637608
rect 489316 637604 489380 637668
rect 58756 637468 58820 637532
rect 485820 637060 485884 637124
rect 58572 636788 58636 636852
rect 178908 636924 178972 636988
rect 282868 636924 282932 636988
rect 52132 636516 52196 636580
rect 177620 636380 177684 636444
rect 479380 636380 479444 636444
rect 541020 636244 541084 636308
rect 48452 635564 48516 635628
rect 44956 635156 45020 635220
rect 177804 635020 177868 635084
rect 48084 634748 48148 634812
rect 296484 634748 296548 634812
rect 296668 634748 296732 634812
rect 484348 634612 484412 634676
rect 121868 634340 121932 634404
rect 121868 633796 121932 633860
rect 543780 633524 543844 633588
rect 177436 633388 177500 633452
rect 486004 633388 486068 633452
rect 179092 632164 179156 632228
rect 545068 632164 545132 632228
rect 55628 632088 55692 632092
rect 55628 632032 55642 632088
rect 55642 632032 55692 632088
rect 55628 632028 55692 632032
rect 57836 632028 57900 632092
rect 57652 630940 57716 631004
rect 551140 630804 551204 630868
rect 179276 629988 179340 630052
rect 539548 629444 539612 629508
rect 178908 628900 178972 628964
rect 59676 627744 59740 627808
rect 59860 626656 59924 626720
rect 539732 626724 539796 626788
rect 288388 625908 288452 625972
rect 286180 625092 286244 625156
rect 177804 624548 177868 624612
rect 283420 624276 283484 624340
rect 539916 624004 539980 624068
rect 177436 623460 177500 623524
rect 282132 623460 282196 623524
rect 296852 623460 296916 623524
rect 285628 622644 285692 622708
rect 177804 622372 177868 622436
rect 288572 621828 288636 621892
rect 296484 621692 296548 621756
rect 177252 621284 177316 621348
rect 285812 621012 285876 621076
rect 164004 620196 164068 620260
rect 298140 620060 298204 620124
rect 541204 619924 541268 619988
rect 291148 619380 291212 619444
rect 29132 619108 29196 619172
rect 177620 619108 177684 619172
rect 291332 618564 291396 618628
rect 543964 618564 544028 618628
rect 177436 618020 177500 618084
rect 545252 617204 545316 617268
rect 273852 617068 273916 617132
rect 177620 616932 177684 616996
rect 292804 616932 292868 616996
rect 292620 616116 292684 616180
rect 177068 615844 177132 615908
rect 173940 615300 174004 615364
rect 294460 615300 294524 615364
rect 166764 614756 166828 614820
rect 294828 614484 294892 614548
rect 177988 613668 178052 613732
rect 298508 613804 298572 613868
rect 178172 613532 178236 613596
rect 271092 613532 271156 613596
rect 293172 612852 293236 612916
rect 177804 612716 177868 612780
rect 292804 612716 292868 612780
rect 177804 612580 177868 612644
rect 175780 612036 175844 612100
rect 295564 612036 295628 612100
rect 177620 611628 177684 611692
rect 177252 611492 177316 611556
rect 286364 611492 286428 611556
rect 177436 611356 177500 611420
rect 170260 611220 170324 611284
rect 295380 611220 295444 611284
rect 177068 610676 177132 610740
rect 177620 610404 177684 610468
rect 543228 610404 543292 610468
rect 298324 610268 298388 610332
rect 177988 609724 178052 609788
rect 299612 609588 299676 609652
rect 177804 609316 177868 609380
rect 296852 609316 296916 609380
rect 542860 609044 542924 609108
rect 299244 608772 299308 608836
rect 375420 608772 375484 608836
rect 298140 608500 298204 608564
rect 165476 608228 165540 608292
rect 298692 607956 298756 608020
rect 539364 607684 539428 607748
rect 176884 607140 176948 607204
rect 294644 607140 294708 607204
rect 177252 607004 177316 607068
rect 177988 607004 178052 607068
rect 271276 607004 271340 607068
rect 272012 606324 272076 606388
rect 542676 606324 542740 606388
rect 11652 606052 11716 606116
rect 177436 605780 177500 605844
rect 299060 605508 299124 605572
rect 177068 604964 177132 605028
rect 296668 604964 296732 605028
rect 175964 604692 176028 604756
rect 269804 604692 269868 604756
rect 177620 604420 177684 604484
rect 298508 604420 298572 604484
rect 173756 603876 173820 603940
rect 262812 603876 262876 603940
rect 280660 603876 280724 603940
rect 540100 603604 540164 603668
rect 265940 603060 266004 603124
rect 177620 602788 177684 602852
rect 255820 602788 255884 602852
rect 280844 602244 280908 602308
rect 377628 602244 377692 602308
rect 177804 601700 177868 601764
rect 538260 601836 538324 601900
rect 538444 601700 538508 601764
rect 266860 601428 266924 601492
rect 543044 601080 543108 601084
rect 543044 601024 543094 601080
rect 543094 601024 543108 601080
rect 543044 601020 543108 601024
rect 277900 600612 277964 600676
rect 537340 600476 537404 600540
rect 542676 600476 542740 600540
rect 534580 600068 534644 600132
rect 542676 600204 542740 600268
rect 526300 599932 526364 599996
rect 540100 599932 540164 599996
rect 256740 599796 256804 599860
rect 522252 599660 522316 599724
rect 543964 599660 544028 599724
rect 522436 599524 522500 599588
rect 545068 599524 545132 599588
rect 537524 599388 537588 599452
rect 545252 599388 545316 599452
rect 533292 599116 533356 599180
rect 295748 598980 295812 599044
rect 536052 598300 536116 598364
rect 275140 598164 275204 598228
rect 490420 598164 490484 598228
rect 492996 598164 493060 598228
rect 494100 598164 494164 598228
rect 496860 598164 496924 598228
rect 530532 598164 530596 598228
rect 294828 597484 294892 597548
rect 295012 597212 295076 597276
rect 501460 596804 501524 596868
rect 256924 596532 256988 596596
rect 257108 595716 257172 595780
rect 508452 595444 508516 595508
rect 542860 595444 542924 595508
rect 268148 594900 268212 594964
rect 256740 594764 256804 594828
rect 543596 594764 543660 594828
rect 269620 594084 269684 594148
rect 506980 593948 507044 594012
rect 543228 593948 543292 594012
rect 543412 593464 543476 593468
rect 543412 593408 543426 593464
rect 543426 593408 543476 593464
rect 543412 593404 543476 593408
rect 296300 593268 296364 593332
rect 518020 592588 518084 592652
rect 543044 592588 543108 592652
rect 294828 592452 294892 592516
rect 294460 592044 294524 592108
rect 298876 591636 298940 591700
rect 298324 591364 298388 591428
rect 265756 590820 265820 590884
rect 295564 590548 295628 590612
rect 296116 590004 296180 590068
rect 268332 589188 268396 589252
rect 277164 588372 277228 588436
rect 284892 587556 284956 587620
rect 291516 586740 291580 586804
rect 295932 585924 295996 585988
rect 289124 585108 289188 585172
rect 295380 585108 295444 585172
rect 286548 584292 286612 584356
rect 285812 583748 285876 583812
rect 283604 583476 283668 583540
rect 271460 582660 271524 582724
rect 290596 581844 290660 581908
rect 274036 581028 274100 581092
rect 292252 580212 292316 580276
rect 291332 579532 291396 579596
rect 290964 579396 291028 579460
rect 291884 578580 291948 578644
rect 290596 578172 290660 578236
rect 291148 578172 291212 578236
rect 291700 577628 291764 577692
rect 548380 577628 548444 577692
rect 290780 576948 290844 577012
rect 381308 576948 381372 577012
rect 295564 576132 295628 576196
rect 295748 575452 295812 575516
rect 256740 575316 256804 575380
rect 292988 574364 293052 574428
rect 256924 574092 256988 574156
rect 292620 574092 292684 574156
rect 292068 573684 292132 573748
rect 291516 572868 291580 572932
rect 292436 572868 292500 572932
rect 292252 572792 292316 572796
rect 292252 572736 292266 572792
rect 292266 572736 292316 572792
rect 292252 572732 292316 572736
rect 54892 572324 54956 572388
rect 294460 572052 294524 572116
rect 383700 572052 383764 572116
rect 294644 571372 294708 571436
rect 169524 571100 169588 571164
rect 379468 571236 379532 571300
rect 299796 571100 299860 571164
rect 299428 570420 299492 570484
rect 382228 570420 382292 570484
rect 171548 570148 171612 570212
rect 281028 570148 281092 570212
rect 299244 570012 299308 570076
rect 299612 570012 299676 570076
rect 177252 569876 177316 569940
rect 295564 569604 295628 569668
rect 177804 569060 177868 569124
rect 288940 568788 289004 568852
rect 379652 568788 379716 568852
rect 296300 568652 296364 568716
rect 173572 567972 173636 568036
rect 29500 566884 29564 566948
rect 179276 566884 179340 566948
rect 285260 566884 285324 566948
rect 174860 565796 174924 565860
rect 277164 565796 277228 565860
rect 175044 564708 175108 564772
rect 279372 564708 279436 564772
rect 60412 564640 60476 564704
rect 54524 564300 54588 564364
rect 285076 563620 285140 563684
rect 179092 563484 179156 563548
rect 295748 563212 295812 563276
rect 296484 563212 296548 563276
rect 287836 562532 287900 562596
rect 60596 562464 60660 562528
rect 180564 562464 180628 562528
rect 179276 562124 179340 562188
rect 59124 560356 59188 560420
rect 179828 561376 179892 561440
rect 276980 560764 277044 560828
rect 476620 560492 476684 560556
rect 277164 560356 277228 560420
rect 173940 560220 174004 560284
rect 177988 560220 178052 560284
rect 296484 559948 296548 560012
rect 514156 559948 514220 560012
rect 277900 559812 277964 559876
rect 498516 559812 498580 559876
rect 47900 559268 47964 559332
rect 268148 559268 268212 559332
rect 474412 559268 474476 559332
rect 47716 559132 47780 559196
rect 282684 558996 282748 559060
rect 55996 558860 56060 558924
rect 60596 558860 60660 558924
rect 60412 558724 60476 558788
rect 280844 558860 280908 558924
rect 281396 558860 281460 558924
rect 487292 558996 487356 559060
rect 180564 558316 180628 558380
rect 510844 558316 510908 558380
rect 54892 558180 54956 558244
rect 179092 558180 179156 558244
rect 511028 558180 511092 558244
rect 173756 558044 173820 558108
rect 280844 558044 280908 558108
rect 33732 557636 33796 557700
rect 281396 557772 281460 557836
rect 501276 557772 501340 557836
rect 31524 557500 31588 557564
rect 265940 557092 266004 557156
rect 478092 557092 478156 557156
rect 55444 556548 55508 556612
rect 53604 556412 53668 556476
rect 33916 556276 33980 556340
rect 177804 555324 177868 555388
rect 494284 555324 494348 555388
rect 177436 555188 177500 555252
rect 275140 555052 275204 555116
rect 502748 555052 502812 555116
rect 176884 554644 176948 554708
rect 294828 554372 294892 554436
rect 501092 554372 501156 554436
rect 290780 554236 290844 554300
rect 499804 554236 499868 554300
rect 174860 553964 174924 554028
rect 499620 553964 499684 554028
rect 2820 553828 2884 553892
rect 47532 553420 47596 553484
rect 57652 553284 57716 553348
rect 170996 553148 171060 553212
rect 173572 553148 173636 553212
rect 481772 553148 481836 553212
rect 291884 553012 291948 553076
rect 498332 553012 498396 553076
rect 262812 552876 262876 552940
rect 476068 552876 476132 552940
rect 166764 552740 166828 552804
rect 292436 552740 292500 552804
rect 510660 552740 510724 552804
rect 292068 552604 292132 552668
rect 512132 552604 512196 552668
rect 296116 552468 296180 552532
rect 476804 552468 476868 552532
rect 46612 552060 46676 552124
rect 169524 551516 169588 551580
rect 164004 550972 164068 551036
rect 269804 550972 269868 551036
rect 478276 550972 478340 551036
rect 41092 550700 41156 550764
rect 32996 550292 33060 550356
rect 271276 550292 271340 550356
rect 286548 550292 286612 550356
rect 500908 550292 500972 550356
rect 39436 549476 39500 549540
rect 31156 549340 31220 549404
rect 59124 548932 59188 548996
rect 296300 549204 296364 549268
rect 295748 549068 295812 549132
rect 505140 549068 505204 549132
rect 299060 548932 299124 548996
rect 500172 548932 500236 548996
rect 34284 548796 34348 548860
rect 273852 548796 273916 548860
rect 274036 548796 274100 548860
rect 502380 548796 502444 548860
rect 170260 547708 170324 547772
rect 57836 547572 57900 547636
rect 256740 547572 256804 547636
rect 487476 547572 487540 547636
rect 271460 547436 271524 547500
rect 502564 547436 502628 547500
rect 59676 546348 59740 546412
rect 30236 546076 30300 546140
rect 286364 546076 286428 546140
rect 292988 546076 293052 546140
rect 511212 546076 511276 546140
rect 59676 545804 59740 545868
rect 289124 545532 289188 545596
rect 498700 545532 498764 545596
rect 486372 545124 486436 545188
rect 31340 544308 31404 544372
rect 277164 544308 277228 544372
rect 295012 544308 295076 544372
rect 506612 544308 506676 544372
rect 43852 544172 43916 544236
rect 293172 543356 293236 543420
rect 481956 543356 482020 543420
rect 175964 542948 176028 543012
rect 32812 540500 32876 540564
rect 281028 540500 281092 540564
rect 272012 540092 272076 540156
rect 494468 540092 494532 540156
rect 482140 538052 482204 538116
rect 165476 537372 165540 537436
rect 32444 536828 32508 536892
rect 30052 536012 30116 536076
rect 382228 536012 382292 536076
rect 32628 535196 32692 535260
rect 276980 535196 277044 535260
rect 35756 535060 35820 535124
rect 285260 535060 285324 535124
rect 42380 534788 42444 534852
rect 379652 534788 379716 534852
rect 30972 534652 31036 534716
rect 383700 534652 383764 534716
rect 31708 534108 31772 534172
rect 379836 534108 379900 534172
rect 29132 533292 29196 533356
rect 29868 533156 29932 533220
rect 379468 533292 379532 533356
rect 283420 533156 283484 533220
rect 495388 533156 495452 533220
rect 266860 532340 266924 532404
rect 502932 532340 502996 532404
rect 286180 531796 286244 531860
rect 498148 531796 498212 531860
rect 37044 531388 37108 531452
rect 282132 531252 282196 531316
rect 288572 530436 288636 530500
rect 55628 529816 55692 529820
rect 55628 529760 55678 529816
rect 55678 529760 55692 529816
rect 55628 529756 55692 529760
rect 57836 529348 57900 529412
rect 177068 529348 177132 529412
rect 288388 529348 288452 529412
rect 55996 528940 56060 529004
rect 377628 529076 377692 529140
rect 175780 527716 175844 527780
rect 285628 527580 285692 527644
rect 36492 527172 36556 527236
rect 483244 526628 483308 526692
rect 299796 526220 299860 526284
rect 503668 526220 503732 526284
rect 171548 526084 171612 526148
rect 288940 525948 289004 526012
rect 493180 525948 493244 526012
rect 37228 525812 37292 525876
rect 175044 525676 175108 525740
rect 179828 525676 179892 525740
rect 295932 525676 295996 525740
rect 497044 525676 497108 525740
rect 294460 525540 294524 525604
rect 507900 525540 507964 525604
rect 299244 524860 299308 524924
rect 499988 524860 500052 524924
rect 547092 524452 547156 524516
rect 35204 524044 35268 524108
rect 58572 523772 58636 523836
rect 39620 523636 39684 523700
rect 280844 523636 280908 523700
rect 36676 523364 36740 523428
rect 58388 523092 58452 523156
rect 482324 523092 482388 523156
rect 55812 523016 55876 523020
rect 55812 522960 55826 523016
rect 55826 522960 55876 523016
rect 55812 522956 55876 522960
rect 59492 523016 59556 523020
rect 59492 522960 59542 523016
rect 59542 522960 59556 523016
rect 59492 522956 59556 522960
rect 257108 522820 257172 522884
rect 480300 522820 480364 522884
rect 43668 522548 43732 522612
rect 59860 522548 59924 522612
rect 55996 522412 56060 522476
rect 296852 522412 296916 522476
rect 298692 522412 298756 522476
rect 495572 522412 495636 522476
rect 34100 522276 34164 522340
rect 280660 522276 280724 522340
rect 35388 522140 35452 522204
rect 39252 521732 39316 521796
rect 58940 521596 59004 521660
rect 59308 521052 59372 521116
rect 279372 521052 279436 521116
rect 36860 520916 36924 520980
rect 287836 520916 287900 520980
rect 50476 520644 50540 520708
rect 42564 520236 42628 520300
rect 495388 520100 495452 520164
rect 283604 519964 283668 520028
rect 490052 519964 490116 520028
rect 35572 519828 35636 519892
rect 37412 519556 37476 519620
rect 54892 519556 54956 519620
rect 57652 519556 57716 519620
rect 255820 519556 255884 519620
rect 265756 519556 265820 519620
rect 490236 519556 490300 519620
rect 285076 519420 285140 519484
rect 290964 519420 291028 519484
rect 50292 519284 50356 519348
rect 291700 519284 291764 519348
rect 491340 519284 491404 519348
rect 46428 519148 46492 519212
rect 284892 519148 284956 519212
rect 494652 519148 494716 519212
rect 43484 519012 43548 519076
rect 483428 519012 483492 519076
rect 54524 518876 54588 518940
rect 269620 518876 269684 518940
rect 495204 518876 495268 518940
rect 476068 518740 476132 518804
rect 478092 518740 478156 518804
rect 58572 518604 58636 518668
rect 271092 518604 271156 518668
rect 298876 518604 298940 518668
rect 497228 518604 497292 518668
rect 268332 518468 268396 518532
rect 503852 518468 503916 518532
rect 50660 518332 50724 518396
rect 379836 518332 379900 518396
rect 476804 518332 476868 518396
rect 44588 518196 44652 518260
rect 381308 518196 381372 518260
rect 491524 518196 491588 518260
rect 474412 518060 474476 518124
rect 478276 518060 478340 518124
rect 54524 517924 54588 517988
rect 476620 517924 476684 517988
rect 493364 518060 493428 518124
rect 58756 517516 58820 517580
rect 481772 517244 481836 517308
rect 481772 516836 481836 516900
rect 482324 516700 482388 516764
rect 482140 515884 482204 515948
rect 57836 514932 57900 514996
rect 3004 514796 3068 514860
rect 481956 512348 482020 512412
rect 483060 511940 483124 512004
rect 44772 510580 44836 510644
rect 43300 510444 43364 510508
rect 39804 510036 39868 510100
rect 44036 509492 44100 509556
rect 495572 508948 495636 509012
rect 490420 508540 490484 508604
rect 41276 508404 41340 508468
rect 50292 507860 50356 507924
rect 494468 507860 494532 507924
rect 500172 507316 500236 507380
rect 54524 506772 54588 506836
rect 43668 505684 43732 505748
rect 44036 505200 44100 505204
rect 44036 505144 44050 505200
rect 44050 505144 44100 505200
rect 44036 505140 44100 505144
rect 55628 505140 55692 505204
rect 501276 505140 501340 505204
rect 50476 505004 50540 505068
rect 57468 505004 57532 505068
rect 59492 504596 59556 504660
rect 502932 504596 502996 504660
rect 35204 504052 35268 504116
rect 498516 504052 498580 504116
rect 58756 502420 58820 502484
rect 502748 502420 502812 502484
rect 59124 502288 59188 502352
rect 4660 501740 4724 501804
rect 506612 501876 506676 501940
rect 36492 501332 36556 501396
rect 35388 500788 35452 500852
rect 480300 500652 480364 500716
rect 46428 499020 46492 499084
rect 57468 499020 57532 499084
rect 57284 498612 57348 498676
rect 501092 498612 501156 498676
rect 46244 498204 46308 498268
rect 497228 498068 497292 498132
rect 490236 497524 490300 497588
rect 491524 496980 491588 497044
rect 50660 496708 50724 496772
rect 57284 496708 57348 496772
rect 503852 496436 503916 496500
rect 57468 495892 57532 495956
rect 493364 495892 493428 495956
rect 487660 495484 487724 495548
rect 494652 495348 494716 495412
rect 33732 494804 33796 494868
rect 497044 494260 497108 494324
rect 498700 493716 498764 493780
rect 500908 493172 500972 493236
rect 52132 492628 52196 492692
rect 490052 492628 490116 492692
rect 36676 492084 36740 492148
rect 502564 492084 502628 492148
rect 42564 491132 42628 491196
rect 43484 490996 43548 491060
rect 502380 490996 502444 491060
rect 42748 490452 42812 490516
rect 41092 490044 41156 490108
rect 495388 489908 495452 489972
rect 39252 489364 39316 489428
rect 498332 489364 498396 489428
rect 57284 488820 57348 488884
rect 491340 488820 491404 488884
rect 44588 488276 44652 488340
rect 499804 488276 499868 488340
rect 55444 487732 55508 487796
rect 514156 487732 514220 487796
rect 487476 487324 487540 487388
rect 511396 486644 511460 486708
rect 33916 486100 33980 486164
rect 512132 486100 512196 486164
rect 511212 485828 511276 485892
rect 39436 485556 39500 485620
rect 510660 485556 510724 485620
rect 30972 485012 31036 485076
rect 507900 485012 507964 485076
rect 29868 484468 29932 484532
rect 580212 484604 580276 484668
rect 503668 484468 503732 484532
rect 30052 483924 30116 483988
rect 499988 483924 500052 483988
rect 32444 483380 32508 483444
rect 505140 483380 505204 483444
rect 42380 482972 42444 483036
rect 42380 482836 42444 482900
rect 493180 482836 493244 482900
rect 54708 476852 54772 476916
rect 544332 471412 544396 471476
rect 486188 465836 486252 465900
rect 3372 462572 3436 462636
rect 487108 460124 487172 460188
rect 489500 459036 489564 459100
rect 46244 457812 46308 457876
rect 46796 457268 46860 457332
rect 46428 456860 46492 456924
rect 50844 456180 50908 456244
rect 484348 456316 484412 456380
rect 485820 455772 485884 455836
rect 48452 455092 48516 455156
rect 59676 454548 59740 454612
rect 48636 454004 48700 454068
rect 486004 454004 486068 454068
rect 52316 453460 52380 453524
rect 48084 452916 48148 452980
rect 47532 452372 47596 452436
rect 47716 451828 47780 451892
rect 479380 451828 479444 451892
rect 58388 451284 58452 451348
rect 34284 450740 34348 450804
rect 483428 450604 483492 450668
rect 39620 450196 39684 450260
rect 487292 450060 487356 450124
rect 37228 449652 37292 449716
rect 3556 449516 3620 449580
rect 58572 449108 58636 449172
rect 31524 448564 31588 448628
rect 30236 448020 30300 448084
rect 31156 447476 31220 447540
rect 55996 446932 56060 446996
rect 47900 446388 47964 446452
rect 32996 445844 33060 445908
rect 46612 445300 46676 445364
rect 59124 444756 59188 444820
rect 34100 444212 34164 444276
rect 57652 443668 57716 443732
rect 32628 443124 32692 443188
rect 499620 443124 499684 443188
rect 58940 442580 59004 442644
rect 37412 442036 37476 442100
rect 511028 442036 511092 442100
rect 36860 441492 36924 441556
rect 510844 441492 510908 441556
rect 35572 440948 35636 441012
rect 31340 440404 31404 440468
rect 32812 439860 32876 439924
rect 53604 439316 53668 439380
rect 494284 439316 494348 439380
rect 37044 438772 37108 438836
rect 35756 438228 35820 438292
rect 483244 420684 483308 420748
rect 483612 420140 483676 420204
rect 543412 420140 543476 420204
rect 558132 418236 558196 418300
rect 42380 416468 42444 416532
rect 44036 415924 44100 415988
rect 498148 415924 498212 415988
rect 43300 415380 43364 415444
rect 43852 414836 43916 414900
rect 44956 414292 45020 414356
rect 46428 413748 46492 413812
rect 42564 413204 42628 413268
rect 3740 410484 3804 410548
rect 3004 409940 3068 410004
rect 481772 403004 481836 403068
rect 486372 400012 486436 400076
rect 2820 398108 2884 398172
rect 3924 397428 3988 397492
rect 489316 394844 489380 394908
rect 479564 388724 479628 388788
rect 55076 387500 55140 387564
rect 3556 384236 3620 384300
rect 210372 384236 210436 384300
rect 239812 384236 239876 384300
rect 239628 382740 239692 382804
rect 3924 381516 3988 381580
rect 206140 381516 206204 381580
rect 282132 381516 282196 381580
rect 541204 381516 541268 381580
rect 541388 380972 541452 381036
rect 281764 379476 281828 379540
rect 236132 378388 236196 378452
rect 3740 377980 3804 378044
rect 284340 377980 284404 378044
rect 281948 376756 282012 376820
rect 492996 374716 493060 374780
rect 235764 373220 235828 373284
rect 3372 370500 3436 370564
rect 282868 370500 282932 370564
rect 580396 365060 580460 365124
rect 294460 358396 294524 358460
rect 239444 355404 239508 355468
rect 496860 349964 496924 350028
rect 238524 349828 238588 349892
rect 237236 349692 237300 349756
rect 580212 349692 580276 349756
rect 238340 348332 238404 348396
rect 239260 347108 239324 347172
rect 238156 345748 238220 345812
rect 494100 345748 494164 345812
rect 230980 345340 231044 345404
rect 48084 344524 48148 344588
rect 231164 344388 231228 344452
rect 224356 344116 224420 344180
rect 230060 343980 230124 344044
rect 229876 343844 229940 343908
rect 285996 343844 286060 343908
rect 227484 343572 227548 343636
rect 224908 343436 224972 343500
rect 227116 343028 227180 343092
rect 223252 342620 223316 342684
rect 224540 342484 224604 342548
rect 227300 342348 227364 342412
rect 224172 342212 224236 342276
rect 29500 342076 29564 342140
rect 222884 341940 222948 342004
rect 285628 341940 285692 342004
rect 226196 341804 226260 341868
rect 284524 341804 284588 341868
rect 223068 341260 223132 341324
rect 251036 341260 251100 341324
rect 251036 340444 251100 340508
rect 285812 340444 285876 340508
rect 226932 339900 226996 339964
rect 222700 339492 222764 339556
rect 287100 339492 287164 339556
rect 280660 338812 280724 338876
rect 490052 338676 490116 338740
rect 228220 338268 228284 338332
rect 284708 338268 284772 338332
rect 228404 338132 228468 338196
rect 290596 338132 290660 338196
rect 233740 337588 233804 337652
rect 281580 337588 281644 337652
rect 295932 337316 295996 337380
rect 580396 337316 580460 337380
rect 238524 336228 238588 336292
rect 287652 335956 287716 336020
rect 542676 335956 542740 336020
rect 239260 335140 239324 335204
rect 238340 333916 238404 333980
rect 298692 333236 298756 333300
rect 543596 333236 543660 333300
rect 536052 328748 536116 328812
rect 538444 327932 538508 327996
rect 530532 327116 530596 327180
rect 533292 326300 533356 326364
rect 501460 325484 501524 325548
rect 538260 324668 538324 324732
rect 511212 323852 511276 323916
rect 541388 320588 541452 320652
rect 541020 319772 541084 319836
rect 543780 318140 543844 318204
rect 522436 317324 522500 317388
rect 539548 315692 539612 315756
rect 539732 314060 539796 314124
rect 539916 312428 539980 312492
rect 580212 312020 580276 312084
rect 281764 311612 281828 311676
rect 282316 311068 282380 311132
rect 539364 311068 539428 311132
rect 281948 310796 282012 310860
rect 282132 309980 282196 310044
rect 522252 309164 522316 309228
rect 537524 308348 537588 308412
rect 483612 307532 483676 307596
rect 298692 306716 298756 306780
rect 228404 306172 228468 306236
rect 287652 305900 287716 305964
rect 518020 305084 518084 305148
rect 506980 304268 507044 304332
rect 508452 303452 508516 303516
rect 282316 302636 282380 302700
rect 238156 302500 238220 302564
rect 537340 301820 537404 301884
rect 534580 301004 534644 301068
rect 526300 300188 526364 300252
rect 239444 298012 239508 298076
rect 239628 293728 239692 293792
rect 122052 293116 122116 293180
rect 280660 291212 280724 291276
rect 235948 289716 236012 289780
rect 236132 289580 236196 289644
rect 237972 289580 238036 289644
rect 11652 286316 11716 286380
rect 238156 286316 238220 286380
rect 345612 276660 345676 276724
rect 580212 276660 580276 276724
rect 14412 273804 14476 273868
rect 237420 273804 237484 273868
rect 4660 272444 4724 272508
rect 238524 272444 238588 272508
rect 284524 265916 284588 265980
rect 285996 264284 286060 264348
rect 284708 263468 284772 263532
rect 281580 261020 281644 261084
rect 54892 260068 54956 260132
rect 285812 259252 285876 259316
rect 287652 258844 287716 258908
rect 227484 258572 227548 258636
rect 285628 258708 285692 258772
rect 226748 257756 226812 257820
rect 287100 257892 287164 257956
rect 227300 256940 227364 257004
rect 226564 256668 226628 256732
rect 224908 255308 224972 255372
rect 48636 254084 48700 254148
rect 227116 253676 227180 253740
rect 287100 253812 287164 253876
rect 226196 252044 226260 252108
rect 292620 252044 292684 252108
rect 230060 250412 230124 250476
rect 229876 248780 229940 248844
rect 285812 248644 285876 248708
rect 228220 247148 228284 247212
rect 288388 246196 288452 246260
rect 231164 245516 231228 245580
rect 291332 245380 291396 245444
rect 48084 244972 48148 245036
rect 291148 244564 291212 244628
rect 224540 243884 224604 243948
rect 291516 243884 291580 243948
rect 233740 242252 233804 242316
rect 288572 242252 288636 242316
rect 290780 241436 290844 241500
rect 3372 241028 3436 241092
rect 223252 240620 223316 240684
rect 223068 238988 223132 239052
rect 222884 237356 222948 237420
rect 222700 235724 222764 235788
rect 226932 234092 226996 234156
rect 224356 232460 224420 232524
rect 226564 230828 226628 230892
rect 226380 229196 226444 229260
rect 232268 227564 232332 227628
rect 224172 225932 224236 225996
rect 232084 224300 232148 224364
rect 580212 218996 580276 219060
rect 239812 218656 239876 218720
rect 238340 217772 238404 217836
rect 224172 217636 224236 217700
rect 237420 216684 237484 216748
rect 219940 216548 220004 216612
rect 228220 215460 228284 215524
rect 231164 213284 231228 213348
rect 235212 212876 235276 212940
rect 116532 212196 116596 212260
rect 235396 211244 235460 211308
rect 280844 211244 280908 211308
rect 122052 210972 122116 211036
rect 281764 210428 281828 210492
rect 230980 210020 231044 210084
rect 235580 209612 235644 209676
rect 206140 208932 206204 208996
rect 281948 208796 282012 208860
rect 235028 207980 235092 208044
rect 210372 207844 210436 207908
rect 235764 207028 235828 207092
rect 238524 206756 238588 206820
rect 239260 204716 239324 204780
rect 238156 204580 238220 204644
rect 238156 203084 238220 203148
rect 48452 201860 48516 201924
rect 3372 199140 3436 199204
rect 116532 199140 116596 199204
rect 285628 195740 285692 195804
rect 342852 195196 342916 195260
rect 580212 195196 580276 195260
rect 280660 194924 280724 194988
rect 284524 192476 284588 192540
rect 235948 189348 236012 189412
rect 281580 189212 281644 189276
rect 231164 188804 231228 188868
rect 237236 188260 237300 188324
rect 237972 186084 238036 186148
rect 284708 185132 284772 185196
rect 283420 184316 283484 184380
rect 279372 183500 279436 183564
rect 237788 182684 237852 182748
rect 281028 182684 281092 182748
rect 282132 181868 282196 181932
rect 237972 181596 238036 181660
rect 239628 180576 239692 180640
rect 283052 180236 283116 180300
rect 239812 179488 239876 179552
rect 283236 179420 283300 179484
rect 288940 179148 289004 179212
rect 288756 177788 288820 177852
rect 290596 176156 290660 176220
rect 294460 175340 294524 175404
rect 284340 174524 284404 174588
rect 282868 173708 282932 173772
rect 555372 162284 555436 162348
rect 551140 161468 551204 161532
rect 548380 160652 548444 160716
rect 547092 159836 547156 159900
rect 544332 159020 544396 159084
rect 558132 158204 558196 158268
rect 295932 157388 295996 157452
rect 345612 156572 345676 156636
rect 287652 155756 287716 155820
rect 342852 154940 342916 155004
rect 288940 154124 289004 154188
rect 351132 153308 351196 153372
rect 306972 152492 307036 152556
rect 288940 151676 289004 151740
rect 551140 150860 551204 150924
rect 3372 149772 3436 149836
rect 240364 144672 240428 144736
rect 240180 142496 240244 142560
rect 232084 142020 232148 142084
rect 292620 142020 292684 142084
rect 238340 141476 238404 141540
rect 285812 141476 285876 141540
rect 240180 141340 240244 141404
rect 273300 141340 273364 141404
rect 48636 140660 48700 140724
rect 237788 140720 237852 140724
rect 237788 140664 237802 140720
rect 237802 140664 237852 140720
rect 237788 140660 237852 140664
rect 237972 140660 238036 140724
rect 239628 140720 239692 140724
rect 239628 140664 239678 140720
rect 239678 140664 239692 140720
rect 239628 140660 239692 140664
rect 3372 140524 3436 140588
rect 48452 140388 48516 140452
rect 288756 140388 288820 140452
rect 273300 139708 273364 139772
rect 240916 139572 240980 139636
rect 288756 139436 288820 139500
rect 351132 139300 351196 139364
rect 235028 139164 235092 139228
rect 235764 139028 235828 139092
rect 291516 139028 291580 139092
rect 291332 138892 291396 138956
rect 235948 138756 236012 138820
rect 291148 138756 291212 138820
rect 239260 138484 239324 138548
rect 288572 138484 288636 138548
rect 3372 138076 3436 138140
rect 235396 138076 235460 138140
rect 288388 138212 288452 138276
rect 232268 137804 232332 137868
rect 287100 137804 287164 137868
rect 238156 137668 238220 137732
rect 290780 137668 290844 137732
rect 3372 136716 3436 136780
rect 284708 134404 284772 134468
rect 3372 133044 3436 133108
rect 283236 133044 283300 133108
rect 280844 130460 280908 130524
rect 281948 127740 282012 127804
rect 281028 127604 281092 127668
rect 282132 126244 282196 126308
rect 281764 118084 281828 118148
rect 279372 116452 279436 116516
rect 283420 115092 283484 115156
rect 239812 112780 239876 112844
rect 306972 99452 307036 99516
rect 3372 97548 3436 97612
rect 281580 97140 281644 97204
rect 3740 88980 3804 89044
rect 283052 88980 283116 89044
rect 288940 88980 289004 89044
rect 580212 88980 580276 89044
rect 3372 86260 3436 86324
rect 228220 86260 228284 86324
rect 3372 84628 3436 84692
rect 580212 59604 580276 59668
rect 3372 58516 3436 58580
rect 280660 49268 280724 49332
rect 490420 46276 490484 46340
rect 219940 45460 220004 45524
rect 284524 44916 284588 44980
rect 285628 37980 285692 38044
rect 551140 19756 551204 19820
rect 288756 19348 288820 19412
rect 4108 7652 4172 7716
rect 224172 7652 224236 7716
rect 4108 6428 4172 6492
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 2819 553892 2885 553893
rect 2819 553828 2820 553892
rect 2884 553828 2885 553892
rect 2819 553827 2885 553828
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 2822 398173 2882 553827
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 3003 514860 3069 514861
rect 3003 514796 3004 514860
rect 3068 514796 3069 514860
rect 3003 514795 3069 514796
rect 3006 410005 3066 514795
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 4659 501804 4725 501805
rect 4659 501740 4660 501804
rect 4724 501740 4725 501804
rect 4659 501739 4725 501740
rect 3371 462636 3437 462637
rect 3371 462572 3372 462636
rect 3436 462572 3437 462636
rect 3371 462571 3437 462572
rect 3003 410004 3069 410005
rect 3003 409940 3004 410004
rect 3068 409940 3069 410004
rect 3003 409939 3069 409940
rect 2819 398172 2885 398173
rect 2819 398108 2820 398172
rect 2884 398108 2885 398172
rect 2819 398107 2885 398108
rect 3374 370565 3434 462571
rect 3555 449580 3621 449581
rect 3555 449516 3556 449580
rect 3620 449516 3621 449580
rect 3555 449515 3621 449516
rect 3558 384301 3618 449515
rect 3739 410548 3805 410549
rect 3739 410484 3740 410548
rect 3804 410484 3805 410548
rect 3739 410483 3805 410484
rect 3555 384300 3621 384301
rect 3555 384236 3556 384300
rect 3620 384236 3621 384300
rect 3555 384235 3621 384236
rect 3742 378045 3802 410483
rect 3923 397492 3989 397493
rect 3923 397428 3924 397492
rect 3988 397428 3989 397492
rect 3923 397427 3989 397428
rect 3926 381581 3986 397427
rect 3923 381580 3989 381581
rect 3923 381516 3924 381580
rect 3988 381516 3989 381580
rect 3923 381515 3989 381516
rect 3739 378044 3805 378045
rect 3739 377980 3740 378044
rect 3804 377980 3805 378044
rect 3739 377979 3805 377980
rect 3371 370564 3437 370565
rect 3371 370500 3372 370564
rect 3436 370500 3437 370564
rect 3371 370499 3437 370500
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 4662 272509 4722 501739
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 4659 272508 4725 272509
rect 4659 272444 4660 272508
rect 4724 272444 4725 272508
rect 4659 272443 4725 272444
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 3371 241092 3437 241093
rect 3371 241028 3372 241092
rect 3436 241028 3437 241092
rect 3371 241027 3437 241028
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 3374 199205 3434 241027
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 3371 199204 3437 199205
rect 3371 199140 3372 199204
rect 3436 199140 3437 199204
rect 3371 199139 3437 199140
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 3371 149836 3437 149837
rect 3371 149772 3372 149836
rect 3436 149772 3437 149836
rect 3371 149771 3437 149772
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 3374 140589 3434 149771
rect 3371 140588 3437 140589
rect 3371 140524 3372 140588
rect 3436 140524 3437 140588
rect 3371 140523 3437 140524
rect 3371 138140 3437 138141
rect 3371 138076 3372 138140
rect 3436 138076 3437 138140
rect 3371 138075 3437 138076
rect 3374 136781 3434 138075
rect 3371 136780 3437 136781
rect 3371 136716 3372 136780
rect 3436 136716 3437 136780
rect 3371 136715 3437 136716
rect 3371 133108 3437 133109
rect 3371 133044 3372 133108
rect 3436 133044 3437 133108
rect 3371 133043 3437 133044
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 3374 97613 3434 133043
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3371 97612 3437 97613
rect 3371 97548 3372 97612
rect 3436 97548 3437 97612
rect 3371 97547 3437 97548
rect 3739 89044 3805 89045
rect 3739 88980 3740 89044
rect 3804 88980 3805 89044
rect 3739 88979 3805 88980
rect 3371 86324 3437 86325
rect 3371 86260 3372 86324
rect 3436 86260 3437 86324
rect 3371 86259 3437 86260
rect 3374 84693 3434 86259
rect 3371 84692 3437 84693
rect 3371 84628 3372 84692
rect 3436 84628 3437 84692
rect 3371 84627 3437 84628
rect 3742 84210 3802 88979
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 84150 3802 84210
rect 3374 58581 3434 84150
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3371 58580 3437 58581
rect 3371 58516 3372 58580
rect 3436 58516 3437 58580
rect 3371 58515 3437 58516
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 4107 7716 4173 7717
rect 4107 7652 4108 7716
rect 4172 7652 4173 7716
rect 4107 7651 4173 7652
rect 4110 6493 4170 7651
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 4107 6492 4173 6493
rect 4107 6428 4108 6492
rect 4172 6428 4173 6492
rect 4107 6427 4173 6428
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 14411 658204 14477 658205
rect 14411 658140 14412 658204
rect 14476 658140 14477 658204
rect 14411 658139 14477 658140
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 11651 606116 11717 606117
rect 11651 606052 11652 606116
rect 11716 606052 11717 606116
rect 11651 606051 11717 606052
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 11654 286381 11714 606051
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 11651 286380 11717 286381
rect 11651 286316 11652 286380
rect 11716 286316 11717 286380
rect 11651 286315 11717 286316
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 266614 13574 302058
rect 14414 273869 14474 658139
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 14411 273868 14477 273869
rect 14411 273804 14412 273868
rect 14476 273804 14477 273868
rect 14411 273803 14477 273804
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 31707 671260 31773 671261
rect 31707 671196 31708 671260
rect 31772 671196 31773 671260
rect 31707 671195 31773 671196
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 29131 619172 29197 619173
rect 29131 619108 29132 619172
rect 29196 619108 29197 619172
rect 29131 619107 29197 619108
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 29134 533357 29194 619107
rect 29499 566948 29565 566949
rect 29499 566884 29500 566948
rect 29564 566884 29565 566948
rect 29499 566883 29565 566884
rect 29131 533356 29197 533357
rect 29131 533292 29132 533356
rect 29196 533292 29197 533356
rect 29131 533291 29197 533292
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 29502 342141 29562 566883
rect 31523 557564 31589 557565
rect 31523 557500 31524 557564
rect 31588 557500 31589 557564
rect 31523 557499 31589 557500
rect 31155 549404 31221 549405
rect 31155 549340 31156 549404
rect 31220 549340 31221 549404
rect 31155 549339 31221 549340
rect 30235 546140 30301 546141
rect 30235 546076 30236 546140
rect 30300 546076 30301 546140
rect 30235 546075 30301 546076
rect 30051 536076 30117 536077
rect 30051 536012 30052 536076
rect 30116 536012 30117 536076
rect 30051 536011 30117 536012
rect 29867 533220 29933 533221
rect 29867 533156 29868 533220
rect 29932 533156 29933 533220
rect 29867 533155 29933 533156
rect 29870 484533 29930 533155
rect 29867 484532 29933 484533
rect 29867 484468 29868 484532
rect 29932 484468 29933 484532
rect 29867 484467 29933 484468
rect 30054 483989 30114 536011
rect 30051 483988 30117 483989
rect 30051 483924 30052 483988
rect 30116 483924 30117 483988
rect 30051 483923 30117 483924
rect 30238 448085 30298 546075
rect 30971 534716 31037 534717
rect 30971 534652 30972 534716
rect 31036 534652 31037 534716
rect 30971 534651 31037 534652
rect 30974 485077 31034 534651
rect 30971 485076 31037 485077
rect 30971 485012 30972 485076
rect 31036 485012 31037 485076
rect 30971 485011 31037 485012
rect 30235 448084 30301 448085
rect 30235 448020 30236 448084
rect 30300 448020 30301 448084
rect 30235 448019 30301 448020
rect 31158 447541 31218 549339
rect 31339 544372 31405 544373
rect 31339 544308 31340 544372
rect 31404 544308 31405 544372
rect 31339 544307 31405 544308
rect 31155 447540 31221 447541
rect 31155 447476 31156 447540
rect 31220 447476 31221 447540
rect 31155 447475 31221 447476
rect 31342 440469 31402 544307
rect 31526 448629 31586 557499
rect 31710 534173 31770 671195
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41275 640116 41341 640117
rect 41275 640052 41276 640116
rect 41340 640052 41341 640116
rect 41275 640051 41341 640052
rect 39803 638756 39869 638757
rect 39803 638692 39804 638756
rect 39868 638692 39869 638756
rect 39803 638691 39869 638692
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 33731 557700 33797 557701
rect 33731 557636 33732 557700
rect 33796 557636 33797 557700
rect 33731 557635 33797 557636
rect 32995 550356 33061 550357
rect 32995 550292 32996 550356
rect 33060 550292 33061 550356
rect 32995 550291 33061 550292
rect 32811 540564 32877 540565
rect 32811 540500 32812 540564
rect 32876 540500 32877 540564
rect 32811 540499 32877 540500
rect 32443 536892 32509 536893
rect 32443 536828 32444 536892
rect 32508 536828 32509 536892
rect 32443 536827 32509 536828
rect 31707 534172 31773 534173
rect 31707 534108 31708 534172
rect 31772 534108 31773 534172
rect 31707 534107 31773 534108
rect 32446 483445 32506 536827
rect 32627 535260 32693 535261
rect 32627 535196 32628 535260
rect 32692 535196 32693 535260
rect 32627 535195 32693 535196
rect 32443 483444 32509 483445
rect 32443 483380 32444 483444
rect 32508 483380 32509 483444
rect 32443 483379 32509 483380
rect 31523 448628 31589 448629
rect 31523 448564 31524 448628
rect 31588 448564 31589 448628
rect 31523 448563 31589 448564
rect 32630 443189 32690 535195
rect 32627 443188 32693 443189
rect 32627 443124 32628 443188
rect 32692 443124 32693 443188
rect 32627 443123 32693 443124
rect 31339 440468 31405 440469
rect 31339 440404 31340 440468
rect 31404 440404 31405 440468
rect 31339 440403 31405 440404
rect 32814 439925 32874 540499
rect 32998 445909 33058 550291
rect 33734 494869 33794 557635
rect 33915 556340 33981 556341
rect 33915 556276 33916 556340
rect 33980 556276 33981 556340
rect 33915 556275 33981 556276
rect 33731 494868 33797 494869
rect 33731 494804 33732 494868
rect 33796 494804 33797 494868
rect 33731 494803 33797 494804
rect 33918 486165 33978 556275
rect 34283 548860 34349 548861
rect 34283 548796 34284 548860
rect 34348 548796 34349 548860
rect 34283 548795 34349 548796
rect 34099 522340 34165 522341
rect 34099 522276 34100 522340
rect 34164 522276 34165 522340
rect 34099 522275 34165 522276
rect 33915 486164 33981 486165
rect 33915 486100 33916 486164
rect 33980 486100 33981 486164
rect 33915 486099 33981 486100
rect 32995 445908 33061 445909
rect 32995 445844 32996 445908
rect 33060 445844 33061 445908
rect 32995 445843 33061 445844
rect 34102 444277 34162 522275
rect 34286 450805 34346 548795
rect 37794 543454 38414 578898
rect 39435 549540 39501 549541
rect 39435 549476 39436 549540
rect 39500 549476 39501 549540
rect 39435 549475 39501 549476
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 35755 535124 35821 535125
rect 35755 535060 35756 535124
rect 35820 535060 35821 535124
rect 35755 535059 35821 535060
rect 35203 524108 35269 524109
rect 35203 524044 35204 524108
rect 35268 524044 35269 524108
rect 35203 524043 35269 524044
rect 35206 504117 35266 524043
rect 35387 522204 35453 522205
rect 35387 522140 35388 522204
rect 35452 522140 35453 522204
rect 35387 522139 35453 522140
rect 35203 504116 35269 504117
rect 35203 504052 35204 504116
rect 35268 504052 35269 504116
rect 35203 504051 35269 504052
rect 35390 500853 35450 522139
rect 35571 519892 35637 519893
rect 35571 519828 35572 519892
rect 35636 519828 35637 519892
rect 35571 519827 35637 519828
rect 35387 500852 35453 500853
rect 35387 500788 35388 500852
rect 35452 500788 35453 500852
rect 35387 500787 35453 500788
rect 34283 450804 34349 450805
rect 34283 450740 34284 450804
rect 34348 450740 34349 450804
rect 34283 450739 34349 450740
rect 34099 444276 34165 444277
rect 34099 444212 34100 444276
rect 34164 444212 34165 444276
rect 34099 444211 34165 444212
rect 35574 441013 35634 519827
rect 35571 441012 35637 441013
rect 35571 440948 35572 441012
rect 35636 440948 35637 441012
rect 35571 440947 35637 440948
rect 32811 439924 32877 439925
rect 32811 439860 32812 439924
rect 32876 439860 32877 439924
rect 32811 439859 32877 439860
rect 35758 438293 35818 535059
rect 37043 531452 37109 531453
rect 37043 531388 37044 531452
rect 37108 531388 37109 531452
rect 37043 531387 37109 531388
rect 36491 527236 36557 527237
rect 36491 527172 36492 527236
rect 36556 527172 36557 527236
rect 36491 527171 36557 527172
rect 36494 501397 36554 527171
rect 36675 523428 36741 523429
rect 36675 523364 36676 523428
rect 36740 523364 36741 523428
rect 36675 523363 36741 523364
rect 36491 501396 36557 501397
rect 36491 501332 36492 501396
rect 36556 501332 36557 501396
rect 36491 501331 36557 501332
rect 36678 492149 36738 523363
rect 36859 520980 36925 520981
rect 36859 520916 36860 520980
rect 36924 520916 36925 520980
rect 36859 520915 36925 520916
rect 36675 492148 36741 492149
rect 36675 492084 36676 492148
rect 36740 492084 36741 492148
rect 36675 492083 36741 492084
rect 36862 441557 36922 520915
rect 36859 441556 36925 441557
rect 36859 441492 36860 441556
rect 36924 441492 36925 441556
rect 36859 441491 36925 441492
rect 37046 438837 37106 531387
rect 37227 525876 37293 525877
rect 37227 525812 37228 525876
rect 37292 525812 37293 525876
rect 37227 525811 37293 525812
rect 37230 449717 37290 525811
rect 37411 519620 37477 519621
rect 37411 519556 37412 519620
rect 37476 519556 37477 519620
rect 37411 519555 37477 519556
rect 37227 449716 37293 449717
rect 37227 449652 37228 449716
rect 37292 449652 37293 449716
rect 37227 449651 37293 449652
rect 37414 442101 37474 519555
rect 37794 507454 38414 542898
rect 39251 521796 39317 521797
rect 39251 521732 39252 521796
rect 39316 521732 39317 521796
rect 39251 521731 39317 521732
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 39254 489429 39314 521731
rect 39251 489428 39317 489429
rect 39251 489364 39252 489428
rect 39316 489364 39317 489428
rect 39251 489363 39317 489364
rect 39438 485621 39498 549475
rect 39619 523700 39685 523701
rect 39619 523636 39620 523700
rect 39684 523636 39685 523700
rect 39619 523635 39685 523636
rect 39435 485620 39501 485621
rect 39435 485556 39436 485620
rect 39500 485556 39501 485620
rect 39435 485555 39501 485556
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37411 442100 37477 442101
rect 37411 442036 37412 442100
rect 37476 442036 37477 442100
rect 37411 442035 37477 442036
rect 37043 438836 37109 438837
rect 37043 438772 37044 438836
rect 37108 438772 37109 438836
rect 37043 438771 37109 438772
rect 35755 438292 35821 438293
rect 35755 438228 35756 438292
rect 35820 438228 35821 438292
rect 35755 438227 35821 438228
rect 37794 435454 38414 470898
rect 39622 450261 39682 523635
rect 39806 510101 39866 638691
rect 41091 550764 41157 550765
rect 41091 550700 41092 550764
rect 41156 550700 41157 550764
rect 41091 550699 41157 550700
rect 39803 510100 39869 510101
rect 39803 510036 39804 510100
rect 39868 510036 39869 510100
rect 39803 510035 39869 510036
rect 41094 490109 41154 550699
rect 41278 508469 41338 640051
rect 41514 619174 42134 654618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 44771 645012 44837 645013
rect 44771 644948 44772 645012
rect 44836 644948 44837 645012
rect 44771 644947 44837 644948
rect 44035 644332 44101 644333
rect 44035 644268 44036 644332
rect 44100 644268 44101 644332
rect 44035 644267 44101 644268
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 43851 544236 43917 544237
rect 43851 544172 43852 544236
rect 43916 544172 43917 544236
rect 43851 544171 43917 544172
rect 42379 534852 42445 534853
rect 42379 534788 42380 534852
rect 42444 534788 42445 534852
rect 42379 534787 42445 534788
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41275 508468 41341 508469
rect 41275 508404 41276 508468
rect 41340 508404 41341 508468
rect 41275 508403 41341 508404
rect 41091 490108 41157 490109
rect 41091 490044 41092 490108
rect 41156 490044 41157 490108
rect 41091 490043 41157 490044
rect 41514 475174 42134 510618
rect 42382 483037 42442 534787
rect 43667 522612 43733 522613
rect 43667 522548 43668 522612
rect 43732 522548 43733 522612
rect 43667 522547 43733 522548
rect 42563 520300 42629 520301
rect 42563 520236 42564 520300
rect 42628 520236 42629 520300
rect 42563 520235 42629 520236
rect 42566 499590 42626 520235
rect 43483 519076 43549 519077
rect 43483 519012 43484 519076
rect 43548 519012 43549 519076
rect 43483 519011 43549 519012
rect 43299 510508 43365 510509
rect 43299 510444 43300 510508
rect 43364 510444 43365 510508
rect 43299 510443 43365 510444
rect 42566 499530 42810 499590
rect 42563 491196 42629 491197
rect 42563 491132 42564 491196
rect 42628 491132 42629 491196
rect 42563 491131 42629 491132
rect 42379 483036 42445 483037
rect 42379 482972 42380 483036
rect 42444 482972 42445 483036
rect 42379 482971 42445 482972
rect 42379 482900 42445 482901
rect 42379 482836 42380 482900
rect 42444 482836 42445 482900
rect 42379 482835 42445 482836
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 39619 450260 39685 450261
rect 39619 450196 39620 450260
rect 39684 450196 39685 450260
rect 39619 450195 39685 450196
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 29499 342140 29565 342141
rect 29499 342076 29500 342140
rect 29564 342076 29565 342140
rect 29499 342075 29565 342076
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 42382 416533 42442 482835
rect 42379 416532 42445 416533
rect 42379 416468 42380 416532
rect 42444 416468 42445 416532
rect 42379 416467 42445 416468
rect 42566 413269 42626 491131
rect 42750 490517 42810 499530
rect 42747 490516 42813 490517
rect 42747 490452 42748 490516
rect 42812 490452 42813 490516
rect 42747 490451 42813 490452
rect 43302 415445 43362 510443
rect 43486 491061 43546 519011
rect 43670 505749 43730 522547
rect 43667 505748 43733 505749
rect 43667 505684 43668 505748
rect 43732 505684 43733 505748
rect 43667 505683 43733 505684
rect 43483 491060 43549 491061
rect 43483 490996 43484 491060
rect 43548 490996 43549 491060
rect 43483 490995 43549 490996
rect 43299 415444 43365 415445
rect 43299 415380 43300 415444
rect 43364 415380 43365 415444
rect 43299 415379 43365 415380
rect 43854 414901 43914 544171
rect 44038 509557 44098 644267
rect 44587 518260 44653 518261
rect 44587 518196 44588 518260
rect 44652 518196 44653 518260
rect 44587 518195 44653 518196
rect 44035 509556 44101 509557
rect 44035 509492 44036 509556
rect 44100 509492 44101 509556
rect 44035 509491 44101 509492
rect 44035 505204 44101 505205
rect 44035 505140 44036 505204
rect 44100 505140 44101 505204
rect 44035 505139 44101 505140
rect 44038 415989 44098 505139
rect 44590 488341 44650 518195
rect 44774 510645 44834 644947
rect 44955 635220 45021 635221
rect 44955 635156 44956 635220
rect 45020 635156 45021 635220
rect 44955 635155 45021 635156
rect 44771 510644 44837 510645
rect 44771 510580 44772 510644
rect 44836 510580 44837 510644
rect 44771 510579 44837 510580
rect 44587 488340 44653 488341
rect 44587 488276 44588 488340
rect 44652 488276 44653 488340
rect 44587 488275 44653 488276
rect 44035 415988 44101 415989
rect 44035 415924 44036 415988
rect 44100 415924 44101 415988
rect 44035 415923 44101 415924
rect 43851 414900 43917 414901
rect 43851 414836 43852 414900
rect 43916 414836 43917 414900
rect 43851 414835 43917 414836
rect 44958 414357 45018 635155
rect 45234 622894 45854 658338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 46795 644604 46861 644605
rect 46795 644540 46796 644604
rect 46860 644540 46861 644604
rect 46795 644539 46861 644540
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 46611 552124 46677 552125
rect 46611 552060 46612 552124
rect 46676 552060 46677 552124
rect 46611 552059 46677 552060
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 46427 519212 46493 519213
rect 46427 519148 46428 519212
rect 46492 519148 46493 519212
rect 46427 519147 46493 519148
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 46430 499085 46490 519147
rect 46427 499084 46493 499085
rect 46427 499020 46428 499084
rect 46492 499020 46493 499084
rect 46427 499019 46493 499020
rect 46243 498268 46309 498269
rect 46243 498204 46244 498268
rect 46308 498204 46309 498268
rect 46243 498203 46309 498204
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 46246 457877 46306 498203
rect 46243 457876 46309 457877
rect 46243 457812 46244 457876
rect 46308 457812 46309 457876
rect 46243 457811 46309 457812
rect 46427 456924 46493 456925
rect 46427 456860 46428 456924
rect 46492 456860 46493 456924
rect 46427 456859 46493 456860
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 44955 414356 45021 414357
rect 44955 414292 44956 414356
rect 45020 414292 45021 414356
rect 44955 414291 45021 414292
rect 42563 413268 42629 413269
rect 42563 413204 42564 413268
rect 42628 413204 42629 413268
rect 42563 413203 42629 413204
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 406894 45854 442338
rect 46430 413813 46490 456859
rect 46614 445365 46674 552059
rect 46798 457333 46858 644539
rect 48635 642292 48701 642293
rect 48635 642228 48636 642292
rect 48700 642228 48701 642292
rect 48635 642227 48701 642228
rect 48451 635628 48517 635629
rect 48451 635564 48452 635628
rect 48516 635564 48517 635628
rect 48451 635563 48517 635564
rect 48083 634812 48149 634813
rect 48083 634748 48084 634812
rect 48148 634748 48149 634812
rect 48083 634747 48149 634748
rect 47899 559332 47965 559333
rect 47899 559268 47900 559332
rect 47964 559268 47965 559332
rect 47899 559267 47965 559268
rect 47715 559196 47781 559197
rect 47715 559132 47716 559196
rect 47780 559132 47781 559196
rect 47715 559131 47781 559132
rect 47531 553484 47597 553485
rect 47531 553420 47532 553484
rect 47596 553420 47597 553484
rect 47531 553419 47597 553420
rect 46795 457332 46861 457333
rect 46795 457268 46796 457332
rect 46860 457268 46861 457332
rect 46795 457267 46861 457268
rect 47534 452437 47594 553419
rect 47531 452436 47597 452437
rect 47531 452372 47532 452436
rect 47596 452372 47597 452436
rect 47531 452371 47597 452372
rect 47718 451893 47778 559131
rect 47715 451892 47781 451893
rect 47715 451828 47716 451892
rect 47780 451828 47781 451892
rect 47715 451827 47781 451828
rect 47902 446453 47962 559267
rect 48086 452981 48146 634747
rect 48454 455157 48514 635563
rect 48451 455156 48517 455157
rect 48451 455092 48452 455156
rect 48516 455092 48517 455156
rect 48451 455091 48517 455092
rect 48638 454069 48698 642227
rect 48954 626614 49574 662058
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 55995 700364 56061 700365
rect 55995 700300 55996 700364
rect 56060 700300 56061 700364
rect 55995 700299 56061 700300
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52315 644740 52381 644741
rect 52315 644676 52316 644740
rect 52380 644676 52381 644740
rect 52315 644675 52381 644676
rect 50843 641068 50909 641069
rect 50843 641004 50844 641068
rect 50908 641004 50909 641068
rect 50843 641003 50909 641004
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 50475 520708 50541 520709
rect 50475 520644 50476 520708
rect 50540 520644 50541 520708
rect 50475 520643 50541 520644
rect 50291 519348 50357 519349
rect 50291 519284 50292 519348
rect 50356 519284 50357 519348
rect 50291 519283 50357 519284
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 50294 507925 50354 519283
rect 50291 507924 50357 507925
rect 50291 507860 50292 507924
rect 50356 507860 50357 507924
rect 50291 507859 50357 507860
rect 50478 505069 50538 520643
rect 50659 518396 50725 518397
rect 50659 518332 50660 518396
rect 50724 518332 50725 518396
rect 50659 518331 50725 518332
rect 50475 505068 50541 505069
rect 50475 505004 50476 505068
rect 50540 505004 50541 505068
rect 50475 505003 50541 505004
rect 50662 496773 50722 518331
rect 50659 496772 50725 496773
rect 50659 496708 50660 496772
rect 50724 496708 50725 496772
rect 50659 496707 50725 496708
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48635 454068 48701 454069
rect 48635 454004 48636 454068
rect 48700 454004 48701 454068
rect 48635 454003 48701 454004
rect 48083 452980 48149 452981
rect 48083 452916 48084 452980
rect 48148 452916 48149 452980
rect 48083 452915 48149 452916
rect 48954 446614 49574 482058
rect 50846 456245 50906 641003
rect 52131 636580 52197 636581
rect 52131 636516 52132 636580
rect 52196 636516 52197 636580
rect 52131 636515 52197 636516
rect 52134 492693 52194 636515
rect 52131 492692 52197 492693
rect 52131 492628 52132 492692
rect 52196 492628 52197 492692
rect 52131 492627 52197 492628
rect 50843 456244 50909 456245
rect 50843 456180 50844 456244
rect 50908 456180 50909 456244
rect 50843 456179 50909 456180
rect 52318 453525 52378 644675
rect 52674 630334 53294 665778
rect 55075 657660 55141 657661
rect 55075 657596 55076 657660
rect 55140 657596 55141 657660
rect 55075 657595 55141 657596
rect 54707 642564 54773 642565
rect 54707 642500 54708 642564
rect 54772 642500 54773 642564
rect 54707 642499 54773 642500
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 54523 564364 54589 564365
rect 54523 564300 54524 564364
rect 54588 564300 54589 564364
rect 54523 564299 54589 564300
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52674 522334 53294 557778
rect 53603 556476 53669 556477
rect 53603 556412 53604 556476
rect 53668 556412 53669 556476
rect 53603 556411 53669 556412
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52315 453524 52381 453525
rect 52315 453460 52316 453524
rect 52380 453460 52381 453524
rect 52315 453459 52381 453460
rect 47899 446452 47965 446453
rect 47899 446388 47900 446452
rect 47964 446388 47965 446452
rect 47899 446387 47965 446388
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 46611 445364 46677 445365
rect 46611 445300 46612 445364
rect 46676 445300 46677 445364
rect 46611 445299 46677 445300
rect 46427 413812 46493 413813
rect 46427 413748 46428 413812
rect 46492 413748 46493 413812
rect 46427 413747 46493 413748
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48083 344588 48149 344589
rect 48083 344524 48084 344588
rect 48148 344524 48149 344588
rect 48083 344523 48149 344524
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 48086 245037 48146 344523
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48635 254148 48701 254149
rect 48635 254084 48636 254148
rect 48700 254084 48701 254148
rect 48635 254083 48701 254084
rect 48083 245036 48149 245037
rect 48083 244972 48084 245036
rect 48148 244972 48149 245036
rect 48083 244971 48149 244972
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 48451 201924 48517 201925
rect 48451 201860 48452 201924
rect 48516 201860 48517 201924
rect 48451 201859 48517 201860
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 48454 140453 48514 201859
rect 48638 140725 48698 254083
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48635 140724 48701 140725
rect 48635 140660 48636 140724
rect 48700 140660 48701 140724
rect 48635 140659 48701 140660
rect 48451 140452 48517 140453
rect 48451 140388 48452 140452
rect 48516 140388 48517 140452
rect 48451 140387 48517 140388
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 414334 53294 449778
rect 53606 439381 53666 556411
rect 54526 518941 54586 564299
rect 54523 518940 54589 518941
rect 54523 518876 54524 518940
rect 54588 518876 54589 518940
rect 54523 518875 54589 518876
rect 54523 517988 54589 517989
rect 54523 517924 54524 517988
rect 54588 517924 54589 517988
rect 54523 517923 54589 517924
rect 54526 506837 54586 517923
rect 54523 506836 54589 506837
rect 54523 506772 54524 506836
rect 54588 506772 54589 506836
rect 54523 506771 54589 506772
rect 54710 476917 54770 642499
rect 54891 572388 54957 572389
rect 54891 572324 54892 572388
rect 54956 572324 54957 572388
rect 54891 572323 54957 572324
rect 54894 558245 54954 572323
rect 54891 558244 54957 558245
rect 54891 558180 54892 558244
rect 54956 558180 54957 558244
rect 54891 558179 54957 558180
rect 54891 519620 54957 519621
rect 54891 519556 54892 519620
rect 54956 519556 54957 519620
rect 54891 519555 54957 519556
rect 54707 476916 54773 476917
rect 54707 476852 54708 476916
rect 54772 476852 54773 476916
rect 54707 476851 54773 476852
rect 53603 439380 53669 439381
rect 53603 439316 53604 439380
rect 53668 439316 53669 439380
rect 53603 439315 53669 439316
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 54894 260133 54954 519555
rect 55078 387565 55138 657595
rect 55811 640388 55877 640389
rect 55811 640324 55812 640388
rect 55876 640324 55877 640388
rect 55811 640323 55877 640324
rect 55627 632092 55693 632093
rect 55627 632028 55628 632092
rect 55692 632028 55693 632092
rect 55627 632027 55693 632028
rect 55443 556612 55509 556613
rect 55443 556548 55444 556612
rect 55508 556548 55509 556612
rect 55443 556547 55509 556548
rect 55446 487797 55506 556547
rect 55630 529821 55690 632027
rect 55627 529820 55693 529821
rect 55627 529756 55628 529820
rect 55692 529756 55693 529820
rect 55627 529755 55693 529756
rect 55814 523021 55874 640323
rect 55998 558925 56058 700299
rect 56394 670054 57014 709082
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 59123 699820 59189 699821
rect 59123 699756 59124 699820
rect 59188 699756 59189 699820
rect 59123 699755 59189 699756
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 634054 57014 669498
rect 58939 639844 59005 639845
rect 58939 639780 58940 639844
rect 59004 639780 59005 639844
rect 58939 639779 59005 639780
rect 58755 637532 58821 637533
rect 58755 637468 58756 637532
rect 58820 637468 58821 637532
rect 58755 637467 58821 637468
rect 58571 636852 58637 636853
rect 58571 636788 58572 636852
rect 58636 636788 58637 636852
rect 58571 636787 58637 636788
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 57835 632092 57901 632093
rect 57835 632028 57836 632092
rect 57900 632028 57901 632092
rect 57835 632027 57901 632028
rect 57651 631004 57717 631005
rect 57651 630940 57652 631004
rect 57716 630940 57717 631004
rect 57651 630939 57717 630940
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 55995 558924 56061 558925
rect 55995 558860 55996 558924
rect 56060 558860 56061 558924
rect 55995 558859 56061 558860
rect 55995 529004 56061 529005
rect 55995 528940 55996 529004
rect 56060 528940 56061 529004
rect 55995 528939 56061 528940
rect 55811 523020 55877 523021
rect 55811 522956 55812 523020
rect 55876 522956 55877 523020
rect 55811 522955 55877 522956
rect 55998 522610 56058 528939
rect 55630 522550 56058 522610
rect 56394 526054 57014 561498
rect 57654 553349 57714 630939
rect 57651 553348 57717 553349
rect 57651 553284 57652 553348
rect 57716 553284 57717 553348
rect 57651 553283 57717 553284
rect 57838 547637 57898 632027
rect 57835 547636 57901 547637
rect 57835 547572 57836 547636
rect 57900 547572 57901 547636
rect 57835 547571 57901 547572
rect 57835 529412 57901 529413
rect 57835 529348 57836 529412
rect 57900 529348 57901 529412
rect 57835 529347 57901 529348
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 55630 505205 55690 522550
rect 55995 522476 56061 522477
rect 55995 522412 55996 522476
rect 56060 522412 56061 522476
rect 55995 522411 56061 522412
rect 55627 505204 55693 505205
rect 55627 505140 55628 505204
rect 55692 505140 55693 505204
rect 55627 505139 55693 505140
rect 55443 487796 55509 487797
rect 55443 487732 55444 487796
rect 55508 487732 55509 487796
rect 55443 487731 55509 487732
rect 55998 446997 56058 522411
rect 56394 490054 57014 525498
rect 57651 519620 57717 519621
rect 57651 519556 57652 519620
rect 57716 519556 57717 519620
rect 57651 519555 57717 519556
rect 57467 505068 57533 505069
rect 57467 505004 57468 505068
rect 57532 505004 57533 505068
rect 57467 505003 57533 505004
rect 57470 499590 57530 505003
rect 57286 499530 57530 499590
rect 57286 498677 57346 499530
rect 57467 499084 57533 499085
rect 57467 499020 57468 499084
rect 57532 499020 57533 499084
rect 57467 499019 57533 499020
rect 57283 498676 57349 498677
rect 57283 498612 57284 498676
rect 57348 498612 57349 498676
rect 57283 498611 57349 498612
rect 57283 496772 57349 496773
rect 57283 496708 57284 496772
rect 57348 496708 57349 496772
rect 57283 496707 57349 496708
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 57286 488885 57346 496707
rect 57470 495957 57530 499019
rect 57467 495956 57533 495957
rect 57467 495892 57468 495956
rect 57532 495892 57533 495956
rect 57467 495891 57533 495892
rect 57283 488884 57349 488885
rect 57283 488820 57284 488884
rect 57348 488820 57349 488884
rect 57283 488819 57349 488820
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 55995 446996 56061 446997
rect 55995 446932 55996 446996
rect 56060 446932 56061 446996
rect 55995 446931 56061 446932
rect 56394 418054 57014 453498
rect 57654 443733 57714 519555
rect 57838 514997 57898 529347
rect 58574 523837 58634 636787
rect 58571 523836 58637 523837
rect 58571 523772 58572 523836
rect 58636 523772 58637 523836
rect 58571 523771 58637 523772
rect 58387 523156 58453 523157
rect 58387 523092 58388 523156
rect 58452 523092 58453 523156
rect 58387 523091 58453 523092
rect 57835 514996 57901 514997
rect 57835 514932 57836 514996
rect 57900 514932 57901 514996
rect 57835 514931 57901 514932
rect 58390 451349 58450 523091
rect 58571 518668 58637 518669
rect 58571 518604 58572 518668
rect 58636 518604 58637 518668
rect 58571 518603 58637 518604
rect 58387 451348 58453 451349
rect 58387 451284 58388 451348
rect 58452 451284 58453 451348
rect 58387 451283 58453 451284
rect 58574 449173 58634 518603
rect 58758 517581 58818 637467
rect 58942 521661 59002 639779
rect 59126 560421 59186 699755
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 633097 60734 637218
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 634540 64454 640938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 633097 74414 650898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 633097 78134 654618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 633097 81854 658338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 633097 85574 662058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 633097 89294 665778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 633097 93014 633498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 96114 633097 96734 637218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 633097 100454 640938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 634540 110414 650898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 633097 114134 654618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 633097 117854 658338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 633097 121574 662058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 121867 634404 121933 634405
rect 121867 634340 121868 634404
rect 121932 634340 121933 634404
rect 121867 634339 121933 634340
rect 121870 633861 121930 634339
rect 121867 633860 121933 633861
rect 121867 633796 121868 633860
rect 121932 633796 121933 633860
rect 121867 633795 121933 633796
rect 124674 633097 125294 665778
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 633097 129014 633498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 633097 132734 637218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 59675 627808 59741 627809
rect 59675 627744 59676 627808
rect 59740 627744 59741 627808
rect 59675 627743 59741 627744
rect 59123 560420 59189 560421
rect 59123 560356 59124 560420
rect 59188 560356 59189 560420
rect 59123 560355 59189 560356
rect 59123 548996 59189 548997
rect 59123 548932 59124 548996
rect 59188 548932 59189 548996
rect 59123 548931 59189 548932
rect 58939 521660 59005 521661
rect 58939 521596 58940 521660
rect 59004 521596 59005 521660
rect 58939 521595 59005 521596
rect 58755 517580 58821 517581
rect 58755 517516 58756 517580
rect 58820 517516 58821 517580
rect 58755 517515 58821 517516
rect 59126 512010 59186 548931
rect 59678 546413 59738 627743
rect 59859 626720 59925 626721
rect 59859 626656 59860 626720
rect 59924 626656 59925 626720
rect 59859 626655 59925 626656
rect 59675 546412 59741 546413
rect 59675 546348 59676 546412
rect 59740 546348 59741 546412
rect 59675 546347 59741 546348
rect 59675 545868 59741 545869
rect 59675 545804 59676 545868
rect 59740 545804 59741 545868
rect 59675 545803 59741 545804
rect 59491 523020 59557 523021
rect 59491 522956 59492 523020
rect 59556 522956 59557 523020
rect 59491 522955 59557 522956
rect 59307 521116 59373 521117
rect 59307 521052 59308 521116
rect 59372 521052 59373 521116
rect 59307 521051 59373 521052
rect 58758 511950 59186 512010
rect 58758 502485 58818 511950
rect 59310 506970 59370 521051
rect 58942 506910 59370 506970
rect 58755 502484 58821 502485
rect 58755 502420 58756 502484
rect 58820 502420 58821 502484
rect 58755 502419 58821 502420
rect 58571 449172 58637 449173
rect 58571 449108 58572 449172
rect 58636 449108 58637 449172
rect 58571 449107 58637 449108
rect 57651 443732 57717 443733
rect 57651 443668 57652 443732
rect 57716 443668 57717 443732
rect 57651 443667 57717 443668
rect 58942 442645 59002 506910
rect 59494 504661 59554 522955
rect 59491 504660 59557 504661
rect 59491 504596 59492 504660
rect 59556 504596 59557 504660
rect 59491 504595 59557 504596
rect 59123 502352 59189 502353
rect 59123 502288 59124 502352
rect 59188 502288 59189 502352
rect 59123 502287 59189 502288
rect 59126 444821 59186 502287
rect 59678 454613 59738 545803
rect 59862 522613 59922 626655
rect 79568 619174 79888 619206
rect 79568 618938 79610 619174
rect 79846 618938 79888 619174
rect 79568 618854 79888 618938
rect 79568 618618 79610 618854
rect 79846 618618 79888 618854
rect 79568 618586 79888 618618
rect 110288 619174 110608 619206
rect 110288 618938 110330 619174
rect 110566 618938 110608 619174
rect 110288 618854 110608 618938
rect 110288 618618 110330 618854
rect 110566 618618 110608 618854
rect 110288 618586 110608 618618
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 125648 615454 125968 615486
rect 125648 615218 125690 615454
rect 125926 615218 125968 615454
rect 125648 615134 125968 615218
rect 125648 614898 125690 615134
rect 125926 614898 125968 615134
rect 125648 614866 125968 614898
rect 135834 605494 136454 640938
rect 135834 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 136454 605494
rect 135834 605174 136454 605258
rect 135834 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 136454 605174
rect 79568 583174 79888 583206
rect 79568 582938 79610 583174
rect 79846 582938 79888 583174
rect 79568 582854 79888 582938
rect 79568 582618 79610 582854
rect 79846 582618 79888 582854
rect 79568 582586 79888 582618
rect 110288 583174 110608 583206
rect 110288 582938 110330 583174
rect 110566 582938 110608 583174
rect 110288 582854 110608 582938
rect 110288 582618 110330 582854
rect 110566 582618 110608 582854
rect 110288 582586 110608 582618
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 125648 579454 125968 579486
rect 125648 579218 125690 579454
rect 125926 579218 125968 579454
rect 125648 579134 125968 579218
rect 125648 578898 125690 579134
rect 125926 578898 125968 579134
rect 125648 578866 125968 578898
rect 135834 569494 136454 604938
rect 135834 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 136454 569494
rect 135834 569174 136454 569258
rect 135834 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 136454 569174
rect 60411 564704 60477 564705
rect 60411 564640 60412 564704
rect 60476 564640 60477 564704
rect 60411 564639 60477 564640
rect 60414 558789 60474 564639
rect 60595 562528 60661 562529
rect 60595 562464 60596 562528
rect 60660 562464 60661 562528
rect 60595 562463 60661 562464
rect 60598 558925 60658 562463
rect 60595 558924 60661 558925
rect 60595 558860 60596 558924
rect 60660 558860 60661 558924
rect 60595 558859 60661 558860
rect 60411 558788 60477 558789
rect 60411 558724 60412 558788
rect 60476 558724 60477 558788
rect 60411 558723 60477 558724
rect 60114 529774 60734 558575
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 59859 522612 59925 522613
rect 59859 522548 59860 522612
rect 59924 522548 59925 522612
rect 59859 522547 59925 522548
rect 60114 493774 60734 529218
rect 73794 543454 74414 558575
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 64208 471454 64528 471486
rect 64208 471218 64250 471454
rect 64486 471218 64528 471454
rect 64208 471134 64528 471218
rect 64208 470898 64250 471134
rect 64486 470898 64528 471134
rect 64208 470866 64528 470898
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 59675 454612 59741 454613
rect 59675 454548 59676 454612
rect 59740 454548 59741 454612
rect 59675 454547 59741 454548
rect 59123 444820 59189 444821
rect 59123 444756 59124 444820
rect 59188 444756 59189 444820
rect 59123 444755 59189 444756
rect 58939 442644 59005 442645
rect 58939 442580 58940 442644
rect 59004 442580 59005 442644
rect 58939 442579 59005 442580
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 55075 387564 55141 387565
rect 55075 387500 55076 387564
rect 55140 387500 55141 387564
rect 55075 387499 55141 387500
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 54891 260132 54957 260133
rect 54891 260068 54892 260132
rect 54956 260068 54957 260132
rect 54891 260067 54957 260068
rect 54208 255454 54528 255486
rect 54208 255218 54250 255454
rect 54486 255218 54528 255454
rect 54208 255134 54528 255218
rect 54208 254898 54250 255134
rect 54486 254898 54528 255134
rect 54208 254866 54528 254898
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 56394 238054 57014 273498
rect 60114 421774 60734 457218
rect 64208 435454 64528 435486
rect 64208 435218 64250 435454
rect 64486 435218 64528 435454
rect 64208 435134 64528 435218
rect 64208 434898 64250 435134
rect 64486 434898 64528 435134
rect 64208 434866 64528 434898
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 64208 399454 64528 399486
rect 64208 399218 64250 399454
rect 64486 399218 64528 399454
rect 64208 399134 64528 399218
rect 64208 398898 64250 399134
rect 64486 398898 64528 399134
rect 64208 398866 64528 398898
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 260449 60734 277218
rect 63834 389494 64454 389988
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 281494 64454 316938
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 63834 260449 64454 280938
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 260449 74414 290898
rect 77514 547174 78134 558575
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 81234 550894 81854 558575
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 79568 511174 79888 511206
rect 79568 510938 79610 511174
rect 79846 510938 79888 511174
rect 79568 510854 79888 510938
rect 79568 510618 79610 510854
rect 79846 510618 79888 510854
rect 79568 510586 79888 510618
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 79568 475174 79888 475206
rect 79568 474938 79610 475174
rect 79846 474938 79888 475174
rect 79568 474854 79888 474938
rect 79568 474618 79610 474854
rect 79846 474618 79888 474854
rect 79568 474586 79888 474618
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 79568 439174 79888 439206
rect 79568 438938 79610 439174
rect 79846 438938 79888 439174
rect 79568 438854 79888 438938
rect 79568 438618 79610 438854
rect 79846 438618 79888 438854
rect 79568 438586 79888 438618
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 79568 403174 79888 403206
rect 79568 402938 79610 403174
rect 79846 402938 79888 403174
rect 79568 402854 79888 402938
rect 79568 402618 79610 402854
rect 79846 402618 79888 402854
rect 79568 402586 79888 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 260449 78134 294618
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 260449 81854 262338
rect 84954 554614 85574 558575
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 260449 85574 266058
rect 88674 558334 89294 558575
rect 88674 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 89294 558334
rect 88674 558014 89294 558098
rect 88674 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 89294 558014
rect 88674 522334 89294 557778
rect 88674 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 89294 522334
rect 88674 522014 89294 522098
rect 88674 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 89294 522014
rect 88674 486334 89294 521778
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 88674 450334 89294 485778
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 414334 89294 449778
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 306334 89294 341778
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 88674 270334 89294 305778
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 88674 260449 89294 269778
rect 92394 526054 93014 558575
rect 92394 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 93014 526054
rect 92394 525734 93014 525818
rect 92394 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 93014 525734
rect 92394 490054 93014 525498
rect 96114 529774 96734 558575
rect 96114 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 96734 529774
rect 96114 529454 96734 529538
rect 96114 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 96734 529454
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 92394 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 93014 490054
rect 92394 489734 93014 489818
rect 92394 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 93014 489734
rect 92394 454054 93014 489498
rect 96114 493774 96734 529218
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 94928 471454 95248 471486
rect 94928 471218 94970 471454
rect 95206 471218 95248 471454
rect 94928 471134 95248 471218
rect 94928 470898 94970 471134
rect 95206 470898 95248 471134
rect 94928 470866 95248 470898
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 418054 93014 453498
rect 96114 457774 96734 493218
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 94928 435454 95248 435486
rect 94928 435218 94970 435454
rect 95206 435218 95248 435454
rect 94928 435134 95248 435218
rect 94928 434898 94970 435134
rect 95206 434898 95248 435134
rect 94928 434866 95248 434898
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 96114 421774 96734 457218
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 94928 399454 95248 399486
rect 94928 399218 94970 399454
rect 95206 399218 95248 399454
rect 94928 399134 95248 399218
rect 94928 398898 94970 399134
rect 95206 398898 95248 399134
rect 94928 398866 95248 398898
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 310054 93014 345498
rect 92394 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 93014 310054
rect 92394 309734 93014 309818
rect 92394 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 93014 309734
rect 92394 274054 93014 309498
rect 92394 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 93014 274054
rect 92394 273734 93014 273818
rect 92394 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 93014 273734
rect 92394 260449 93014 273498
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 313774 96734 349218
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 96114 277774 96734 313218
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 96114 260449 96734 277218
rect 99834 533494 100454 558575
rect 99834 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 100454 533494
rect 99834 533174 100454 533258
rect 99834 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 100454 533174
rect 99834 497494 100454 532938
rect 113514 547174 114134 558575
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 110288 511174 110608 511206
rect 110288 510938 110330 511174
rect 110566 510938 110608 511174
rect 110288 510854 110608 510938
rect 110288 510618 110330 510854
rect 110566 510618 110608 510854
rect 110288 510586 110608 510618
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 99834 461494 100454 496938
rect 110288 475174 110608 475206
rect 110288 474938 110330 475174
rect 110566 474938 110608 475174
rect 110288 474854 110608 474938
rect 110288 474618 110330 474854
rect 110566 474618 110608 474854
rect 110288 474586 110608 474618
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 425494 100454 460938
rect 110288 439174 110608 439206
rect 110288 438938 110330 439174
rect 110566 438938 110608 439174
rect 110288 438854 110608 438938
rect 110288 438618 110330 438854
rect 110566 438618 110608 438854
rect 110288 438586 110608 438618
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 110288 403174 110608 403206
rect 110288 402938 110330 403174
rect 110566 402938 110608 403174
rect 110288 402854 110608 402938
rect 110288 402618 110330 402854
rect 110566 402618 110608 402854
rect 110288 402586 110608 402618
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 317494 100454 352938
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 99834 281494 100454 316938
rect 99834 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 100454 281494
rect 99834 281174 100454 281258
rect 99834 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 100454 281174
rect 99834 260449 100454 280938
rect 109794 363454 110414 389988
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 260449 110414 290898
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 84928 255454 85248 255486
rect 84928 255218 84970 255454
rect 85206 255218 85248 255454
rect 84928 255134 85248 255218
rect 84928 254898 84970 255134
rect 85206 254898 85248 255134
rect 84928 254866 85248 254898
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 54208 219454 54528 219486
rect 54208 219218 54250 219454
rect 54486 219218 54528 219454
rect 54208 219134 54528 219218
rect 54208 218898 54250 219134
rect 54486 218898 54528 219134
rect 54208 218866 54528 218898
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 56394 202054 57014 237498
rect 69568 223174 69888 223206
rect 69568 222938 69610 223174
rect 69846 222938 69888 223174
rect 69568 222854 69888 222938
rect 69568 222618 69610 222854
rect 69846 222618 69888 222854
rect 69568 222586 69888 222618
rect 100288 223174 100608 223206
rect 100288 222938 100330 223174
rect 100566 222938 100608 223174
rect 100288 222854 100608 222938
rect 100288 222618 100330 222854
rect 100566 222618 100608 222854
rect 100288 222586 100608 222618
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 84928 219454 85248 219486
rect 84928 219218 84970 219454
rect 85206 219218 85248 219454
rect 84928 219134 85248 219218
rect 84928 218898 84970 219134
rect 85206 218898 85248 219134
rect 84928 218866 85248 218898
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 130054 57014 165498
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 56394 94054 57014 129498
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 55038 75454 55358 75486
rect 55038 75218 55080 75454
rect 55316 75218 55358 75454
rect 55038 75134 55358 75218
rect 55038 74898 55080 75134
rect 55316 74898 55358 75134
rect 55038 74866 55358 74898
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 58054 57014 93498
rect 60114 169774 60734 198167
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 97774 60734 133218
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 59132 79174 59452 79206
rect 59132 78938 59174 79174
rect 59410 78938 59452 79174
rect 59132 78854 59452 78938
rect 59132 78618 59174 78854
rect 59410 78618 59452 78854
rect 59132 78586 59452 78618
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 61774 60734 97218
rect 63834 173494 64454 198167
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 63834 137494 64454 172938
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 63834 101494 64454 136938
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63226 75454 63546 75486
rect 63226 75218 63268 75454
rect 63504 75218 63546 75454
rect 63226 75134 63546 75218
rect 63226 74898 63268 75134
rect 63504 74898 63546 75134
rect 63226 74866 63546 74898
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 65494 64454 100938
rect 73794 183454 74414 198167
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 67320 79174 67640 79206
rect 67320 78938 67362 79174
rect 67598 78938 67640 79174
rect 67320 78854 67640 78938
rect 67320 78618 67362 78854
rect 67598 78618 67640 78854
rect 67320 78586 67640 78618
rect 71414 75454 71734 75486
rect 71414 75218 71456 75454
rect 71692 75218 71734 75454
rect 71414 75134 71734 75218
rect 71414 74898 71456 75134
rect 71692 74898 71734 75134
rect 71414 74866 71734 74898
rect 73794 75454 74414 110898
rect 77514 187174 78134 198167
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 75508 79174 75828 79206
rect 75508 78938 75550 79174
rect 75786 78938 75828 79174
rect 75508 78854 75828 78938
rect 75508 78618 75550 78854
rect 75786 78618 75828 78854
rect 75508 78586 75828 78618
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 78618
rect 81234 190894 81854 198167
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 79602 75454 79922 75486
rect 79602 75218 79644 75454
rect 79880 75218 79922 75454
rect 79602 75134 79922 75218
rect 79602 74898 79644 75134
rect 79880 74898 79922 75134
rect 79602 74866 79922 74898
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 82338
rect 84954 194614 85574 198167
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 83696 79174 84016 79206
rect 83696 78938 83738 79174
rect 83974 78938 84016 79174
rect 83696 78854 84016 78938
rect 83696 78618 83738 78854
rect 83974 78618 84016 78854
rect 83696 78586 84016 78618
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 162334 89294 198167
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 88674 126334 89294 161778
rect 88674 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 89294 126334
rect 88674 126014 89294 126098
rect 88674 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 89294 126014
rect 88674 90334 89294 125778
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 88674 54334 89294 89778
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 166054 93014 198167
rect 92394 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 93014 166054
rect 92394 165734 93014 165818
rect 92394 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 93014 165734
rect 92394 130054 93014 165498
rect 92394 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 93014 130054
rect 92394 129734 93014 129818
rect 92394 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 93014 129734
rect 92394 94054 93014 129498
rect 92394 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 93014 94054
rect 92394 93734 93014 93818
rect 92394 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 93014 93734
rect 92394 58054 93014 93498
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 169774 96734 198167
rect 96114 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 96734 169774
rect 96114 169454 96734 169538
rect 96114 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 96734 169454
rect 96114 133774 96734 169218
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 96114 97774 96734 133218
rect 96114 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 96734 97774
rect 96114 97454 96734 97538
rect 96114 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 96734 97454
rect 96114 61774 96734 97218
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 96114 25774 96734 61218
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 173494 100454 198167
rect 99834 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 100454 173494
rect 99834 173174 100454 173258
rect 99834 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 100454 173174
rect 99834 137494 100454 172938
rect 99834 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 100454 137494
rect 99834 137174 100454 137258
rect 99834 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 100454 137174
rect 99834 101494 100454 136938
rect 99834 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 100454 101494
rect 99834 101174 100454 101258
rect 99834 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 100454 101174
rect 99834 65494 100454 100938
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 99834 29494 100454 64938
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 183454 110414 198167
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 187174 114134 222618
rect 117234 550894 117854 558575
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 116531 212260 116597 212261
rect 116531 212196 116532 212260
rect 116596 212196 116597 212260
rect 116531 212195 116597 212196
rect 116534 199205 116594 212195
rect 116531 199204 116597 199205
rect 116531 199140 116532 199204
rect 116596 199140 116597 199204
rect 116531 199139 116597 199140
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 554614 121574 558575
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 124674 558334 125294 558575
rect 124674 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 125294 558334
rect 124674 558014 125294 558098
rect 124674 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 125294 558014
rect 124674 522334 125294 557778
rect 124674 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 125294 522334
rect 124674 522014 125294 522098
rect 124674 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 125294 522014
rect 124674 486334 125294 521778
rect 135834 533494 136454 568938
rect 135834 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 136454 533494
rect 135834 533174 136454 533258
rect 135834 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 136454 533174
rect 135834 519809 136454 532938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 519809 146414 542898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 519809 150134 546618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 519809 153854 550338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 519809 157574 554058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 594334 161294 629778
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164003 620260 164069 620261
rect 164003 620196 164004 620260
rect 164068 620196 164069 620260
rect 164003 620195 164069 620196
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 160674 558334 161294 593778
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 160674 522334 161294 557778
rect 164006 551037 164066 620195
rect 164394 598054 165014 633498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 170995 657524 171061 657525
rect 170995 657460 170996 657524
rect 171060 657460 171061 657524
rect 170995 657459 171061 657460
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 166763 614820 166829 614821
rect 166763 614756 166764 614820
rect 166828 614756 166829 614820
rect 166763 614755 166829 614756
rect 165475 608292 165541 608293
rect 165475 608228 165476 608292
rect 165540 608228 165541 608292
rect 165475 608227 165541 608228
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 164394 562054 165014 597498
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 164003 551036 164069 551037
rect 164003 550972 164004 551036
rect 164068 550972 164069 551036
rect 164003 550971 164069 550972
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 160674 519809 161294 521778
rect 164394 526054 165014 561498
rect 165478 537437 165538 608227
rect 166766 552805 166826 614755
rect 168114 601774 168734 637218
rect 170259 611284 170325 611285
rect 170259 611220 170260 611284
rect 170324 611220 170325 611284
rect 170259 611219 170325 611220
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 169523 571164 169589 571165
rect 169523 571100 169524 571164
rect 169588 571100 169589 571164
rect 169523 571099 169589 571100
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 166763 552804 166829 552805
rect 166763 552740 166764 552804
rect 166828 552740 166829 552804
rect 166763 552739 166829 552740
rect 165475 537436 165541 537437
rect 165475 537372 165476 537436
rect 165540 537372 165541 537436
rect 165475 537371 165541 537372
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 164394 519809 165014 525498
rect 168114 529774 168734 565218
rect 169526 551581 169586 571099
rect 169523 551580 169589 551581
rect 169523 551516 169524 551580
rect 169588 551516 169589 551580
rect 169523 551515 169589 551516
rect 170262 547773 170322 611219
rect 170998 553213 171058 657459
rect 171834 641494 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 179275 643244 179341 643245
rect 179275 643180 179276 643244
rect 179340 643180 179341 643244
rect 179275 643179 179341 643180
rect 177251 641748 177317 641749
rect 177251 641684 177252 641748
rect 177316 641684 177317 641748
rect 177251 641683 177317 641684
rect 179091 641748 179157 641749
rect 179091 641684 179092 641748
rect 179156 641684 179157 641748
rect 179091 641683 179157 641684
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 177254 621349 177314 641683
rect 178907 636988 178973 636989
rect 178907 636924 178908 636988
rect 178972 636924 178973 636988
rect 178907 636923 178973 636924
rect 177619 636444 177685 636445
rect 177619 636380 177620 636444
rect 177684 636380 177685 636444
rect 177619 636379 177685 636380
rect 177435 633452 177501 633453
rect 177435 633388 177436 633452
rect 177500 633388 177501 633452
rect 177435 633387 177501 633388
rect 177438 623525 177498 633387
rect 177435 623524 177501 623525
rect 177435 623460 177436 623524
rect 177500 623460 177501 623524
rect 177435 623459 177501 623460
rect 177251 621348 177317 621349
rect 177251 621284 177252 621348
rect 177316 621284 177317 621348
rect 177251 621283 177317 621284
rect 177622 619173 177682 636379
rect 177803 635084 177869 635085
rect 177803 635020 177804 635084
rect 177868 635020 177869 635084
rect 177803 635019 177869 635020
rect 177806 624613 177866 635019
rect 178910 628965 178970 636923
rect 179094 632229 179154 641683
rect 179091 632228 179157 632229
rect 179091 632164 179092 632228
rect 179156 632164 179157 632228
rect 179091 632163 179157 632164
rect 179278 630053 179338 643179
rect 181794 633097 182414 650898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 633097 186134 654618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 633097 189854 658338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 633097 193574 662058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 633097 197294 665778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 633097 201014 633498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 633097 204734 637218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 633097 208454 640938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 633097 218414 650898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 633097 222134 654618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 633097 225854 658338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 633097 229574 662058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 633097 233294 665778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 633097 237014 633498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 633097 240734 637218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 633097 244454 640938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 633097 254414 650898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 179275 630052 179341 630053
rect 179275 629988 179276 630052
rect 179340 629988 179341 630052
rect 179275 629987 179341 629988
rect 178907 628964 178973 628965
rect 178907 628900 178908 628964
rect 178972 628900 178973 628964
rect 178907 628899 178973 628900
rect 177803 624612 177869 624613
rect 177803 624548 177804 624612
rect 177868 624548 177869 624612
rect 177803 624547 177869 624548
rect 177803 622436 177869 622437
rect 177803 622372 177804 622436
rect 177868 622372 177869 622436
rect 177803 622371 177869 622372
rect 177619 619172 177685 619173
rect 177619 619108 177620 619172
rect 177684 619108 177685 619172
rect 177619 619107 177685 619108
rect 177435 618084 177501 618085
rect 177435 618020 177436 618084
rect 177500 618020 177501 618084
rect 177435 618019 177501 618020
rect 177067 615908 177133 615909
rect 177067 615844 177068 615908
rect 177132 615844 177133 615908
rect 177067 615843 177133 615844
rect 173939 615364 174005 615365
rect 173939 615300 173940 615364
rect 174004 615300 174005 615364
rect 173939 615299 174005 615300
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171547 570212 171613 570213
rect 171547 570148 171548 570212
rect 171612 570148 171613 570212
rect 171547 570147 171613 570148
rect 170995 553212 171061 553213
rect 170995 553148 170996 553212
rect 171060 553148 171061 553212
rect 170995 553147 171061 553148
rect 170259 547772 170325 547773
rect 170259 547708 170260 547772
rect 170324 547708 170325 547772
rect 170259 547707 170325 547708
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 519809 168734 529218
rect 171550 526149 171610 570147
rect 171834 569494 172454 604938
rect 173755 603940 173821 603941
rect 173755 603876 173756 603940
rect 173820 603876 173821 603940
rect 173755 603875 173821 603876
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171834 533494 172454 568938
rect 173571 568036 173637 568037
rect 173571 567972 173572 568036
rect 173636 567972 173637 568036
rect 173571 567971 173637 567972
rect 173574 553213 173634 567971
rect 173758 558109 173818 603875
rect 173942 560285 174002 615299
rect 175779 612100 175845 612101
rect 175779 612036 175780 612100
rect 175844 612036 175845 612100
rect 175779 612035 175845 612036
rect 174859 565860 174925 565861
rect 174859 565796 174860 565860
rect 174924 565796 174925 565860
rect 174859 565795 174925 565796
rect 173939 560284 174005 560285
rect 173939 560220 173940 560284
rect 174004 560220 174005 560284
rect 173939 560219 174005 560220
rect 173755 558108 173821 558109
rect 173755 558044 173756 558108
rect 173820 558044 173821 558108
rect 173755 558043 173821 558044
rect 174862 554029 174922 565795
rect 175043 564772 175109 564773
rect 175043 564708 175044 564772
rect 175108 564708 175109 564772
rect 175043 564707 175109 564708
rect 174859 554028 174925 554029
rect 174859 553964 174860 554028
rect 174924 553964 174925 554028
rect 174859 553963 174925 553964
rect 173571 553212 173637 553213
rect 173571 553148 173572 553212
rect 173636 553148 173637 553212
rect 173571 553147 173637 553148
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171547 526148 171613 526149
rect 171547 526084 171548 526148
rect 171612 526084 171613 526148
rect 171547 526083 171613 526084
rect 171834 519809 172454 532938
rect 175046 525741 175106 564707
rect 175782 527781 175842 612035
rect 177070 610741 177130 615843
rect 177251 611556 177317 611557
rect 177251 611492 177252 611556
rect 177316 611492 177317 611556
rect 177251 611491 177317 611492
rect 177067 610740 177133 610741
rect 177067 610676 177068 610740
rect 177132 610676 177133 610740
rect 177067 610675 177133 610676
rect 176883 607204 176949 607205
rect 176883 607140 176884 607204
rect 176948 607140 176949 607204
rect 176883 607139 176949 607140
rect 175963 604756 176029 604757
rect 175963 604692 175964 604756
rect 176028 604692 176029 604756
rect 175963 604691 176029 604692
rect 175966 543013 176026 604691
rect 176886 554709 176946 607139
rect 177254 607069 177314 611491
rect 177438 611421 177498 618019
rect 177619 616996 177685 616997
rect 177619 616932 177620 616996
rect 177684 616932 177685 616996
rect 177619 616931 177685 616932
rect 177622 611693 177682 616931
rect 177806 612781 177866 622371
rect 199568 619174 199888 619206
rect 199568 618938 199610 619174
rect 199846 618938 199888 619174
rect 199568 618854 199888 618938
rect 199568 618618 199610 618854
rect 199846 618618 199888 618854
rect 199568 618586 199888 618618
rect 230288 619174 230608 619206
rect 230288 618938 230330 619174
rect 230566 618938 230608 619174
rect 230288 618854 230608 618938
rect 230288 618618 230330 618854
rect 230566 618618 230608 618854
rect 230288 618586 230608 618618
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 184208 615454 184528 615486
rect 184208 615218 184250 615454
rect 184486 615218 184528 615454
rect 184208 615134 184528 615218
rect 184208 614898 184250 615134
rect 184486 614898 184528 615134
rect 184208 614866 184528 614898
rect 214928 615454 215248 615486
rect 214928 615218 214970 615454
rect 215206 615218 215248 615454
rect 214928 615134 215248 615218
rect 214928 614898 214970 615134
rect 215206 614898 215248 615134
rect 214928 614866 215248 614898
rect 245648 615454 245968 615486
rect 245648 615218 245690 615454
rect 245926 615218 245968 615454
rect 245648 615134 245968 615218
rect 245648 614898 245690 615134
rect 245926 614898 245968 615134
rect 245648 614866 245968 614898
rect 177987 613732 178053 613733
rect 177987 613668 177988 613732
rect 178052 613668 178053 613732
rect 177987 613667 178053 613668
rect 177803 612780 177869 612781
rect 177803 612716 177804 612780
rect 177868 612716 177869 612780
rect 177803 612715 177869 612716
rect 177803 612644 177869 612645
rect 177803 612580 177804 612644
rect 177868 612580 177869 612644
rect 177803 612579 177869 612580
rect 177619 611692 177685 611693
rect 177619 611628 177620 611692
rect 177684 611628 177685 611692
rect 177619 611627 177685 611628
rect 177435 611420 177501 611421
rect 177435 611356 177436 611420
rect 177500 611356 177501 611420
rect 177435 611355 177501 611356
rect 177619 610468 177685 610469
rect 177619 610404 177620 610468
rect 177684 610404 177685 610468
rect 177619 610403 177685 610404
rect 177251 607068 177317 607069
rect 177251 607004 177252 607068
rect 177316 607004 177317 607068
rect 177251 607003 177317 607004
rect 177435 605844 177501 605845
rect 177435 605780 177436 605844
rect 177500 605780 177501 605844
rect 177435 605779 177501 605780
rect 177067 605028 177133 605029
rect 177067 604964 177068 605028
rect 177132 604964 177133 605028
rect 177067 604963 177133 604964
rect 176883 554708 176949 554709
rect 176883 554644 176884 554708
rect 176948 554644 176949 554708
rect 176883 554643 176949 554644
rect 175963 543012 176029 543013
rect 175963 542948 175964 543012
rect 176028 542948 176029 543012
rect 175963 542947 176029 542948
rect 177070 529413 177130 604963
rect 177438 600810 177498 605779
rect 177622 604485 177682 610403
rect 177806 609650 177866 612579
rect 177990 609789 178050 613667
rect 178171 613596 178237 613597
rect 178171 613532 178172 613596
rect 178236 613532 178237 613596
rect 178171 613531 178237 613532
rect 177987 609788 178053 609789
rect 177987 609724 177988 609788
rect 178052 609724 178053 609788
rect 177987 609723 178053 609724
rect 177806 609590 178050 609650
rect 177803 609380 177869 609381
rect 177803 609316 177804 609380
rect 177868 609316 177869 609380
rect 177803 609315 177869 609316
rect 177619 604484 177685 604485
rect 177619 604420 177620 604484
rect 177684 604420 177685 604484
rect 177619 604419 177685 604420
rect 177619 602852 177685 602853
rect 177619 602788 177620 602852
rect 177684 602788 177685 602852
rect 177619 602787 177685 602788
rect 177254 600750 177498 600810
rect 177254 569941 177314 600750
rect 177622 586530 177682 602787
rect 177806 601765 177866 609315
rect 177990 607069 178050 609590
rect 177987 607068 178053 607069
rect 177987 607004 177988 607068
rect 178052 607004 178053 607068
rect 177987 607003 178053 607004
rect 178174 605850 178234 613531
rect 177990 605790 178234 605850
rect 177803 601764 177869 601765
rect 177803 601700 177804 601764
rect 177868 601700 177869 601764
rect 177803 601699 177869 601700
rect 177438 586470 177682 586530
rect 177251 569940 177317 569941
rect 177251 569876 177252 569940
rect 177316 569876 177317 569940
rect 177251 569875 177317 569876
rect 177438 555253 177498 586470
rect 177803 569124 177869 569125
rect 177803 569060 177804 569124
rect 177868 569060 177869 569124
rect 177803 569059 177869 569060
rect 177806 555389 177866 569059
rect 177990 560285 178050 605790
rect 255819 602852 255885 602853
rect 255819 602788 255820 602852
rect 255884 602788 255885 602852
rect 255819 602787 255885 602788
rect 199568 583174 199888 583206
rect 199568 582938 199610 583174
rect 199846 582938 199888 583174
rect 199568 582854 199888 582938
rect 199568 582618 199610 582854
rect 199846 582618 199888 582854
rect 199568 582586 199888 582618
rect 230288 583174 230608 583206
rect 230288 582938 230330 583174
rect 230566 582938 230608 583174
rect 230288 582854 230608 582938
rect 230288 582618 230330 582854
rect 230566 582618 230608 582854
rect 230288 582586 230608 582618
rect 184208 579454 184528 579486
rect 184208 579218 184250 579454
rect 184486 579218 184528 579454
rect 184208 579134 184528 579218
rect 184208 578898 184250 579134
rect 184486 578898 184528 579134
rect 184208 578866 184528 578898
rect 214928 579454 215248 579486
rect 214928 579218 214970 579454
rect 215206 579218 215248 579454
rect 214928 579134 215248 579218
rect 214928 578898 214970 579134
rect 215206 578898 215248 579134
rect 214928 578866 215248 578898
rect 245648 579454 245968 579486
rect 245648 579218 245690 579454
rect 245926 579218 245968 579454
rect 245648 579134 245968 579218
rect 245648 578898 245690 579134
rect 245926 578898 245968 579134
rect 245648 578866 245968 578898
rect 179275 566948 179341 566949
rect 179275 566884 179276 566948
rect 179340 566884 179341 566948
rect 179275 566883 179341 566884
rect 179091 563548 179157 563549
rect 179091 563484 179092 563548
rect 179156 563484 179157 563548
rect 179091 563483 179157 563484
rect 177987 560284 178053 560285
rect 177987 560220 177988 560284
rect 178052 560220 178053 560284
rect 177987 560219 178053 560220
rect 179094 558245 179154 563483
rect 179278 562189 179338 566883
rect 180563 562528 180629 562529
rect 180563 562464 180564 562528
rect 180628 562464 180629 562528
rect 180563 562463 180629 562464
rect 179275 562188 179341 562189
rect 179275 562124 179276 562188
rect 179340 562124 179341 562188
rect 179275 562123 179341 562124
rect 179827 561440 179893 561441
rect 179827 561376 179828 561440
rect 179892 561376 179893 561440
rect 179827 561375 179893 561376
rect 179091 558244 179157 558245
rect 179091 558180 179092 558244
rect 179156 558180 179157 558244
rect 179091 558179 179157 558180
rect 177803 555388 177869 555389
rect 177803 555324 177804 555388
rect 177868 555324 177869 555388
rect 177803 555323 177869 555324
rect 177435 555252 177501 555253
rect 177435 555188 177436 555252
rect 177500 555188 177501 555252
rect 177435 555187 177501 555188
rect 177067 529412 177133 529413
rect 177067 529348 177068 529412
rect 177132 529348 177133 529412
rect 177067 529347 177133 529348
rect 175779 527780 175845 527781
rect 175779 527716 175780 527780
rect 175844 527716 175845 527780
rect 175779 527715 175845 527716
rect 179830 525741 179890 561375
rect 180566 558381 180626 562463
rect 180563 558380 180629 558381
rect 180563 558316 180564 558380
rect 180628 558316 180629 558380
rect 180563 558315 180629 558316
rect 196674 558334 197294 558575
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 175043 525740 175109 525741
rect 175043 525676 175044 525740
rect 175108 525676 175109 525740
rect 175043 525675 175109 525676
rect 179827 525740 179893 525741
rect 179827 525676 179828 525740
rect 179892 525676 179893 525740
rect 179827 525675 179893 525676
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 519809 197294 521778
rect 232674 558334 233294 558575
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522334 233294 557778
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 232674 519809 233294 521778
rect 255822 519621 255882 602787
rect 256739 599860 256805 599861
rect 256739 599796 256740 599860
rect 256804 599796 256805 599860
rect 256739 599795 256805 599796
rect 256742 594829 256802 599795
rect 256923 596596 256989 596597
rect 256923 596532 256924 596596
rect 256988 596532 256989 596596
rect 256923 596531 256989 596532
rect 256739 594828 256805 594829
rect 256739 594764 256740 594828
rect 256804 594764 256805 594828
rect 256739 594763 256805 594764
rect 256739 575380 256805 575381
rect 256739 575316 256740 575380
rect 256804 575316 256805 575380
rect 256739 575315 256805 575316
rect 256742 547637 256802 575315
rect 256926 574157 256986 596531
rect 257107 595780 257173 595781
rect 257107 595716 257108 595780
rect 257172 595716 257173 595780
rect 257107 595715 257173 595716
rect 256923 574156 256989 574157
rect 256923 574092 256924 574156
rect 256988 574092 256989 574156
rect 256923 574091 256989 574092
rect 256739 547636 256805 547637
rect 256739 547572 256740 547636
rect 256804 547572 256805 547636
rect 256739 547571 256805 547572
rect 257110 522885 257170 595715
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257107 522884 257173 522885
rect 257107 522820 257108 522884
rect 257172 522820 257173 522884
rect 257107 522819 257173 522820
rect 257514 519809 258134 546618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 262811 603940 262877 603941
rect 262811 603876 262812 603940
rect 262876 603876 262877 603940
rect 262811 603875 262877 603876
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 262814 552941 262874 603875
rect 264954 590614 265574 626058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 265939 603124 266005 603125
rect 265939 603060 265940 603124
rect 266004 603060 266005 603124
rect 265939 603059 266005 603060
rect 265755 590884 265821 590885
rect 265755 590820 265756 590884
rect 265820 590820 265821 590884
rect 265755 590819 265821 590820
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 262811 552940 262877 552941
rect 262811 552876 262812 552940
rect 262876 552876 262877 552940
rect 262811 552875 262877 552876
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 519809 261854 550338
rect 264954 519809 265574 554058
rect 265758 519621 265818 590819
rect 265942 557157 266002 603059
rect 266859 601492 266925 601493
rect 266859 601428 266860 601492
rect 266924 601428 266925 601492
rect 266859 601427 266925 601428
rect 265939 557156 266005 557157
rect 265939 557092 265940 557156
rect 266004 557092 266005 557156
rect 265939 557091 266005 557092
rect 266862 532405 266922 601427
rect 268147 594964 268213 594965
rect 268147 594900 268148 594964
rect 268212 594900 268213 594964
rect 268147 594899 268213 594900
rect 268150 559333 268210 594899
rect 268674 594334 269294 629778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 271091 613596 271157 613597
rect 271091 613532 271092 613596
rect 271156 613532 271157 613596
rect 271091 613531 271157 613532
rect 269803 604756 269869 604757
rect 269803 604692 269804 604756
rect 269868 604692 269869 604756
rect 269803 604691 269869 604692
rect 268674 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 269294 594334
rect 268674 594014 269294 594098
rect 269619 594148 269685 594149
rect 269619 594084 269620 594148
rect 269684 594084 269685 594148
rect 269619 594083 269685 594084
rect 268674 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 269294 594014
rect 268331 589252 268397 589253
rect 268331 589188 268332 589252
rect 268396 589188 268397 589252
rect 268331 589187 268397 589188
rect 268147 559332 268213 559333
rect 268147 559268 268148 559332
rect 268212 559268 268213 559332
rect 268147 559267 268213 559268
rect 266859 532404 266925 532405
rect 266859 532340 266860 532404
rect 266924 532340 266925 532404
rect 266859 532339 266925 532340
rect 255819 519620 255885 519621
rect 255819 519556 255820 519620
rect 255884 519556 255885 519620
rect 255819 519555 255885 519556
rect 265755 519620 265821 519621
rect 265755 519556 265756 519620
rect 265820 519556 265821 519620
rect 265755 519555 265821 519556
rect 268334 518533 268394 589187
rect 268674 558334 269294 593778
rect 268674 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 269294 558334
rect 268674 558014 269294 558098
rect 268674 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 269294 558014
rect 268674 522334 269294 557778
rect 268674 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 269294 522334
rect 268674 522014 269294 522098
rect 268674 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 269294 522014
rect 268674 519809 269294 521778
rect 269622 518941 269682 594083
rect 269806 551037 269866 604691
rect 269803 551036 269869 551037
rect 269803 550972 269804 551036
rect 269868 550972 269869 551036
rect 269803 550971 269869 550972
rect 269619 518940 269685 518941
rect 269619 518876 269620 518940
rect 269684 518876 269685 518940
rect 269619 518875 269685 518876
rect 271094 518669 271154 613531
rect 271275 607068 271341 607069
rect 271275 607004 271276 607068
rect 271340 607004 271341 607068
rect 271275 607003 271341 607004
rect 271278 550357 271338 607003
rect 272011 606388 272077 606389
rect 272011 606324 272012 606388
rect 272076 606324 272077 606388
rect 272011 606323 272077 606324
rect 271459 582724 271525 582725
rect 271459 582660 271460 582724
rect 271524 582660 271525 582724
rect 271459 582659 271525 582660
rect 271275 550356 271341 550357
rect 271275 550292 271276 550356
rect 271340 550292 271341 550356
rect 271275 550291 271341 550292
rect 271462 547501 271522 582659
rect 271459 547500 271525 547501
rect 271459 547436 271460 547500
rect 271524 547436 271525 547500
rect 271459 547435 271525 547436
rect 272014 540157 272074 606323
rect 272394 598054 273014 633498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 273851 617132 273917 617133
rect 273851 617068 273852 617132
rect 273916 617068 273917 617132
rect 273851 617067 273917 617068
rect 272394 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 273014 598054
rect 272394 597734 273014 597818
rect 272394 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 273014 597734
rect 272394 562054 273014 597498
rect 272394 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 273014 562054
rect 272394 561734 273014 561818
rect 272394 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 273014 561734
rect 272011 540156 272077 540157
rect 272011 540092 272012 540156
rect 272076 540092 272077 540156
rect 272011 540091 272077 540092
rect 272394 526054 273014 561498
rect 273854 548861 273914 617067
rect 276114 601774 276734 637218
rect 276114 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 276734 601774
rect 276114 601454 276734 601538
rect 276114 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 276734 601454
rect 275139 598228 275205 598229
rect 275139 598164 275140 598228
rect 275204 598164 275205 598228
rect 275139 598163 275205 598164
rect 274035 581092 274101 581093
rect 274035 581028 274036 581092
rect 274100 581028 274101 581092
rect 274035 581027 274101 581028
rect 274038 548861 274098 581027
rect 275142 555117 275202 598163
rect 276114 565774 276734 601218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 605494 280454 640938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 282867 636988 282933 636989
rect 282867 636924 282868 636988
rect 282932 636924 282933 636988
rect 282867 636923 282933 636924
rect 282131 623524 282197 623525
rect 282131 623460 282132 623524
rect 282196 623460 282197 623524
rect 282131 623459 282197 623460
rect 279834 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 280454 605494
rect 279834 605174 280454 605258
rect 279834 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 280454 605174
rect 277899 600676 277965 600677
rect 277899 600612 277900 600676
rect 277964 600612 277965 600676
rect 277899 600611 277965 600612
rect 277163 588436 277229 588437
rect 277163 588372 277164 588436
rect 277228 588372 277229 588436
rect 277163 588371 277229 588372
rect 277166 567210 277226 588371
rect 276114 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 276734 565774
rect 276114 565454 276734 565538
rect 276114 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 276734 565454
rect 275139 555116 275205 555117
rect 275139 555052 275140 555116
rect 275204 555052 275205 555116
rect 275139 555051 275205 555052
rect 273851 548860 273917 548861
rect 273851 548796 273852 548860
rect 273916 548796 273917 548860
rect 273851 548795 273917 548796
rect 274035 548860 274101 548861
rect 274035 548796 274036 548860
rect 274100 548796 274101 548860
rect 274035 548795 274101 548796
rect 272394 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 273014 526054
rect 272394 525734 273014 525818
rect 272394 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 273014 525734
rect 272394 519809 273014 525498
rect 276114 529774 276734 565218
rect 276982 567150 277226 567210
rect 276982 560829 277042 567150
rect 277163 565860 277229 565861
rect 277163 565796 277164 565860
rect 277228 565796 277229 565860
rect 277163 565795 277229 565796
rect 276979 560828 277045 560829
rect 276979 560764 276980 560828
rect 277044 560764 277045 560828
rect 276979 560763 277045 560764
rect 277166 560690 277226 565795
rect 276982 560630 277226 560690
rect 276982 535261 277042 560630
rect 277163 560420 277229 560421
rect 277163 560356 277164 560420
rect 277228 560356 277229 560420
rect 277163 560355 277229 560356
rect 277166 544373 277226 560355
rect 277902 559877 277962 600611
rect 279834 569494 280454 604938
rect 280659 603940 280725 603941
rect 280659 603876 280660 603940
rect 280724 603876 280725 603940
rect 280659 603875 280725 603876
rect 279834 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 280454 569494
rect 279834 569174 280454 569258
rect 279834 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 280454 569174
rect 279371 564772 279437 564773
rect 279371 564708 279372 564772
rect 279436 564708 279437 564772
rect 279371 564707 279437 564708
rect 277899 559876 277965 559877
rect 277899 559812 277900 559876
rect 277964 559812 277965 559876
rect 277899 559811 277965 559812
rect 277163 544372 277229 544373
rect 277163 544308 277164 544372
rect 277228 544308 277229 544372
rect 277163 544307 277229 544308
rect 276979 535260 277045 535261
rect 276979 535196 276980 535260
rect 277044 535196 277045 535260
rect 276979 535195 277045 535196
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 276114 519809 276734 529218
rect 279374 521117 279434 564707
rect 279834 533494 280454 568938
rect 279834 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 280454 533494
rect 279834 533174 280454 533258
rect 279834 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 280454 533174
rect 279371 521116 279437 521117
rect 279371 521052 279372 521116
rect 279436 521052 279437 521116
rect 279371 521051 279437 521052
rect 279834 519809 280454 532938
rect 280662 522341 280722 603875
rect 280843 602308 280909 602309
rect 280843 602244 280844 602308
rect 280908 602244 280909 602308
rect 280843 602243 280909 602244
rect 280846 558925 280906 602243
rect 281027 570212 281093 570213
rect 281027 570148 281028 570212
rect 281092 570148 281093 570212
rect 281027 570147 281093 570148
rect 280843 558924 280909 558925
rect 280843 558860 280844 558924
rect 280908 558860 280909 558924
rect 280843 558859 280909 558860
rect 280843 558108 280909 558109
rect 280843 558044 280844 558108
rect 280908 558044 280909 558108
rect 280843 558043 280909 558044
rect 280846 523701 280906 558043
rect 281030 540565 281090 570147
rect 281395 558924 281461 558925
rect 281395 558860 281396 558924
rect 281460 558860 281461 558924
rect 281395 558859 281461 558860
rect 281398 557837 281458 558859
rect 281395 557836 281461 557837
rect 281395 557772 281396 557836
rect 281460 557772 281461 557836
rect 281395 557771 281461 557772
rect 281027 540564 281093 540565
rect 281027 540500 281028 540564
rect 281092 540500 281093 540564
rect 281027 540499 281093 540500
rect 282134 531317 282194 623459
rect 282870 563070 282930 636923
rect 288387 625972 288453 625973
rect 288387 625908 288388 625972
rect 288452 625908 288453 625972
rect 288387 625907 288453 625908
rect 286179 625156 286245 625157
rect 286179 625092 286180 625156
rect 286244 625092 286245 625156
rect 286179 625091 286245 625092
rect 283419 624340 283485 624341
rect 283419 624276 283420 624340
rect 283484 624276 283485 624340
rect 283419 624275 283485 624276
rect 282686 563010 282930 563070
rect 282686 559061 282746 563010
rect 282683 559060 282749 559061
rect 282683 558996 282684 559060
rect 282748 558996 282749 559060
rect 282683 558995 282749 558996
rect 283422 533221 283482 624275
rect 285627 622708 285693 622709
rect 285627 622644 285628 622708
rect 285692 622644 285693 622708
rect 285627 622643 285693 622644
rect 284891 587620 284957 587621
rect 284891 587556 284892 587620
rect 284956 587556 284957 587620
rect 284891 587555 284957 587556
rect 283603 583540 283669 583541
rect 283603 583476 283604 583540
rect 283668 583476 283669 583540
rect 283603 583475 283669 583476
rect 283419 533220 283485 533221
rect 283419 533156 283420 533220
rect 283484 533156 283485 533220
rect 283419 533155 283485 533156
rect 282131 531316 282197 531317
rect 282131 531252 282132 531316
rect 282196 531252 282197 531316
rect 282131 531251 282197 531252
rect 280843 523700 280909 523701
rect 280843 523636 280844 523700
rect 280908 523636 280909 523700
rect 280843 523635 280909 523636
rect 280659 522340 280725 522341
rect 280659 522276 280660 522340
rect 280724 522276 280725 522340
rect 280659 522275 280725 522276
rect 283606 520029 283666 583475
rect 283603 520028 283669 520029
rect 283603 519964 283604 520028
rect 283668 519964 283669 520028
rect 283603 519963 283669 519964
rect 284894 519213 284954 587555
rect 285259 566948 285325 566949
rect 285259 566884 285260 566948
rect 285324 566884 285325 566948
rect 285259 566883 285325 566884
rect 285075 563684 285141 563685
rect 285075 563620 285076 563684
rect 285140 563620 285141 563684
rect 285075 563619 285141 563620
rect 285078 519485 285138 563619
rect 285262 535125 285322 566883
rect 285259 535124 285325 535125
rect 285259 535060 285260 535124
rect 285324 535060 285325 535124
rect 285259 535059 285325 535060
rect 285630 527645 285690 622643
rect 285811 621076 285877 621077
rect 285811 621012 285812 621076
rect 285876 621012 285877 621076
rect 285811 621011 285877 621012
rect 285814 583813 285874 621011
rect 285811 583812 285877 583813
rect 285811 583748 285812 583812
rect 285876 583748 285877 583812
rect 285811 583747 285877 583748
rect 286182 531861 286242 625091
rect 286363 611556 286429 611557
rect 286363 611492 286364 611556
rect 286428 611492 286429 611556
rect 286363 611491 286429 611492
rect 286366 546141 286426 611491
rect 286547 584356 286613 584357
rect 286547 584292 286548 584356
rect 286612 584292 286613 584356
rect 286547 584291 286613 584292
rect 286550 550357 286610 584291
rect 287835 562596 287901 562597
rect 287835 562532 287836 562596
rect 287900 562532 287901 562596
rect 287835 562531 287901 562532
rect 286547 550356 286613 550357
rect 286547 550292 286548 550356
rect 286612 550292 286613 550356
rect 286547 550291 286613 550292
rect 286363 546140 286429 546141
rect 286363 546076 286364 546140
rect 286428 546076 286429 546140
rect 286363 546075 286429 546076
rect 286179 531860 286245 531861
rect 286179 531796 286180 531860
rect 286244 531796 286245 531860
rect 286179 531795 286245 531796
rect 285627 527644 285693 527645
rect 285627 527580 285628 527644
rect 285692 527580 285693 527644
rect 285627 527579 285693 527580
rect 287838 520981 287898 562531
rect 288390 529413 288450 625907
rect 288571 621892 288637 621893
rect 288571 621828 288572 621892
rect 288636 621828 288637 621892
rect 288571 621827 288637 621828
rect 288574 530501 288634 621827
rect 289794 615454 290414 650898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 291147 619444 291213 619445
rect 291147 619380 291148 619444
rect 291212 619380 291213 619444
rect 291147 619379 291213 619380
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289123 585172 289189 585173
rect 289123 585108 289124 585172
rect 289188 585108 289189 585172
rect 289123 585107 289189 585108
rect 288939 568852 289005 568853
rect 288939 568788 288940 568852
rect 289004 568788 289005 568852
rect 288939 568787 289005 568788
rect 288571 530500 288637 530501
rect 288571 530436 288572 530500
rect 288636 530436 288637 530500
rect 288571 530435 288637 530436
rect 288387 529412 288453 529413
rect 288387 529348 288388 529412
rect 288452 529348 288453 529412
rect 288387 529347 288453 529348
rect 288942 526013 289002 568787
rect 289126 545597 289186 585107
rect 289794 579454 290414 614898
rect 290595 581908 290661 581909
rect 290595 581844 290596 581908
rect 290660 581844 290661 581908
rect 290595 581843 290661 581844
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289123 545596 289189 545597
rect 289123 545532 289124 545596
rect 289188 545532 289189 545596
rect 289123 545531 289189 545532
rect 289794 543454 290414 578898
rect 290598 578237 290658 581843
rect 290963 579460 291029 579461
rect 290963 579396 290964 579460
rect 291028 579396 291029 579460
rect 290963 579395 291029 579396
rect 290595 578236 290661 578237
rect 290595 578172 290596 578236
rect 290660 578172 290661 578236
rect 290595 578171 290661 578172
rect 290779 577012 290845 577013
rect 290779 576948 290780 577012
rect 290844 576948 290845 577012
rect 290779 576947 290845 576948
rect 290782 554301 290842 576947
rect 290779 554300 290845 554301
rect 290779 554236 290780 554300
rect 290844 554236 290845 554300
rect 290779 554235 290845 554236
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 288939 526012 289005 526013
rect 288939 525948 288940 526012
rect 289004 525948 289005 526012
rect 288939 525947 289005 525948
rect 287835 520980 287901 520981
rect 287835 520916 287836 520980
rect 287900 520916 287901 520980
rect 287835 520915 287901 520916
rect 289794 519809 290414 542898
rect 290966 519485 291026 579395
rect 291150 578237 291210 619379
rect 293514 619174 294134 654618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 296483 644740 296549 644741
rect 296483 644676 296484 644740
rect 296548 644676 296549 644740
rect 296483 644675 296549 644676
rect 296486 635490 296546 644675
rect 296851 642292 296917 642293
rect 296851 642228 296852 642292
rect 296916 642228 296917 642292
rect 296851 642227 296917 642228
rect 296486 635430 296730 635490
rect 296670 634813 296730 635430
rect 296483 634812 296549 634813
rect 296483 634748 296484 634812
rect 296548 634748 296549 634812
rect 296483 634747 296549 634748
rect 296667 634812 296733 634813
rect 296667 634748 296668 634812
rect 296732 634748 296733 634812
rect 296667 634747 296733 634748
rect 296486 621757 296546 634747
rect 296854 623525 296914 642227
rect 296851 623524 296917 623525
rect 296851 623460 296852 623524
rect 296916 623460 296917 623524
rect 296851 623459 296917 623460
rect 297234 622894 297854 658338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 633097 301574 662058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 633097 305294 665778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 633097 309014 633498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 312114 633097 312734 637218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 633097 316454 640938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 633097 326414 650898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 633097 330134 654618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 633097 333854 658338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 633097 337574 662058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 633097 341294 665778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 633097 345014 633498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 633097 348734 637218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 633097 352454 640938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 633097 362414 650898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 634540 366134 654618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 633097 369854 658338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 633097 373574 662058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 375419 644332 375485 644333
rect 375419 644268 375420 644332
rect 375484 644268 375485 644332
rect 375419 644267 375485 644268
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 296483 621756 296549 621757
rect 296483 621692 296484 621756
rect 296548 621692 296549 621756
rect 296483 621691 296549 621692
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 291331 618628 291397 618629
rect 291331 618564 291332 618628
rect 291396 618564 291397 618628
rect 291331 618563 291397 618564
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 291334 579597 291394 618563
rect 292803 616996 292869 616997
rect 292803 616932 292804 616996
rect 292868 616932 292869 616996
rect 292803 616931 292869 616932
rect 292619 616180 292685 616181
rect 292619 616116 292620 616180
rect 292684 616116 292685 616180
rect 292619 616115 292685 616116
rect 291515 586804 291581 586805
rect 291515 586740 291516 586804
rect 291580 586740 291581 586804
rect 291515 586739 291581 586740
rect 291331 579596 291397 579597
rect 291331 579532 291332 579596
rect 291396 579532 291397 579596
rect 291331 579531 291397 579532
rect 291147 578236 291213 578237
rect 291147 578172 291148 578236
rect 291212 578172 291213 578236
rect 291147 578171 291213 578172
rect 291518 572933 291578 586739
rect 292251 580276 292317 580277
rect 292251 580212 292252 580276
rect 292316 580212 292317 580276
rect 292251 580211 292317 580212
rect 291883 578644 291949 578645
rect 291883 578580 291884 578644
rect 291948 578580 291949 578644
rect 291883 578579 291949 578580
rect 291699 577692 291765 577693
rect 291699 577628 291700 577692
rect 291764 577628 291765 577692
rect 291699 577627 291765 577628
rect 291515 572932 291581 572933
rect 291515 572868 291516 572932
rect 291580 572868 291581 572932
rect 291515 572867 291581 572868
rect 285075 519484 285141 519485
rect 285075 519420 285076 519484
rect 285140 519420 285141 519484
rect 285075 519419 285141 519420
rect 290963 519484 291029 519485
rect 290963 519420 290964 519484
rect 291028 519420 291029 519484
rect 290963 519419 291029 519420
rect 291702 519349 291762 577627
rect 291886 553077 291946 578579
rect 292067 573748 292133 573749
rect 292067 573684 292068 573748
rect 292132 573684 292133 573748
rect 292067 573683 292133 573684
rect 291883 553076 291949 553077
rect 291883 553012 291884 553076
rect 291948 553012 291949 553076
rect 291883 553011 291949 553012
rect 292070 552669 292130 573683
rect 292254 572797 292314 580211
rect 292622 574157 292682 616115
rect 292806 612781 292866 616931
rect 293171 612916 293237 612917
rect 293171 612852 293172 612916
rect 293236 612852 293237 612916
rect 293171 612851 293237 612852
rect 292803 612780 292869 612781
rect 292803 612716 292804 612780
rect 292868 612716 292869 612780
rect 292803 612715 292869 612716
rect 292987 574428 293053 574429
rect 292987 574364 292988 574428
rect 293052 574364 293053 574428
rect 292987 574363 293053 574364
rect 292619 574156 292685 574157
rect 292619 574092 292620 574156
rect 292684 574092 292685 574156
rect 292619 574091 292685 574092
rect 292435 572932 292501 572933
rect 292435 572868 292436 572932
rect 292500 572868 292501 572932
rect 292435 572867 292501 572868
rect 292251 572796 292317 572797
rect 292251 572732 292252 572796
rect 292316 572732 292317 572796
rect 292251 572731 292317 572732
rect 292438 552805 292498 572867
rect 292435 552804 292501 552805
rect 292435 552740 292436 552804
rect 292500 552740 292501 552804
rect 292435 552739 292501 552740
rect 292067 552668 292133 552669
rect 292067 552604 292068 552668
rect 292132 552604 292133 552668
rect 292067 552603 292133 552604
rect 292990 546141 293050 574363
rect 292987 546140 293053 546141
rect 292987 546076 292988 546140
rect 293052 546076 293053 546140
rect 292987 546075 293053 546076
rect 293174 543421 293234 612851
rect 293514 583174 294134 618618
rect 294459 615364 294525 615365
rect 294459 615300 294460 615364
rect 294524 615300 294525 615364
rect 294459 615299 294525 615300
rect 294462 592109 294522 615299
rect 294827 614548 294893 614549
rect 294827 614484 294828 614548
rect 294892 614484 294893 614548
rect 294827 614483 294893 614484
rect 294643 607204 294709 607205
rect 294643 607140 294644 607204
rect 294708 607140 294709 607204
rect 294643 607139 294709 607140
rect 294459 592108 294525 592109
rect 294459 592044 294460 592108
rect 294524 592044 294525 592108
rect 294459 592043 294525 592044
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 294459 572116 294525 572117
rect 294459 572052 294460 572116
rect 294524 572052 294525 572116
rect 294459 572051 294525 572052
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293171 543420 293237 543421
rect 293171 543356 293172 543420
rect 293236 543356 293237 543420
rect 293171 543355 293237 543356
rect 293514 519809 294134 546618
rect 294462 525605 294522 572051
rect 294646 571437 294706 607139
rect 294830 597549 294890 614483
rect 295563 612100 295629 612101
rect 295563 612036 295564 612100
rect 295628 612036 295629 612100
rect 295563 612035 295629 612036
rect 295379 611284 295445 611285
rect 295379 611220 295380 611284
rect 295444 611220 295445 611284
rect 295379 611219 295445 611220
rect 294827 597548 294893 597549
rect 294827 597484 294828 597548
rect 294892 597484 294893 597548
rect 294827 597483 294893 597484
rect 295011 597276 295077 597277
rect 295011 597212 295012 597276
rect 295076 597212 295077 597276
rect 295011 597211 295077 597212
rect 294827 592516 294893 592517
rect 294827 592452 294828 592516
rect 294892 592452 294893 592516
rect 294827 592451 294893 592452
rect 294643 571436 294709 571437
rect 294643 571372 294644 571436
rect 294708 571372 294709 571436
rect 294643 571371 294709 571372
rect 294830 554437 294890 592451
rect 294827 554436 294893 554437
rect 294827 554372 294828 554436
rect 294892 554372 294893 554436
rect 294827 554371 294893 554372
rect 295014 544373 295074 597211
rect 295382 585173 295442 611219
rect 295566 590613 295626 612035
rect 296851 609380 296917 609381
rect 296851 609316 296852 609380
rect 296916 609316 296917 609380
rect 296851 609315 296917 609316
rect 296667 605028 296733 605029
rect 296667 604964 296668 605028
rect 296732 604964 296733 605028
rect 296667 604963 296733 604964
rect 296670 604890 296730 604963
rect 296486 604830 296730 604890
rect 295747 599044 295813 599045
rect 295747 598980 295748 599044
rect 295812 598980 295813 599044
rect 295747 598979 295813 598980
rect 295563 590612 295629 590613
rect 295563 590548 295564 590612
rect 295628 590548 295629 590612
rect 295563 590547 295629 590548
rect 295379 585172 295445 585173
rect 295379 585108 295380 585172
rect 295444 585108 295445 585172
rect 295379 585107 295445 585108
rect 295563 576196 295629 576197
rect 295563 576132 295564 576196
rect 295628 576132 295629 576196
rect 295563 576131 295629 576132
rect 295566 572730 295626 576131
rect 295750 575517 295810 598979
rect 296299 593332 296365 593333
rect 296299 593268 296300 593332
rect 296364 593268 296365 593332
rect 296299 593267 296365 593268
rect 296115 590068 296181 590069
rect 296115 590004 296116 590068
rect 296180 590004 296181 590068
rect 296115 590003 296181 590004
rect 295931 585988 295997 585989
rect 295931 585924 295932 585988
rect 295996 585924 295997 585988
rect 295931 585923 295997 585924
rect 295747 575516 295813 575517
rect 295747 575452 295748 575516
rect 295812 575452 295813 575516
rect 295747 575451 295813 575452
rect 295566 572670 295810 572730
rect 295563 569668 295629 569669
rect 295563 569604 295564 569668
rect 295628 569604 295629 569668
rect 295563 569603 295629 569604
rect 295566 563070 295626 569603
rect 295750 563277 295810 572670
rect 295747 563276 295813 563277
rect 295747 563212 295748 563276
rect 295812 563212 295813 563276
rect 295747 563211 295813 563212
rect 295566 563010 295810 563070
rect 295750 549133 295810 563010
rect 295747 549132 295813 549133
rect 295747 549068 295748 549132
rect 295812 549068 295813 549132
rect 295747 549067 295813 549068
rect 295011 544372 295077 544373
rect 295011 544308 295012 544372
rect 295076 544308 295077 544372
rect 295011 544307 295077 544308
rect 295934 525741 295994 585923
rect 296118 552533 296178 590003
rect 296302 568717 296362 593267
rect 296486 572730 296546 604830
rect 296486 572670 296730 572730
rect 296299 568716 296365 568717
rect 296299 568652 296300 568716
rect 296364 568652 296365 568716
rect 296299 568651 296365 568652
rect 296670 563410 296730 572670
rect 296302 563350 296730 563410
rect 296115 552532 296181 552533
rect 296115 552468 296116 552532
rect 296180 552468 296181 552532
rect 296115 552467 296181 552468
rect 296302 549269 296362 563350
rect 296483 563276 296549 563277
rect 296483 563212 296484 563276
rect 296548 563212 296549 563276
rect 296483 563211 296549 563212
rect 296486 560013 296546 563211
rect 296483 560012 296549 560013
rect 296483 559948 296484 560012
rect 296548 559948 296549 560012
rect 296483 559947 296549 559948
rect 296299 549268 296365 549269
rect 296299 549204 296300 549268
rect 296364 549204 296365 549268
rect 296299 549203 296365 549204
rect 295931 525740 295997 525741
rect 295931 525676 295932 525740
rect 295996 525676 295997 525740
rect 295931 525675 295997 525676
rect 294459 525604 294525 525605
rect 294459 525540 294460 525604
rect 294524 525540 294525 525604
rect 294459 525539 294525 525540
rect 296854 522477 296914 609315
rect 297234 586894 297854 622338
rect 298139 620124 298205 620125
rect 298139 620060 298140 620124
rect 298204 620060 298205 620124
rect 298139 620059 298205 620060
rect 298142 608565 298202 620059
rect 319568 619174 319888 619206
rect 319568 618938 319610 619174
rect 319846 618938 319888 619174
rect 319568 618854 319888 618938
rect 319568 618618 319610 618854
rect 319846 618618 319888 618854
rect 319568 618586 319888 618618
rect 350288 619174 350608 619206
rect 350288 618938 350330 619174
rect 350566 618938 350608 619174
rect 350288 618854 350608 618938
rect 350288 618618 350330 618854
rect 350566 618618 350608 618854
rect 350288 618586 350608 618618
rect 304208 615454 304528 615486
rect 304208 615218 304250 615454
rect 304486 615218 304528 615454
rect 304208 615134 304528 615218
rect 304208 614898 304250 615134
rect 304486 614898 304528 615134
rect 304208 614866 304528 614898
rect 334928 615454 335248 615486
rect 334928 615218 334970 615454
rect 335206 615218 335248 615454
rect 334928 615134 335248 615218
rect 334928 614898 334970 615134
rect 335206 614898 335248 615134
rect 334928 614866 335248 614898
rect 365648 615454 365968 615486
rect 365648 615218 365690 615454
rect 365926 615218 365968 615454
rect 365648 615134 365968 615218
rect 365648 614898 365690 615134
rect 365926 614898 365968 615134
rect 365648 614866 365968 614898
rect 298507 613868 298573 613869
rect 298507 613804 298508 613868
rect 298572 613804 298573 613868
rect 298507 613803 298573 613804
rect 298323 610332 298389 610333
rect 298323 610268 298324 610332
rect 298388 610268 298389 610332
rect 298323 610267 298389 610268
rect 298139 608564 298205 608565
rect 298139 608500 298140 608564
rect 298204 608500 298205 608564
rect 298139 608499 298205 608500
rect 298326 591429 298386 610267
rect 298510 604485 298570 613803
rect 299611 609652 299677 609653
rect 299611 609588 299612 609652
rect 299676 609588 299677 609652
rect 299611 609587 299677 609588
rect 299243 608836 299309 608837
rect 299243 608772 299244 608836
rect 299308 608772 299309 608836
rect 299243 608771 299309 608772
rect 298691 608020 298757 608021
rect 298691 607956 298692 608020
rect 298756 607956 298757 608020
rect 298691 607955 298757 607956
rect 298507 604484 298573 604485
rect 298507 604420 298508 604484
rect 298572 604420 298573 604484
rect 298507 604419 298573 604420
rect 298323 591428 298389 591429
rect 298323 591364 298324 591428
rect 298388 591364 298389 591428
rect 298323 591363 298389 591364
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 296851 522476 296917 522477
rect 296851 522412 296852 522476
rect 296916 522412 296917 522476
rect 296851 522411 296917 522412
rect 297234 519809 297854 550338
rect 298694 522477 298754 607955
rect 299059 605572 299125 605573
rect 299059 605508 299060 605572
rect 299124 605508 299125 605572
rect 299059 605507 299125 605508
rect 298875 591700 298941 591701
rect 298875 591636 298876 591700
rect 298940 591636 298941 591700
rect 298875 591635 298941 591636
rect 298691 522476 298757 522477
rect 298691 522412 298692 522476
rect 298756 522412 298757 522476
rect 298691 522411 298757 522412
rect 291699 519348 291765 519349
rect 291699 519284 291700 519348
rect 291764 519284 291765 519348
rect 291699 519283 291765 519284
rect 284891 519212 284957 519213
rect 284891 519148 284892 519212
rect 284956 519148 284957 519212
rect 284891 519147 284957 519148
rect 298878 518669 298938 591635
rect 299062 548997 299122 605507
rect 299246 570077 299306 608771
rect 299427 570484 299493 570485
rect 299427 570420 299428 570484
rect 299492 570420 299493 570484
rect 299427 570419 299493 570420
rect 299243 570076 299309 570077
rect 299243 570012 299244 570076
rect 299308 570012 299309 570076
rect 299243 570011 299309 570012
rect 299430 563070 299490 570419
rect 299614 570077 299674 609587
rect 375422 608837 375482 644267
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 375419 608836 375485 608837
rect 375419 608772 375420 608836
rect 375484 608772 375485 608836
rect 375419 608771 375485 608772
rect 376674 594334 377294 629778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 377627 602308 377693 602309
rect 377627 602244 377628 602308
rect 377692 602244 377693 602308
rect 377627 602243 377693 602244
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 319568 583174 319888 583206
rect 319568 582938 319610 583174
rect 319846 582938 319888 583174
rect 319568 582854 319888 582938
rect 319568 582618 319610 582854
rect 319846 582618 319888 582854
rect 319568 582586 319888 582618
rect 350288 583174 350608 583206
rect 350288 582938 350330 583174
rect 350566 582938 350608 583174
rect 350288 582854 350608 582938
rect 350288 582618 350330 582854
rect 350566 582618 350608 582854
rect 350288 582586 350608 582618
rect 304208 579454 304528 579486
rect 304208 579218 304250 579454
rect 304486 579218 304528 579454
rect 304208 579134 304528 579218
rect 304208 578898 304250 579134
rect 304486 578898 304528 579134
rect 304208 578866 304528 578898
rect 334928 579454 335248 579486
rect 334928 579218 334970 579454
rect 335206 579218 335248 579454
rect 334928 579134 335248 579218
rect 334928 578898 334970 579134
rect 335206 578898 335248 579134
rect 334928 578866 335248 578898
rect 365648 579454 365968 579486
rect 365648 579218 365690 579454
rect 365926 579218 365968 579454
rect 365648 579134 365968 579218
rect 365648 578898 365690 579134
rect 365926 578898 365968 579134
rect 365648 578866 365968 578898
rect 299795 571164 299861 571165
rect 299795 571100 299796 571164
rect 299860 571100 299861 571164
rect 299795 571099 299861 571100
rect 299611 570076 299677 570077
rect 299611 570012 299612 570076
rect 299676 570012 299677 570076
rect 299611 570011 299677 570012
rect 299246 563010 299490 563070
rect 299059 548996 299125 548997
rect 299059 548932 299060 548996
rect 299124 548932 299125 548996
rect 299059 548931 299125 548932
rect 299246 524925 299306 563010
rect 299798 526285 299858 571099
rect 304674 558334 305294 558575
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 299795 526284 299861 526285
rect 299795 526220 299796 526284
rect 299860 526220 299861 526284
rect 299795 526219 299861 526220
rect 299243 524924 299309 524925
rect 299243 524860 299244 524924
rect 299308 524860 299309 524924
rect 299243 524859 299309 524860
rect 304674 522334 305294 557778
rect 304674 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 305294 522334
rect 304674 522014 305294 522098
rect 304674 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 305294 522014
rect 304674 519809 305294 521778
rect 340674 558334 341294 558575
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522334 341294 557778
rect 340674 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 341294 522334
rect 340674 522014 341294 522098
rect 340674 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 341294 522014
rect 340674 519809 341294 521778
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 377630 529141 377690 602243
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 379467 571300 379533 571301
rect 379467 571236 379468 571300
rect 379532 571236 379533 571300
rect 379467 571235 379533 571236
rect 379470 533357 379530 571235
rect 379651 568852 379717 568853
rect 379651 568788 379652 568852
rect 379716 568788 379717 568852
rect 379651 568787 379717 568788
rect 379654 534853 379714 568787
rect 380394 562054 381014 597498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 381307 577012 381373 577013
rect 381307 576948 381308 577012
rect 381372 576948 381373 577012
rect 381307 576947 381373 576948
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 379651 534852 379717 534853
rect 379651 534788 379652 534852
rect 379716 534788 379717 534852
rect 379651 534787 379717 534788
rect 379835 534172 379901 534173
rect 379835 534108 379836 534172
rect 379900 534108 379901 534172
rect 379835 534107 379901 534108
rect 379467 533356 379533 533357
rect 379467 533292 379468 533356
rect 379532 533292 379533 533356
rect 379467 533291 379533 533292
rect 377627 529140 377693 529141
rect 377627 529076 377628 529140
rect 377692 529076 377693 529140
rect 377627 529075 377693 529076
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 519809 377294 521778
rect 271091 518668 271157 518669
rect 271091 518604 271092 518668
rect 271156 518604 271157 518668
rect 271091 518603 271157 518604
rect 298875 518668 298941 518669
rect 298875 518604 298876 518668
rect 298940 518604 298941 518668
rect 298875 518603 298941 518604
rect 268331 518532 268397 518533
rect 268331 518468 268332 518532
rect 268396 518468 268397 518532
rect 268331 518467 268397 518468
rect 379838 518397 379898 534107
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 519809 381014 525498
rect 379835 518396 379901 518397
rect 379835 518332 379836 518396
rect 379900 518332 379901 518396
rect 379835 518331 379901 518332
rect 381310 518261 381370 576947
rect 383699 572116 383765 572117
rect 383699 572052 383700 572116
rect 383764 572052 383765 572116
rect 383699 572051 383765 572052
rect 382227 570484 382293 570485
rect 382227 570420 382228 570484
rect 382292 570420 382293 570484
rect 382227 570419 382293 570420
rect 382230 536077 382290 570419
rect 382227 536076 382293 536077
rect 382227 536012 382228 536076
rect 382292 536012 382293 536076
rect 382227 536011 382293 536012
rect 383702 534717 383762 572051
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 383699 534716 383765 534717
rect 383699 534652 383700 534716
rect 383764 534652 383765 534716
rect 383699 534651 383765 534652
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 519809 384734 529218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 519809 388454 532938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 519809 398414 542898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 519809 402134 546618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 519809 405854 550338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 519809 409574 554058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 519809 413294 521778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 519809 417014 525498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 519809 420734 529218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 519809 424454 532938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 519809 434414 542898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 519809 438134 546618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 519809 441854 550338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 519809 445574 554058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 519809 449294 521778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 519809 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 519809 456734 529218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 569494 460454 604938
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 519809 460454 532938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 519809 470414 542898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 479563 700364 479629 700365
rect 479563 700300 479564 700364
rect 479628 700300 479629 700364
rect 479563 700299 479629 700300
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 479379 636444 479445 636445
rect 479379 636380 479380 636444
rect 479444 636380 479445 636444
rect 479379 636379 479445 636380
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 476619 560556 476685 560557
rect 476619 560492 476620 560556
rect 476684 560492 476685 560556
rect 476619 560491 476685 560492
rect 474411 559332 474477 559333
rect 474411 559268 474412 559332
rect 474476 559268 474477 559332
rect 474411 559267 474477 559268
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 519809 474134 546618
rect 381307 518260 381373 518261
rect 381307 518196 381308 518260
rect 381372 518196 381373 518260
rect 381307 518195 381373 518196
rect 474414 518125 474474 559267
rect 476067 552940 476133 552941
rect 476067 552876 476068 552940
rect 476132 552876 476133 552940
rect 476067 552875 476133 552876
rect 476070 518805 476130 552875
rect 476067 518804 476133 518805
rect 476067 518740 476068 518804
rect 476132 518740 476133 518804
rect 476067 518739 476133 518740
rect 474411 518124 474477 518125
rect 474411 518060 474412 518124
rect 474476 518060 474477 518124
rect 474411 518059 474477 518060
rect 476622 517989 476682 560491
rect 476803 552532 476869 552533
rect 476803 552468 476804 552532
rect 476868 552468 476869 552532
rect 476803 552467 476869 552468
rect 476806 518397 476866 552467
rect 477234 550894 477854 586338
rect 478091 557156 478157 557157
rect 478091 557092 478092 557156
rect 478156 557092 478157 557156
rect 478091 557091 478157 557092
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 519809 477854 550338
rect 478094 518805 478154 557091
rect 478275 551036 478341 551037
rect 478275 550972 478276 551036
rect 478340 550972 478341 551036
rect 478275 550971 478341 550972
rect 478091 518804 478157 518805
rect 478091 518740 478092 518804
rect 478156 518740 478157 518804
rect 478091 518739 478157 518740
rect 476803 518396 476869 518397
rect 476803 518332 476804 518396
rect 476868 518332 476869 518396
rect 476803 518331 476869 518332
rect 478278 518125 478338 550971
rect 478275 518124 478341 518125
rect 478275 518060 478276 518124
rect 478340 518060 478341 518124
rect 478275 518059 478341 518060
rect 476619 517988 476685 517989
rect 476619 517924 476620 517988
rect 476684 517924 476685 517988
rect 476619 517923 476685 517924
rect 141008 511174 141328 511206
rect 141008 510938 141050 511174
rect 141286 510938 141328 511174
rect 141008 510854 141328 510938
rect 141008 510618 141050 510854
rect 141286 510618 141328 510854
rect 141008 510586 141328 510618
rect 171728 511174 172048 511206
rect 171728 510938 171770 511174
rect 172006 510938 172048 511174
rect 171728 510854 172048 510938
rect 171728 510618 171770 510854
rect 172006 510618 172048 510854
rect 171728 510586 172048 510618
rect 202448 511174 202768 511206
rect 202448 510938 202490 511174
rect 202726 510938 202768 511174
rect 202448 510854 202768 510938
rect 202448 510618 202490 510854
rect 202726 510618 202768 510854
rect 202448 510586 202768 510618
rect 233168 511174 233488 511206
rect 233168 510938 233210 511174
rect 233446 510938 233488 511174
rect 233168 510854 233488 510938
rect 233168 510618 233210 510854
rect 233446 510618 233488 510854
rect 233168 510586 233488 510618
rect 263888 511174 264208 511206
rect 263888 510938 263930 511174
rect 264166 510938 264208 511174
rect 263888 510854 264208 510938
rect 263888 510618 263930 510854
rect 264166 510618 264208 510854
rect 263888 510586 264208 510618
rect 294608 511174 294928 511206
rect 294608 510938 294650 511174
rect 294886 510938 294928 511174
rect 294608 510854 294928 510938
rect 294608 510618 294650 510854
rect 294886 510618 294928 510854
rect 294608 510586 294928 510618
rect 325328 511174 325648 511206
rect 325328 510938 325370 511174
rect 325606 510938 325648 511174
rect 325328 510854 325648 510938
rect 325328 510618 325370 510854
rect 325606 510618 325648 510854
rect 325328 510586 325648 510618
rect 356048 511174 356368 511206
rect 356048 510938 356090 511174
rect 356326 510938 356368 511174
rect 356048 510854 356368 510938
rect 356048 510618 356090 510854
rect 356326 510618 356368 510854
rect 356048 510586 356368 510618
rect 386768 511174 387088 511206
rect 386768 510938 386810 511174
rect 387046 510938 387088 511174
rect 386768 510854 387088 510938
rect 386768 510618 386810 510854
rect 387046 510618 387088 510854
rect 386768 510586 387088 510618
rect 417488 511174 417808 511206
rect 417488 510938 417530 511174
rect 417766 510938 417808 511174
rect 417488 510854 417808 510938
rect 417488 510618 417530 510854
rect 417766 510618 417808 510854
rect 417488 510586 417808 510618
rect 448208 511174 448528 511206
rect 448208 510938 448250 511174
rect 448486 510938 448528 511174
rect 448208 510854 448528 510938
rect 448208 510618 448250 510854
rect 448486 510618 448528 510854
rect 448208 510586 448528 510618
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 309968 507454 310288 507486
rect 309968 507218 310010 507454
rect 310246 507218 310288 507454
rect 309968 507134 310288 507218
rect 309968 506898 310010 507134
rect 310246 506898 310288 507134
rect 309968 506866 310288 506898
rect 340688 507454 341008 507486
rect 340688 507218 340730 507454
rect 340966 507218 341008 507454
rect 340688 507134 341008 507218
rect 340688 506898 340730 507134
rect 340966 506898 341008 507134
rect 340688 506866 341008 506898
rect 371408 507454 371728 507486
rect 371408 507218 371450 507454
rect 371686 507218 371728 507454
rect 371408 507134 371728 507218
rect 371408 506898 371450 507134
rect 371686 506898 371728 507134
rect 371408 506866 371728 506898
rect 402128 507454 402448 507486
rect 402128 507218 402170 507454
rect 402406 507218 402448 507454
rect 402128 507134 402448 507218
rect 402128 506898 402170 507134
rect 402406 506898 402448 507134
rect 402128 506866 402448 506898
rect 432848 507454 433168 507486
rect 432848 507218 432890 507454
rect 433126 507218 433168 507454
rect 432848 507134 433168 507218
rect 432848 506898 432890 507134
rect 433126 506898 433168 507134
rect 432848 506866 433168 506898
rect 463568 507454 463888 507486
rect 463568 507218 463610 507454
rect 463846 507218 463888 507454
rect 463568 507134 463888 507218
rect 463568 506898 463610 507134
rect 463846 506898 463888 507134
rect 463568 506866 463888 506898
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 141008 475174 141328 475206
rect 141008 474938 141050 475174
rect 141286 474938 141328 475174
rect 141008 474854 141328 474938
rect 141008 474618 141050 474854
rect 141286 474618 141328 474854
rect 141008 474586 141328 474618
rect 171728 475174 172048 475206
rect 171728 474938 171770 475174
rect 172006 474938 172048 475174
rect 171728 474854 172048 474938
rect 171728 474618 171770 474854
rect 172006 474618 172048 474854
rect 171728 474586 172048 474618
rect 202448 475174 202768 475206
rect 202448 474938 202490 475174
rect 202726 474938 202768 475174
rect 202448 474854 202768 474938
rect 202448 474618 202490 474854
rect 202726 474618 202768 474854
rect 202448 474586 202768 474618
rect 233168 475174 233488 475206
rect 233168 474938 233210 475174
rect 233446 474938 233488 475174
rect 233168 474854 233488 474938
rect 233168 474618 233210 474854
rect 233446 474618 233488 474854
rect 233168 474586 233488 474618
rect 263888 475174 264208 475206
rect 263888 474938 263930 475174
rect 264166 474938 264208 475174
rect 263888 474854 264208 474938
rect 263888 474618 263930 474854
rect 264166 474618 264208 474854
rect 263888 474586 264208 474618
rect 294608 475174 294928 475206
rect 294608 474938 294650 475174
rect 294886 474938 294928 475174
rect 294608 474854 294928 474938
rect 294608 474618 294650 474854
rect 294886 474618 294928 474854
rect 294608 474586 294928 474618
rect 325328 475174 325648 475206
rect 325328 474938 325370 475174
rect 325606 474938 325648 475174
rect 325328 474854 325648 474938
rect 325328 474618 325370 474854
rect 325606 474618 325648 474854
rect 325328 474586 325648 474618
rect 356048 475174 356368 475206
rect 356048 474938 356090 475174
rect 356326 474938 356368 475174
rect 356048 474854 356368 474938
rect 356048 474618 356090 474854
rect 356326 474618 356368 474854
rect 356048 474586 356368 474618
rect 386768 475174 387088 475206
rect 386768 474938 386810 475174
rect 387046 474938 387088 475174
rect 386768 474854 387088 474938
rect 386768 474618 386810 474854
rect 387046 474618 387088 474854
rect 386768 474586 387088 474618
rect 417488 475174 417808 475206
rect 417488 474938 417530 475174
rect 417766 474938 417808 475174
rect 417488 474854 417808 474938
rect 417488 474618 417530 474854
rect 417766 474618 417808 474854
rect 417488 474586 417808 474618
rect 448208 475174 448528 475206
rect 448208 474938 448250 475174
rect 448486 474938 448528 475174
rect 448208 474854 448528 474938
rect 448208 474618 448250 474854
rect 448486 474618 448528 474854
rect 448208 474586 448528 474618
rect 125648 471454 125968 471486
rect 125648 471218 125690 471454
rect 125926 471218 125968 471454
rect 125648 471134 125968 471218
rect 125648 470898 125690 471134
rect 125926 470898 125968 471134
rect 125648 470866 125968 470898
rect 156368 471454 156688 471486
rect 156368 471218 156410 471454
rect 156646 471218 156688 471454
rect 156368 471134 156688 471218
rect 156368 470898 156410 471134
rect 156646 470898 156688 471134
rect 156368 470866 156688 470898
rect 187088 471454 187408 471486
rect 187088 471218 187130 471454
rect 187366 471218 187408 471454
rect 187088 471134 187408 471218
rect 187088 470898 187130 471134
rect 187366 470898 187408 471134
rect 187088 470866 187408 470898
rect 217808 471454 218128 471486
rect 217808 471218 217850 471454
rect 218086 471218 218128 471454
rect 217808 471134 218128 471218
rect 217808 470898 217850 471134
rect 218086 470898 218128 471134
rect 217808 470866 218128 470898
rect 248528 471454 248848 471486
rect 248528 471218 248570 471454
rect 248806 471218 248848 471454
rect 248528 471134 248848 471218
rect 248528 470898 248570 471134
rect 248806 470898 248848 471134
rect 248528 470866 248848 470898
rect 279248 471454 279568 471486
rect 279248 471218 279290 471454
rect 279526 471218 279568 471454
rect 279248 471134 279568 471218
rect 279248 470898 279290 471134
rect 279526 470898 279568 471134
rect 279248 470866 279568 470898
rect 309968 471454 310288 471486
rect 309968 471218 310010 471454
rect 310246 471218 310288 471454
rect 309968 471134 310288 471218
rect 309968 470898 310010 471134
rect 310246 470898 310288 471134
rect 309968 470866 310288 470898
rect 340688 471454 341008 471486
rect 340688 471218 340730 471454
rect 340966 471218 341008 471454
rect 340688 471134 341008 471218
rect 340688 470898 340730 471134
rect 340966 470898 341008 471134
rect 340688 470866 341008 470898
rect 371408 471454 371728 471486
rect 371408 471218 371450 471454
rect 371686 471218 371728 471454
rect 371408 471134 371728 471218
rect 371408 470898 371450 471134
rect 371686 470898 371728 471134
rect 371408 470866 371728 470898
rect 402128 471454 402448 471486
rect 402128 471218 402170 471454
rect 402406 471218 402448 471454
rect 402128 471134 402448 471218
rect 402128 470898 402170 471134
rect 402406 470898 402448 471134
rect 402128 470866 402448 470898
rect 432848 471454 433168 471486
rect 432848 471218 432890 471454
rect 433126 471218 433168 471454
rect 432848 471134 433168 471218
rect 432848 470898 432890 471134
rect 433126 470898 433168 471134
rect 432848 470866 433168 470898
rect 463568 471454 463888 471486
rect 463568 471218 463610 471454
rect 463846 471218 463888 471454
rect 463568 471134 463888 471218
rect 463568 470898 463610 471134
rect 463846 470898 463888 471134
rect 463568 470866 463888 470898
rect 479382 451893 479442 636379
rect 479379 451892 479445 451893
rect 479379 451828 479380 451892
rect 479444 451828 479445 451892
rect 479379 451827 479445 451828
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 141008 439174 141328 439206
rect 141008 438938 141050 439174
rect 141286 438938 141328 439174
rect 141008 438854 141328 438938
rect 141008 438618 141050 438854
rect 141286 438618 141328 438854
rect 141008 438586 141328 438618
rect 171728 439174 172048 439206
rect 171728 438938 171770 439174
rect 172006 438938 172048 439174
rect 171728 438854 172048 438938
rect 171728 438618 171770 438854
rect 172006 438618 172048 438854
rect 171728 438586 172048 438618
rect 202448 439174 202768 439206
rect 202448 438938 202490 439174
rect 202726 438938 202768 439174
rect 202448 438854 202768 438938
rect 202448 438618 202490 438854
rect 202726 438618 202768 438854
rect 202448 438586 202768 438618
rect 233168 439174 233488 439206
rect 233168 438938 233210 439174
rect 233446 438938 233488 439174
rect 233168 438854 233488 438938
rect 233168 438618 233210 438854
rect 233446 438618 233488 438854
rect 233168 438586 233488 438618
rect 263888 439174 264208 439206
rect 263888 438938 263930 439174
rect 264166 438938 264208 439174
rect 263888 438854 264208 438938
rect 263888 438618 263930 438854
rect 264166 438618 264208 438854
rect 263888 438586 264208 438618
rect 294608 439174 294928 439206
rect 294608 438938 294650 439174
rect 294886 438938 294928 439174
rect 294608 438854 294928 438938
rect 294608 438618 294650 438854
rect 294886 438618 294928 438854
rect 294608 438586 294928 438618
rect 325328 439174 325648 439206
rect 325328 438938 325370 439174
rect 325606 438938 325648 439174
rect 325328 438854 325648 438938
rect 325328 438618 325370 438854
rect 325606 438618 325648 438854
rect 325328 438586 325648 438618
rect 356048 439174 356368 439206
rect 356048 438938 356090 439174
rect 356326 438938 356368 439174
rect 356048 438854 356368 438938
rect 356048 438618 356090 438854
rect 356326 438618 356368 438854
rect 356048 438586 356368 438618
rect 386768 439174 387088 439206
rect 386768 438938 386810 439174
rect 387046 438938 387088 439174
rect 386768 438854 387088 438938
rect 386768 438618 386810 438854
rect 387046 438618 387088 438854
rect 386768 438586 387088 438618
rect 417488 439174 417808 439206
rect 417488 438938 417530 439174
rect 417766 438938 417808 439174
rect 417488 438854 417808 438938
rect 417488 438618 417530 438854
rect 417766 438618 417808 438854
rect 417488 438586 417808 438618
rect 448208 439174 448528 439206
rect 448208 438938 448250 439174
rect 448486 438938 448528 439174
rect 448208 438854 448528 438938
rect 448208 438618 448250 438854
rect 448486 438618 448528 438854
rect 448208 438586 448528 438618
rect 125648 435454 125968 435486
rect 125648 435218 125690 435454
rect 125926 435218 125968 435454
rect 125648 435134 125968 435218
rect 125648 434898 125690 435134
rect 125926 434898 125968 435134
rect 125648 434866 125968 434898
rect 156368 435454 156688 435486
rect 156368 435218 156410 435454
rect 156646 435218 156688 435454
rect 156368 435134 156688 435218
rect 156368 434898 156410 435134
rect 156646 434898 156688 435134
rect 156368 434866 156688 434898
rect 187088 435454 187408 435486
rect 187088 435218 187130 435454
rect 187366 435218 187408 435454
rect 187088 435134 187408 435218
rect 187088 434898 187130 435134
rect 187366 434898 187408 435134
rect 187088 434866 187408 434898
rect 217808 435454 218128 435486
rect 217808 435218 217850 435454
rect 218086 435218 218128 435454
rect 217808 435134 218128 435218
rect 217808 434898 217850 435134
rect 218086 434898 218128 435134
rect 217808 434866 218128 434898
rect 248528 435454 248848 435486
rect 248528 435218 248570 435454
rect 248806 435218 248848 435454
rect 248528 435134 248848 435218
rect 248528 434898 248570 435134
rect 248806 434898 248848 435134
rect 248528 434866 248848 434898
rect 279248 435454 279568 435486
rect 279248 435218 279290 435454
rect 279526 435218 279568 435454
rect 279248 435134 279568 435218
rect 279248 434898 279290 435134
rect 279526 434898 279568 435134
rect 279248 434866 279568 434898
rect 309968 435454 310288 435486
rect 309968 435218 310010 435454
rect 310246 435218 310288 435454
rect 309968 435134 310288 435218
rect 309968 434898 310010 435134
rect 310246 434898 310288 435134
rect 309968 434866 310288 434898
rect 340688 435454 341008 435486
rect 340688 435218 340730 435454
rect 340966 435218 341008 435454
rect 340688 435134 341008 435218
rect 340688 434898 340730 435134
rect 340966 434898 341008 435134
rect 340688 434866 341008 434898
rect 371408 435454 371728 435486
rect 371408 435218 371450 435454
rect 371686 435218 371728 435454
rect 371408 435134 371728 435218
rect 371408 434898 371450 435134
rect 371686 434898 371728 435134
rect 371408 434866 371728 434898
rect 402128 435454 402448 435486
rect 402128 435218 402170 435454
rect 402406 435218 402448 435454
rect 402128 435134 402448 435218
rect 402128 434898 402170 435134
rect 402406 434898 402448 435134
rect 402128 434866 402448 434898
rect 432848 435454 433168 435486
rect 432848 435218 432890 435454
rect 433126 435218 433168 435454
rect 432848 435134 433168 435218
rect 432848 434898 432890 435134
rect 433126 434898 433168 435134
rect 432848 434866 433168 434898
rect 463568 435454 463888 435486
rect 463568 435218 463610 435454
rect 463846 435218 463888 435454
rect 463568 435134 463888 435218
rect 463568 434898 463610 435134
rect 463846 434898 463888 435134
rect 463568 434866 463888 434898
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 141008 403174 141328 403206
rect 141008 402938 141050 403174
rect 141286 402938 141328 403174
rect 141008 402854 141328 402938
rect 141008 402618 141050 402854
rect 141286 402618 141328 402854
rect 141008 402586 141328 402618
rect 171728 403174 172048 403206
rect 171728 402938 171770 403174
rect 172006 402938 172048 403174
rect 171728 402854 172048 402938
rect 171728 402618 171770 402854
rect 172006 402618 172048 402854
rect 171728 402586 172048 402618
rect 202448 403174 202768 403206
rect 202448 402938 202490 403174
rect 202726 402938 202768 403174
rect 202448 402854 202768 402938
rect 202448 402618 202490 402854
rect 202726 402618 202768 402854
rect 202448 402586 202768 402618
rect 233168 403174 233488 403206
rect 233168 402938 233210 403174
rect 233446 402938 233488 403174
rect 233168 402854 233488 402938
rect 233168 402618 233210 402854
rect 233446 402618 233488 402854
rect 233168 402586 233488 402618
rect 263888 403174 264208 403206
rect 263888 402938 263930 403174
rect 264166 402938 264208 403174
rect 263888 402854 264208 402938
rect 263888 402618 263930 402854
rect 264166 402618 264208 402854
rect 263888 402586 264208 402618
rect 294608 403174 294928 403206
rect 294608 402938 294650 403174
rect 294886 402938 294928 403174
rect 294608 402854 294928 402938
rect 294608 402618 294650 402854
rect 294886 402618 294928 402854
rect 294608 402586 294928 402618
rect 325328 403174 325648 403206
rect 325328 402938 325370 403174
rect 325606 402938 325648 403174
rect 325328 402854 325648 402938
rect 325328 402618 325370 402854
rect 325606 402618 325648 402854
rect 325328 402586 325648 402618
rect 356048 403174 356368 403206
rect 356048 402938 356090 403174
rect 356326 402938 356368 403174
rect 356048 402854 356368 402938
rect 356048 402618 356090 402854
rect 356326 402618 356368 402854
rect 356048 402586 356368 402618
rect 386768 403174 387088 403206
rect 386768 402938 386810 403174
rect 387046 402938 387088 403174
rect 386768 402854 387088 402938
rect 386768 402618 386810 402854
rect 387046 402618 387088 402854
rect 386768 402586 387088 402618
rect 417488 403174 417808 403206
rect 417488 402938 417530 403174
rect 417766 402938 417808 403174
rect 417488 402854 417808 402938
rect 417488 402618 417530 402854
rect 417766 402618 417808 402854
rect 417488 402586 417808 402618
rect 448208 403174 448528 403206
rect 448208 402938 448250 403174
rect 448486 402938 448528 403174
rect 448208 402854 448528 402938
rect 448208 402618 448250 402854
rect 448486 402618 448528 402854
rect 448208 402586 448528 402618
rect 125648 399454 125968 399486
rect 125648 399218 125690 399454
rect 125926 399218 125968 399454
rect 125648 399134 125968 399218
rect 125648 398898 125690 399134
rect 125926 398898 125968 399134
rect 125648 398866 125968 398898
rect 156368 399454 156688 399486
rect 156368 399218 156410 399454
rect 156646 399218 156688 399454
rect 156368 399134 156688 399218
rect 156368 398898 156410 399134
rect 156646 398898 156688 399134
rect 156368 398866 156688 398898
rect 187088 399454 187408 399486
rect 187088 399218 187130 399454
rect 187366 399218 187408 399454
rect 187088 399134 187408 399218
rect 187088 398898 187130 399134
rect 187366 398898 187408 399134
rect 187088 398866 187408 398898
rect 217808 399454 218128 399486
rect 217808 399218 217850 399454
rect 218086 399218 218128 399454
rect 217808 399134 218128 399218
rect 217808 398898 217850 399134
rect 218086 398898 218128 399134
rect 217808 398866 218128 398898
rect 248528 399454 248848 399486
rect 248528 399218 248570 399454
rect 248806 399218 248848 399454
rect 248528 399134 248848 399218
rect 248528 398898 248570 399134
rect 248806 398898 248848 399134
rect 248528 398866 248848 398898
rect 279248 399454 279568 399486
rect 279248 399218 279290 399454
rect 279526 399218 279568 399454
rect 279248 399134 279568 399218
rect 279248 398898 279290 399134
rect 279526 398898 279568 399134
rect 279248 398866 279568 398898
rect 309968 399454 310288 399486
rect 309968 399218 310010 399454
rect 310246 399218 310288 399454
rect 309968 399134 310288 399218
rect 309968 398898 310010 399134
rect 310246 398898 310288 399134
rect 309968 398866 310288 398898
rect 340688 399454 341008 399486
rect 340688 399218 340730 399454
rect 340966 399218 341008 399454
rect 340688 399134 341008 399218
rect 340688 398898 340730 399134
rect 340966 398898 341008 399134
rect 340688 398866 341008 398898
rect 371408 399454 371728 399486
rect 371408 399218 371450 399454
rect 371686 399218 371728 399454
rect 371408 399134 371728 399218
rect 371408 398898 371450 399134
rect 371686 398898 371728 399134
rect 371408 398866 371728 398898
rect 402128 399454 402448 399486
rect 402128 399218 402170 399454
rect 402406 399218 402448 399454
rect 402128 399134 402448 399218
rect 402128 398898 402170 399134
rect 402406 398898 402448 399134
rect 402128 398866 402448 398898
rect 432848 399454 433168 399486
rect 432848 399218 432890 399454
rect 433126 399218 433168 399454
rect 432848 399134 433168 399218
rect 432848 398898 432890 399134
rect 433126 398898 433168 399134
rect 432848 398866 433168 398898
rect 463568 399454 463888 399486
rect 463568 399218 463610 399454
rect 463846 399218 463888 399454
rect 463568 399134 463888 399218
rect 463568 398898 463610 399134
rect 463846 398898 463888 399134
rect 463568 398866 463888 398898
rect 479566 388789 479626 700299
rect 480954 698614 481574 707162
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 483059 700500 483125 700501
rect 483059 700436 483060 700500
rect 483124 700436 483125 700500
rect 483059 700435 483125 700436
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480299 522884 480365 522885
rect 480299 522820 480300 522884
rect 480364 522820 480365 522884
rect 480299 522819 480365 522820
rect 480302 500717 480362 522819
rect 480954 518614 481574 554058
rect 481771 553212 481837 553213
rect 481771 553148 481772 553212
rect 481836 553148 481837 553212
rect 481771 553147 481837 553148
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480299 500716 480365 500717
rect 480299 500652 480300 500716
rect 480364 500652 480365 500716
rect 480299 500651 480365 500652
rect 480954 482614 481574 518058
rect 481774 517309 481834 553147
rect 481955 543420 482021 543421
rect 481955 543356 481956 543420
rect 482020 543356 482021 543420
rect 481955 543355 482021 543356
rect 481771 517308 481837 517309
rect 481771 517244 481772 517308
rect 481836 517244 481837 517308
rect 481771 517243 481837 517244
rect 481771 516900 481837 516901
rect 481771 516836 481772 516900
rect 481836 516836 481837 516900
rect 481771 516835 481837 516836
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 479563 388788 479629 388789
rect 479563 388724 479564 388788
rect 479628 388724 479629 388788
rect 479563 388723 479629 388724
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 122051 293180 122117 293181
rect 122051 293116 122052 293180
rect 122116 293116 122117 293180
rect 122051 293115 122117 293116
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 122054 211037 122114 293115
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 122051 211036 122117 211037
rect 122051 210972 122052 211036
rect 122116 210972 122117 211036
rect 122051 210971 122117 210972
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124674 126334 125294 161778
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 124674 90334 125294 125778
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 124674 54334 125294 89778
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 382054 129014 388167
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 128394 130054 129014 165498
rect 128394 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 129014 130054
rect 128394 129734 129014 129818
rect 128394 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 129014 129734
rect 128394 94054 129014 129498
rect 128394 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 129014 94054
rect 128394 93734 129014 93818
rect 128394 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 129014 93734
rect 128394 58054 129014 93498
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 385774 132734 388167
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 97774 132734 133218
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 132114 61774 132734 97218
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 132114 25774 132734 61218
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 353494 136454 388167
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 173494 136454 208938
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 135834 137494 136454 172938
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 135834 101494 136454 136938
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 363454 146414 388167
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 367174 150134 388167
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 370894 153854 388167
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 374614 157574 388167
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 378334 161294 388167
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 382054 165014 388167
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 385774 168734 388167
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 353494 172454 388167
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 363454 182414 388167
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 367174 186134 388167
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 370894 189854 388167
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 374614 193574 388167
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 378334 197294 388167
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 196674 234334 197294 269778
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 196674 162334 197294 197778
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 382054 201014 388167
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 200394 238054 201014 273498
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 385774 204734 388167
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 206139 381580 206205 381581
rect 206139 381516 206140 381580
rect 206204 381516 206205 381580
rect 206139 381515 206205 381516
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 206142 208997 206202 381515
rect 207834 353494 208454 388167
rect 210371 384300 210437 384301
rect 210371 384236 210372 384300
rect 210436 384236 210437 384300
rect 210371 384235 210437 384236
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 206139 208996 206205 208997
rect 206139 208932 206140 208996
rect 206204 208932 206205 208996
rect 206139 208931 206205 208932
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 173494 208454 208938
rect 210374 207909 210434 384235
rect 217794 363454 218414 388167
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 210371 207908 210437 207909
rect 210371 207844 210372 207908
rect 210436 207844 210437 207908
rect 210371 207843 210437 207844
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 183454 218414 218898
rect 221514 367174 222134 388167
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 225234 370894 225854 388167
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 224355 344180 224421 344181
rect 224355 344116 224356 344180
rect 224420 344116 224421 344180
rect 224355 344115 224421 344116
rect 223251 342684 223317 342685
rect 223251 342620 223252 342684
rect 223316 342620 223317 342684
rect 223251 342619 223317 342620
rect 222883 342004 222949 342005
rect 222883 341940 222884 342004
rect 222948 341940 222949 342004
rect 222883 341939 222949 341940
rect 222699 339556 222765 339557
rect 222699 339492 222700 339556
rect 222764 339492 222765 339556
rect 222699 339491 222765 339492
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 222702 235789 222762 339491
rect 222886 237421 222946 341939
rect 223067 341324 223133 341325
rect 223067 341260 223068 341324
rect 223132 341260 223133 341324
rect 223067 341259 223133 341260
rect 223070 239053 223130 341259
rect 223254 240685 223314 342619
rect 224171 342276 224237 342277
rect 224171 342212 224172 342276
rect 224236 342212 224237 342276
rect 224171 342211 224237 342212
rect 223251 240684 223317 240685
rect 223251 240620 223252 240684
rect 223316 240620 223317 240684
rect 223251 240619 223317 240620
rect 223067 239052 223133 239053
rect 223067 238988 223068 239052
rect 223132 238988 223133 239052
rect 223067 238987 223133 238988
rect 222883 237420 222949 237421
rect 222883 237356 222884 237420
rect 222948 237356 222949 237420
rect 222883 237355 222949 237356
rect 222699 235788 222765 235789
rect 222699 235724 222700 235788
rect 222764 235724 222765 235788
rect 222699 235723 222765 235724
rect 224174 225997 224234 342211
rect 224358 232525 224418 344115
rect 224907 343500 224973 343501
rect 224907 343436 224908 343500
rect 224972 343436 224973 343500
rect 224907 343435 224973 343436
rect 224539 342548 224605 342549
rect 224539 342484 224540 342548
rect 224604 342484 224605 342548
rect 224539 342483 224605 342484
rect 224542 243949 224602 342483
rect 224910 255373 224970 343435
rect 225234 334894 225854 370338
rect 228954 374614 229574 388167
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 227483 343636 227549 343637
rect 227483 343572 227484 343636
rect 227548 343572 227549 343636
rect 227483 343571 227549 343572
rect 227115 343092 227181 343093
rect 227115 343028 227116 343092
rect 227180 343028 227181 343092
rect 227115 343027 227181 343028
rect 226195 341868 226261 341869
rect 226195 341804 226196 341868
rect 226260 341804 226261 341868
rect 226195 341803 226261 341804
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 224907 255372 224973 255373
rect 224907 255308 224908 255372
rect 224972 255308 224973 255372
rect 224907 255307 224973 255308
rect 224539 243948 224605 243949
rect 224539 243884 224540 243948
rect 224604 243884 224605 243948
rect 224539 243883 224605 243884
rect 224355 232524 224421 232525
rect 224355 232460 224356 232524
rect 224420 232460 224421 232524
rect 224355 232459 224421 232460
rect 225234 226894 225854 262338
rect 226198 252109 226258 341803
rect 226931 339964 226997 339965
rect 226931 339900 226932 339964
rect 226996 339900 226997 339964
rect 226931 339899 226997 339900
rect 226747 257820 226813 257821
rect 226747 257756 226748 257820
rect 226812 257756 226813 257820
rect 226747 257755 226813 257756
rect 226750 257410 226810 257755
rect 226382 257350 226810 257410
rect 226195 252108 226261 252109
rect 226195 252044 226196 252108
rect 226260 252044 226261 252108
rect 226195 252043 226261 252044
rect 226382 229261 226442 257350
rect 226563 256732 226629 256733
rect 226563 256668 226564 256732
rect 226628 256668 226629 256732
rect 226563 256667 226629 256668
rect 226566 230893 226626 256667
rect 226934 234157 226994 339899
rect 227118 253741 227178 343027
rect 227299 342412 227365 342413
rect 227299 342348 227300 342412
rect 227364 342348 227365 342412
rect 227299 342347 227365 342348
rect 227302 257005 227362 342347
rect 227486 258637 227546 343571
rect 228954 338614 229574 374058
rect 232674 378334 233294 388167
rect 236394 382054 237014 388167
rect 240114 385774 240734 388167
rect 240114 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 240734 385774
rect 240114 385454 240734 385538
rect 240114 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 240734 385454
rect 239811 384300 239877 384301
rect 239811 384236 239812 384300
rect 239876 384236 239877 384300
rect 239811 384235 239877 384236
rect 239627 382804 239693 382805
rect 239627 382740 239628 382804
rect 239692 382740 239693 382804
rect 239627 382739 239693 382740
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236131 378452 236197 378453
rect 236131 378388 236132 378452
rect 236196 378388 236197 378452
rect 236131 378387 236197 378388
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 230979 345404 231045 345405
rect 230979 345340 230980 345404
rect 231044 345340 231045 345404
rect 230979 345339 231045 345340
rect 230059 344044 230125 344045
rect 230059 343980 230060 344044
rect 230124 343980 230125 344044
rect 230059 343979 230125 343980
rect 229875 343908 229941 343909
rect 229875 343844 229876 343908
rect 229940 343844 229941 343908
rect 229875 343843 229941 343844
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228219 338332 228285 338333
rect 228219 338268 228220 338332
rect 228284 338268 228285 338332
rect 228219 338267 228285 338268
rect 228954 338294 229574 338378
rect 227483 258636 227549 258637
rect 227483 258572 227484 258636
rect 227548 258572 227549 258636
rect 227483 258571 227549 258572
rect 227299 257004 227365 257005
rect 227299 256940 227300 257004
rect 227364 256940 227365 257004
rect 227299 256939 227365 256940
rect 227115 253740 227181 253741
rect 227115 253676 227116 253740
rect 227180 253676 227181 253740
rect 227115 253675 227181 253676
rect 228222 247213 228282 338267
rect 228403 338196 228469 338197
rect 228403 338132 228404 338196
rect 228468 338132 228469 338196
rect 228403 338131 228469 338132
rect 228406 306237 228466 338131
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228403 306236 228469 306237
rect 228403 306172 228404 306236
rect 228468 306172 228469 306236
rect 228403 306171 228469 306172
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228219 247212 228285 247213
rect 228219 247148 228220 247212
rect 228284 247148 228285 247212
rect 228219 247147 228285 247148
rect 226931 234156 226997 234157
rect 226931 234092 226932 234156
rect 226996 234092 226997 234156
rect 226931 234091 226997 234092
rect 226563 230892 226629 230893
rect 226563 230828 226564 230892
rect 226628 230828 226629 230892
rect 226563 230827 226629 230828
rect 228954 230614 229574 266058
rect 229878 248845 229938 343843
rect 230062 250477 230122 343979
rect 230059 250476 230125 250477
rect 230059 250412 230060 250476
rect 230124 250412 230125 250476
rect 230059 250411 230125 250412
rect 229875 248844 229941 248845
rect 229875 248780 229876 248844
rect 229940 248780 229941 248844
rect 229875 248779 229941 248780
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 226379 229260 226445 229261
rect 226379 229196 226380 229260
rect 226444 229196 226445 229260
rect 226379 229195 226445 229196
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 224171 225996 224237 225997
rect 224171 225932 224172 225996
rect 224236 225932 224237 225996
rect 224171 225931 224237 225932
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 219939 216612 220005 216613
rect 219939 216548 219940 216612
rect 220004 216548 220005 216612
rect 219939 216547 220005 216548
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 219942 45525 220002 216547
rect 221514 187174 222134 222618
rect 224171 217700 224237 217701
rect 224171 217636 224172 217700
rect 224236 217636 224237 217700
rect 224171 217635 224237 217636
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 219939 45524 220005 45525
rect 219939 45460 219940 45524
rect 220004 45460 220005 45524
rect 219939 45459 220005 45460
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 224174 7717 224234 217635
rect 225234 190894 225854 226338
rect 228219 215524 228285 215525
rect 228219 215460 228220 215524
rect 228284 215460 228285 215524
rect 228219 215459 228285 215460
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 228222 86325 228282 215459
rect 228954 194614 229574 230058
rect 230982 210085 231042 345339
rect 231163 344452 231229 344453
rect 231163 344388 231164 344452
rect 231228 344388 231229 344452
rect 231163 344387 231229 344388
rect 231166 245581 231226 344387
rect 232674 342334 233294 377778
rect 235763 373284 235829 373285
rect 235763 373220 235764 373284
rect 235828 373220 235829 373284
rect 235763 373219 235829 373220
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 233739 337652 233805 337653
rect 233739 337588 233740 337652
rect 233804 337588 233805 337652
rect 233739 337587 233805 337588
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 270334 233294 305778
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 231163 245580 231229 245581
rect 231163 245516 231164 245580
rect 231228 245516 231229 245580
rect 231163 245515 231229 245516
rect 232674 234334 233294 269778
rect 233742 242317 233802 337587
rect 233739 242316 233805 242317
rect 233739 242252 233740 242316
rect 233804 242252 233805 242316
rect 233739 242251 233805 242252
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232267 227628 232333 227629
rect 232267 227564 232268 227628
rect 232332 227564 232333 227628
rect 232267 227563 232333 227564
rect 232083 224364 232149 224365
rect 232083 224300 232084 224364
rect 232148 224300 232149 224364
rect 232083 224299 232149 224300
rect 231163 213348 231229 213349
rect 231163 213284 231164 213348
rect 231228 213284 231229 213348
rect 231163 213283 231229 213284
rect 230979 210084 231045 210085
rect 230979 210020 230980 210084
rect 231044 210020 231045 210084
rect 230979 210019 231045 210020
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 231166 188869 231226 213283
rect 231163 188868 231229 188869
rect 231163 188804 231164 188868
rect 231228 188804 231229 188868
rect 231163 188803 231229 188804
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 232086 142085 232146 224299
rect 232083 142084 232149 142085
rect 232083 142020 232084 142084
rect 232148 142020 232149 142084
rect 232083 142019 232149 142020
rect 232270 137869 232330 227563
rect 232674 198334 233294 233778
rect 235211 212940 235277 212941
rect 235211 212876 235212 212940
rect 235276 212876 235277 212940
rect 235211 212875 235277 212876
rect 235027 208044 235093 208045
rect 235027 207980 235028 208044
rect 235092 207980 235093 208044
rect 235027 207979 235093 207980
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232267 137868 232333 137869
rect 232267 137804 232268 137868
rect 232332 137804 232333 137868
rect 232267 137803 232333 137804
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228219 86324 228285 86325
rect 228219 86260 228220 86324
rect 228284 86260 228285 86324
rect 228219 86259 228285 86260
rect 228954 86294 229574 86378
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 224171 7716 224237 7717
rect 224171 7652 224172 7716
rect 224236 7652 224237 7716
rect 224171 7651 224237 7652
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 126334 233294 161778
rect 235030 139229 235090 207979
rect 235214 143850 235274 212875
rect 235395 211308 235461 211309
rect 235395 211244 235396 211308
rect 235460 211244 235461 211308
rect 235395 211243 235461 211244
rect 235398 144530 235458 211243
rect 235579 209676 235645 209677
rect 235579 209612 235580 209676
rect 235644 209612 235645 209676
rect 235579 209611 235645 209612
rect 235582 151830 235642 209611
rect 235766 207093 235826 373219
rect 235947 289780 236013 289781
rect 235947 289716 235948 289780
rect 236012 289716 236013 289780
rect 235947 289715 236013 289716
rect 235763 207092 235829 207093
rect 235763 207028 235764 207092
rect 235828 207028 235829 207092
rect 235763 207027 235829 207028
rect 235950 189413 236010 289715
rect 236134 289645 236194 378387
rect 236394 346054 237014 381498
rect 239443 355468 239509 355469
rect 239443 355404 239444 355468
rect 239508 355404 239509 355468
rect 239443 355403 239509 355404
rect 238523 349892 238589 349893
rect 238523 349828 238524 349892
rect 238588 349828 238589 349892
rect 238523 349827 238589 349828
rect 237235 349756 237301 349757
rect 237235 349692 237236 349756
rect 237300 349692 237301 349756
rect 237235 349691 237301 349692
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236131 289644 236197 289645
rect 236131 289580 236132 289644
rect 236196 289580 236197 289644
rect 236131 289579 236197 289580
rect 236394 274054 237014 309498
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236394 238054 237014 273498
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 235947 189412 236013 189413
rect 235947 189348 235948 189412
rect 236012 189348 236013 189412
rect 235947 189347 236013 189348
rect 236394 166054 237014 201498
rect 237238 188325 237298 349691
rect 238339 348396 238405 348397
rect 238339 348332 238340 348396
rect 238404 348332 238405 348396
rect 238339 348331 238405 348332
rect 238155 345812 238221 345813
rect 238155 345748 238156 345812
rect 238220 345748 238221 345812
rect 238155 345747 238221 345748
rect 238158 302565 238218 345747
rect 238342 333981 238402 348331
rect 238526 336293 238586 349827
rect 239259 347172 239325 347173
rect 239259 347108 239260 347172
rect 239324 347108 239325 347172
rect 239259 347107 239325 347108
rect 238523 336292 238589 336293
rect 238523 336228 238524 336292
rect 238588 336228 238589 336292
rect 238523 336227 238589 336228
rect 239262 335205 239322 347107
rect 239259 335204 239325 335205
rect 239259 335140 239260 335204
rect 239324 335140 239325 335204
rect 239259 335139 239325 335140
rect 238339 333980 238405 333981
rect 238339 333916 238340 333980
rect 238404 333916 238405 333980
rect 238339 333915 238405 333916
rect 238155 302564 238221 302565
rect 238155 302500 238156 302564
rect 238220 302500 238221 302564
rect 238155 302499 238221 302500
rect 239446 298077 239506 355403
rect 239443 298076 239509 298077
rect 239443 298012 239444 298076
rect 239508 298012 239509 298076
rect 239443 298011 239509 298012
rect 239630 293793 239690 382739
rect 239627 293792 239693 293793
rect 239627 293728 239628 293792
rect 239692 293728 239693 293792
rect 239627 293727 239693 293728
rect 237971 289644 238037 289645
rect 237971 289580 237972 289644
rect 238036 289580 238037 289644
rect 237971 289579 238037 289580
rect 237419 273868 237485 273869
rect 237419 273804 237420 273868
rect 237484 273804 237485 273868
rect 237419 273803 237485 273804
rect 237422 216749 237482 273803
rect 237419 216748 237485 216749
rect 237419 216684 237420 216748
rect 237484 216684 237485 216748
rect 237419 216683 237485 216684
rect 237235 188324 237301 188325
rect 237235 188260 237236 188324
rect 237300 188260 237301 188324
rect 237235 188259 237301 188260
rect 237974 186149 238034 289579
rect 238155 286380 238221 286381
rect 238155 286316 238156 286380
rect 238220 286316 238221 286380
rect 238155 286315 238221 286316
rect 238158 204645 238218 286315
rect 238523 272508 238589 272509
rect 238523 272444 238524 272508
rect 238588 272444 238589 272508
rect 238523 272443 238589 272444
rect 238339 217836 238405 217837
rect 238339 217772 238340 217836
rect 238404 217772 238405 217836
rect 238339 217771 238405 217772
rect 238155 204644 238221 204645
rect 238155 204580 238156 204644
rect 238220 204580 238221 204644
rect 238155 204579 238221 204580
rect 238155 203148 238221 203149
rect 238155 203084 238156 203148
rect 238220 203084 238221 203148
rect 238155 203083 238221 203084
rect 237971 186148 238037 186149
rect 237971 186084 237972 186148
rect 238036 186084 238037 186148
rect 237971 186083 238037 186084
rect 237787 182748 237853 182749
rect 237787 182684 237788 182748
rect 237852 182684 237853 182748
rect 237787 182683 237853 182684
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 235582 151770 236010 151830
rect 235398 144470 235826 144530
rect 235214 143790 235458 143850
rect 235027 139228 235093 139229
rect 235027 139164 235028 139228
rect 235092 139164 235093 139228
rect 235027 139163 235093 139164
rect 235398 138141 235458 143790
rect 235766 139093 235826 144470
rect 235763 139092 235829 139093
rect 235763 139028 235764 139092
rect 235828 139028 235829 139092
rect 235763 139027 235829 139028
rect 235950 138821 236010 151770
rect 235947 138820 236013 138821
rect 235947 138756 235948 138820
rect 236012 138756 236013 138820
rect 235947 138755 236013 138756
rect 235395 138140 235461 138141
rect 235395 138076 235396 138140
rect 235460 138076 235461 138140
rect 235395 138075 235461 138076
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 130054 237014 165498
rect 237790 140725 237850 182683
rect 237971 181660 238037 181661
rect 237971 181596 237972 181660
rect 238036 181596 238037 181660
rect 237971 181595 238037 181596
rect 237974 140725 238034 181595
rect 237787 140724 237853 140725
rect 237787 140660 237788 140724
rect 237852 140660 237853 140724
rect 237787 140659 237853 140660
rect 237971 140724 238037 140725
rect 237971 140660 237972 140724
rect 238036 140660 238037 140724
rect 237971 140659 238037 140660
rect 238158 137733 238218 203083
rect 238342 141541 238402 217771
rect 238526 206821 238586 272443
rect 239814 218721 239874 384235
rect 240114 349774 240734 385218
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 240114 318905 240734 349218
rect 253794 363454 254414 388167
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 251035 341324 251101 341325
rect 251035 341260 251036 341324
rect 251100 341260 251101 341324
rect 251035 341259 251101 341260
rect 251038 340509 251098 341259
rect 251035 340508 251101 340509
rect 251035 340444 251036 340508
rect 251100 340444 251101 340508
rect 251035 340443 251101 340444
rect 244208 327454 244528 327486
rect 244208 327218 244250 327454
rect 244486 327218 244528 327454
rect 244208 327134 244528 327218
rect 244208 326898 244250 327134
rect 244486 326898 244528 327134
rect 244208 326866 244528 326898
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 318905 254414 326898
rect 257514 367174 258134 388167
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 261234 370894 261854 388167
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 318905 258134 330618
rect 259568 331174 259888 331206
rect 259568 330938 259610 331174
rect 259846 330938 259888 331174
rect 259568 330854 259888 330938
rect 259568 330618 259610 330854
rect 259846 330618 259888 330854
rect 259568 330586 259888 330618
rect 261234 318905 261854 334338
rect 264954 374614 265574 388167
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 318905 265574 338058
rect 268674 378334 269294 388167
rect 268674 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 269294 378334
rect 268674 378014 269294 378098
rect 268674 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 269294 378014
rect 268674 342334 269294 377778
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 268674 318905 269294 341778
rect 272394 382054 273014 388167
rect 272394 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 273014 382054
rect 272394 381734 273014 381818
rect 272394 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 273014 381734
rect 272394 346054 273014 381498
rect 272394 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 273014 346054
rect 272394 345734 273014 345818
rect 272394 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 273014 345734
rect 272394 318905 273014 345498
rect 276114 385774 276734 388167
rect 276114 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 276734 385774
rect 276114 385454 276734 385538
rect 276114 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 276734 385454
rect 276114 349774 276734 385218
rect 276114 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 276734 349774
rect 276114 349454 276734 349538
rect 276114 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 276734 349454
rect 274928 327454 275248 327486
rect 274928 327218 274970 327454
rect 275206 327218 275248 327454
rect 274928 327134 275248 327218
rect 274928 326898 274970 327134
rect 275206 326898 275248 327134
rect 274928 326866 275248 326898
rect 276114 318905 276734 349218
rect 279834 353494 280454 388167
rect 282131 381580 282197 381581
rect 282131 381516 282132 381580
rect 282196 381516 282197 381580
rect 282131 381515 282197 381516
rect 281763 379540 281829 379541
rect 281763 379476 281764 379540
rect 281828 379476 281829 379540
rect 281763 379475 281829 379476
rect 279834 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 280454 353494
rect 279834 353174 280454 353258
rect 279834 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 280454 353174
rect 279834 317494 280454 352938
rect 280659 338876 280725 338877
rect 280659 338812 280660 338876
rect 280724 338812 280725 338876
rect 280659 338811 280725 338812
rect 279834 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 280454 317494
rect 279834 317174 280454 317258
rect 279834 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 280454 317174
rect 259568 295174 259888 295206
rect 259568 294938 259610 295174
rect 259846 294938 259888 295174
rect 259568 294854 259888 294938
rect 259568 294618 259610 294854
rect 259846 294618 259888 294854
rect 259568 294586 259888 294618
rect 244208 291454 244528 291486
rect 244208 291218 244250 291454
rect 244486 291218 244528 291454
rect 244208 291134 244528 291218
rect 244208 290898 244250 291134
rect 244486 290898 244528 291134
rect 244208 290866 244528 290898
rect 274928 291454 275248 291486
rect 274928 291218 274970 291454
rect 275206 291218 275248 291454
rect 274928 291134 275248 291218
rect 274928 290898 274970 291134
rect 275206 290898 275248 291134
rect 274928 290866 275248 290898
rect 279834 281494 280454 316938
rect 280662 291277 280722 338811
rect 281579 337652 281645 337653
rect 281579 337588 281580 337652
rect 281644 337588 281645 337652
rect 281579 337587 281645 337588
rect 280659 291276 280725 291277
rect 280659 291212 280660 291276
rect 280724 291212 280725 291276
rect 280659 291211 280725 291212
rect 279834 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 280454 281494
rect 279834 281174 280454 281258
rect 279834 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 280454 281174
rect 259568 259174 259888 259206
rect 259568 258938 259610 259174
rect 259846 258938 259888 259174
rect 259568 258854 259888 258938
rect 259568 258618 259610 258854
rect 259846 258618 259888 258854
rect 259568 258586 259888 258618
rect 244208 255454 244528 255486
rect 244208 255218 244250 255454
rect 244486 255218 244528 255454
rect 244208 255134 244528 255218
rect 244208 254898 244250 255134
rect 244486 254898 244528 255134
rect 244208 254866 244528 254898
rect 274928 255454 275248 255486
rect 274928 255218 274970 255454
rect 275206 255218 275248 255454
rect 274928 255134 275248 255218
rect 274928 254898 274970 255134
rect 275206 254898 275248 255134
rect 274928 254866 275248 254898
rect 279834 245494 280454 280938
rect 281582 261085 281642 337587
rect 281766 311677 281826 379475
rect 281947 376820 282013 376821
rect 281947 376756 281948 376820
rect 282012 376756 282013 376820
rect 281947 376755 282013 376756
rect 281763 311676 281829 311677
rect 281763 311612 281764 311676
rect 281828 311612 281829 311676
rect 281763 311611 281829 311612
rect 281950 310861 282010 376755
rect 281947 310860 282013 310861
rect 281947 310796 281948 310860
rect 282012 310796 282013 310860
rect 281947 310795 282013 310796
rect 282134 310045 282194 381515
rect 284339 378044 284405 378045
rect 284339 377980 284340 378044
rect 284404 377980 284405 378044
rect 284339 377979 284405 377980
rect 282867 370564 282933 370565
rect 282867 370500 282868 370564
rect 282932 370500 282933 370564
rect 282867 370499 282933 370500
rect 282315 311132 282381 311133
rect 282315 311068 282316 311132
rect 282380 311068 282381 311132
rect 282315 311067 282381 311068
rect 282131 310044 282197 310045
rect 282131 309980 282132 310044
rect 282196 309980 282197 310044
rect 282131 309979 282197 309980
rect 282318 302701 282378 311067
rect 282315 302700 282381 302701
rect 282315 302636 282316 302700
rect 282380 302636 282381 302700
rect 282315 302635 282381 302636
rect 282870 263610 282930 370499
rect 282870 263550 283114 263610
rect 281579 261084 281645 261085
rect 281579 261020 281580 261084
rect 281644 261020 281645 261084
rect 281579 261019 281645 261020
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 259568 223174 259888 223206
rect 259568 222938 259610 223174
rect 259846 222938 259888 223174
rect 259568 222854 259888 222938
rect 259568 222618 259610 222854
rect 259846 222618 259888 222854
rect 259568 222586 259888 222618
rect 244208 219454 244528 219486
rect 244208 219218 244250 219454
rect 244486 219218 244528 219454
rect 244208 219134 244528 219218
rect 244208 218898 244250 219134
rect 244486 218898 244528 219134
rect 244208 218866 244528 218898
rect 274928 219454 275248 219486
rect 274928 219218 274970 219454
rect 275206 219218 275248 219454
rect 274928 219134 275248 219218
rect 274928 218898 274970 219134
rect 275206 218898 275248 219134
rect 274928 218866 275248 218898
rect 239811 218720 239877 218721
rect 239811 218656 239812 218720
rect 239876 218656 239877 218720
rect 239811 218655 239877 218656
rect 279834 209494 280454 244938
rect 283054 244290 283114 263550
rect 282870 244230 283114 244290
rect 280843 211308 280909 211309
rect 280843 211244 280844 211308
rect 280908 211244 280909 211308
rect 280843 211243 280909 211244
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 238523 206820 238589 206821
rect 238523 206756 238524 206820
rect 238588 206756 238589 206820
rect 238523 206755 238589 206756
rect 239259 204780 239325 204781
rect 239259 204716 239260 204780
rect 239324 204716 239325 204780
rect 239259 204715 239325 204716
rect 238339 141540 238405 141541
rect 238339 141476 238340 141540
rect 238404 141476 238405 141540
rect 238339 141475 238405 141476
rect 239262 138549 239322 204715
rect 259568 187174 259888 187206
rect 259568 186938 259610 187174
rect 259846 186938 259888 187174
rect 259568 186854 259888 186938
rect 259568 186618 259610 186854
rect 259846 186618 259888 186854
rect 259568 186586 259888 186618
rect 279371 183564 279437 183565
rect 279371 183500 279372 183564
rect 279436 183500 279437 183564
rect 279371 183499 279437 183500
rect 244208 183454 244528 183486
rect 244208 183218 244250 183454
rect 244486 183218 244528 183454
rect 244208 183134 244528 183218
rect 244208 182898 244250 183134
rect 244486 182898 244528 183134
rect 244208 182866 244528 182898
rect 274928 183454 275248 183486
rect 274928 183218 274970 183454
rect 275206 183218 275248 183454
rect 274928 183134 275248 183218
rect 274928 182898 274970 183134
rect 275206 182898 275248 183134
rect 274928 182866 275248 182898
rect 239627 180640 239693 180641
rect 239627 180576 239628 180640
rect 239692 180576 239693 180640
rect 239627 180575 239693 180576
rect 239630 140725 239690 180575
rect 239811 179552 239877 179553
rect 239811 179488 239812 179552
rect 239876 179488 239877 179552
rect 239811 179487 239877 179488
rect 239627 140724 239693 140725
rect 239627 140660 239628 140724
rect 239692 140660 239693 140724
rect 239627 140659 239693 140660
rect 239259 138548 239325 138549
rect 239259 138484 239260 138548
rect 239324 138484 239325 138548
rect 239259 138483 239325 138484
rect 238155 137732 238221 137733
rect 238155 137668 238156 137732
rect 238220 137668 238221 137732
rect 238155 137667 238221 137668
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 94054 237014 129498
rect 239814 112845 239874 179487
rect 259568 151174 259888 151206
rect 259568 150938 259610 151174
rect 259846 150938 259888 151174
rect 259568 150854 259888 150938
rect 259568 150618 259610 150854
rect 259846 150618 259888 150854
rect 259568 150586 259888 150618
rect 244208 147454 244528 147486
rect 244208 147218 244250 147454
rect 244486 147218 244528 147454
rect 244208 147134 244528 147218
rect 244208 146898 244250 147134
rect 244486 146898 244528 147134
rect 244208 146866 244528 146898
rect 274928 147454 275248 147486
rect 274928 147218 274970 147454
rect 275206 147218 275248 147454
rect 274928 147134 275248 147218
rect 274928 146898 274970 147134
rect 275206 146898 275248 147134
rect 274928 146866 275248 146898
rect 240363 144736 240429 144737
rect 240363 144672 240364 144736
rect 240428 144672 240429 144736
rect 240363 144671 240429 144672
rect 240179 142560 240245 142561
rect 240179 142496 240180 142560
rect 240244 142496 240245 142560
rect 240179 142495 240245 142496
rect 240182 141405 240242 142495
rect 240366 142082 240426 144671
rect 240366 142022 240978 142082
rect 240179 141404 240245 141405
rect 240179 141340 240180 141404
rect 240244 141340 240245 141404
rect 240179 141339 240245 141340
rect 240114 133774 240734 140887
rect 240918 139637 240978 142022
rect 273299 141404 273365 141405
rect 273299 141340 273300 141404
rect 273364 141340 273365 141404
rect 273299 141339 273365 141340
rect 240915 139636 240981 139637
rect 240915 139572 240916 139636
rect 240980 139572 240981 139636
rect 240915 139571 240981 139572
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 239811 112844 239877 112845
rect 239811 112780 239812 112844
rect 239876 112780 239877 112844
rect 239811 112779 239877 112780
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 97774 240734 133218
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 137494 244454 139988
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 101494 244454 136938
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 111454 254414 140887
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 115174 258134 140887
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 118894 261854 140887
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 122614 265574 140887
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 126334 269294 140887
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 90334 269294 125778
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 268674 54334 269294 89778
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 130054 273014 140887
rect 273302 139773 273362 141339
rect 273299 139772 273365 139773
rect 273299 139708 273300 139772
rect 273364 139708 273365 139772
rect 273299 139707 273365 139708
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 272394 94054 273014 129498
rect 272394 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 273014 94054
rect 272394 93734 273014 93818
rect 272394 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 273014 93734
rect 272394 58054 273014 93498
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 133774 276734 140887
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 276114 97774 276734 133218
rect 279374 116517 279434 183499
rect 279834 173494 280454 208938
rect 280659 194988 280725 194989
rect 280659 194924 280660 194988
rect 280724 194924 280725 194988
rect 280659 194923 280725 194924
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 279834 137494 280454 172938
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 279371 116516 279437 116517
rect 279371 116452 279372 116516
rect 279436 116452 279437 116516
rect 279371 116451 279437 116452
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 276114 61774 276734 97218
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 101494 280454 136938
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 279834 65494 280454 100938
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 280662 49333 280722 194923
rect 280846 130525 280906 211243
rect 281763 210492 281829 210493
rect 281763 210428 281764 210492
rect 281828 210428 281829 210492
rect 281763 210427 281829 210428
rect 281579 189276 281645 189277
rect 281579 189212 281580 189276
rect 281644 189212 281645 189276
rect 281579 189211 281645 189212
rect 281027 182748 281093 182749
rect 281027 182684 281028 182748
rect 281092 182684 281093 182748
rect 281027 182683 281093 182684
rect 280843 130524 280909 130525
rect 280843 130460 280844 130524
rect 280908 130460 280909 130524
rect 280843 130459 280909 130460
rect 281030 127669 281090 182683
rect 281027 127668 281093 127669
rect 281027 127604 281028 127668
rect 281092 127604 281093 127668
rect 281027 127603 281093 127604
rect 281582 97205 281642 189211
rect 281766 118149 281826 210427
rect 281947 208860 282013 208861
rect 281947 208796 281948 208860
rect 282012 208796 282013 208860
rect 281947 208795 282013 208796
rect 281950 127805 282010 208795
rect 282131 181932 282197 181933
rect 282131 181868 282132 181932
rect 282196 181868 282197 181932
rect 282131 181867 282197 181868
rect 281947 127804 282013 127805
rect 281947 127740 281948 127804
rect 282012 127740 282013 127804
rect 281947 127739 282013 127740
rect 282134 126309 282194 181867
rect 282870 173773 282930 244230
rect 283419 184380 283485 184381
rect 283419 184316 283420 184380
rect 283484 184316 283485 184380
rect 283419 184315 283485 184316
rect 283051 180300 283117 180301
rect 283051 180236 283052 180300
rect 283116 180236 283117 180300
rect 283051 180235 283117 180236
rect 282867 173772 282933 173773
rect 282867 173708 282868 173772
rect 282932 173708 282933 173772
rect 282867 173707 282933 173708
rect 282131 126308 282197 126309
rect 282131 126244 282132 126308
rect 282196 126244 282197 126308
rect 282131 126243 282197 126244
rect 281763 118148 281829 118149
rect 281763 118084 281764 118148
rect 281828 118084 281829 118148
rect 281763 118083 281829 118084
rect 281579 97204 281645 97205
rect 281579 97140 281580 97204
rect 281644 97140 281645 97204
rect 281579 97139 281645 97140
rect 283054 89045 283114 180235
rect 283235 179484 283301 179485
rect 283235 179420 283236 179484
rect 283300 179420 283301 179484
rect 283235 179419 283301 179420
rect 283238 133109 283298 179419
rect 283235 133108 283301 133109
rect 283235 133044 283236 133108
rect 283300 133044 283301 133108
rect 283235 133043 283301 133044
rect 283422 115157 283482 184315
rect 284342 174589 284402 377979
rect 289794 363454 290414 388167
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 285995 343908 286061 343909
rect 285995 343844 285996 343908
rect 286060 343844 286061 343908
rect 285995 343843 286061 343844
rect 285627 342004 285693 342005
rect 285627 341940 285628 342004
rect 285692 341940 285693 342004
rect 285627 341939 285693 341940
rect 284523 341868 284589 341869
rect 284523 341804 284524 341868
rect 284588 341804 284589 341868
rect 284523 341803 284589 341804
rect 284526 265981 284586 341803
rect 284707 338332 284773 338333
rect 284707 338268 284708 338332
rect 284772 338268 284773 338332
rect 284707 338267 284773 338268
rect 284523 265980 284589 265981
rect 284523 265916 284524 265980
rect 284588 265916 284589 265980
rect 284523 265915 284589 265916
rect 284710 263533 284770 338267
rect 284707 263532 284773 263533
rect 284707 263468 284708 263532
rect 284772 263468 284773 263532
rect 284707 263467 284773 263468
rect 285630 258773 285690 341939
rect 285811 340508 285877 340509
rect 285811 340444 285812 340508
rect 285876 340444 285877 340508
rect 285811 340443 285877 340444
rect 285814 259317 285874 340443
rect 285998 264349 286058 343843
rect 287099 339556 287165 339557
rect 287099 339492 287100 339556
rect 287164 339492 287165 339556
rect 287099 339491 287165 339492
rect 285995 264348 286061 264349
rect 285995 264284 285996 264348
rect 286060 264284 286061 264348
rect 285995 264283 286061 264284
rect 285811 259316 285877 259317
rect 285811 259252 285812 259316
rect 285876 259252 285877 259316
rect 285811 259251 285877 259252
rect 285627 258772 285693 258773
rect 285627 258708 285628 258772
rect 285692 258708 285693 258772
rect 285627 258707 285693 258708
rect 287102 257957 287162 339491
rect 287651 336020 287717 336021
rect 287651 335956 287652 336020
rect 287716 335956 287717 336020
rect 287651 335955 287717 335956
rect 287654 305965 287714 335955
rect 289794 327454 290414 362898
rect 293514 367174 294134 388167
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 290595 338196 290661 338197
rect 290595 338132 290596 338196
rect 290660 338132 290661 338196
rect 290595 338131 290661 338132
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 287651 305964 287717 305965
rect 287651 305900 287652 305964
rect 287716 305900 287717 305964
rect 287651 305899 287717 305900
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 287651 258908 287717 258909
rect 287651 258844 287652 258908
rect 287716 258844 287717 258908
rect 287651 258843 287717 258844
rect 287099 257956 287165 257957
rect 287099 257892 287100 257956
rect 287164 257892 287165 257956
rect 287099 257891 287165 257892
rect 287099 253876 287165 253877
rect 287099 253812 287100 253876
rect 287164 253812 287165 253876
rect 287099 253811 287165 253812
rect 285811 248708 285877 248709
rect 285811 248644 285812 248708
rect 285876 248644 285877 248708
rect 285811 248643 285877 248644
rect 285627 195804 285693 195805
rect 285627 195740 285628 195804
rect 285692 195740 285693 195804
rect 285627 195739 285693 195740
rect 284523 192540 284589 192541
rect 284523 192476 284524 192540
rect 284588 192476 284589 192540
rect 284523 192475 284589 192476
rect 284339 174588 284405 174589
rect 284339 174524 284340 174588
rect 284404 174524 284405 174588
rect 284339 174523 284405 174524
rect 283419 115156 283485 115157
rect 283419 115092 283420 115156
rect 283484 115092 283485 115156
rect 283419 115091 283485 115092
rect 283051 89044 283117 89045
rect 283051 88980 283052 89044
rect 283116 88980 283117 89044
rect 283051 88979 283117 88980
rect 280659 49332 280725 49333
rect 280659 49268 280660 49332
rect 280724 49268 280725 49332
rect 280659 49267 280725 49268
rect 284526 44981 284586 192475
rect 284707 185196 284773 185197
rect 284707 185132 284708 185196
rect 284772 185132 284773 185196
rect 284707 185131 284773 185132
rect 284710 134469 284770 185131
rect 284707 134468 284773 134469
rect 284707 134404 284708 134468
rect 284772 134404 284773 134468
rect 284707 134403 284773 134404
rect 284523 44980 284589 44981
rect 284523 44916 284524 44980
rect 284588 44916 284589 44980
rect 284523 44915 284589 44916
rect 285630 38045 285690 195739
rect 285814 141541 285874 248643
rect 285811 141540 285877 141541
rect 285811 141476 285812 141540
rect 285876 141476 285877 141540
rect 285811 141475 285877 141476
rect 287102 137869 287162 253811
rect 287654 155821 287714 258843
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 288387 246260 288453 246261
rect 288387 246196 288388 246260
rect 288452 246196 288453 246260
rect 288387 246195 288453 246196
rect 287651 155820 287717 155821
rect 287651 155756 287652 155820
rect 287716 155756 287717 155820
rect 287651 155755 287717 155756
rect 288390 138277 288450 246195
rect 288571 242316 288637 242317
rect 288571 242252 288572 242316
rect 288636 242252 288637 242316
rect 288571 242251 288637 242252
rect 288574 138549 288634 242251
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 288939 179212 289005 179213
rect 288939 179148 288940 179212
rect 289004 179148 289005 179212
rect 288939 179147 289005 179148
rect 288755 177852 288821 177853
rect 288755 177788 288756 177852
rect 288820 177788 288821 177852
rect 288755 177787 288821 177788
rect 288758 140453 288818 177787
rect 288942 154189 289002 179147
rect 288939 154188 289005 154189
rect 288939 154124 288940 154188
rect 289004 154124 289005 154188
rect 288939 154123 289005 154124
rect 288939 151740 289005 151741
rect 288939 151676 288940 151740
rect 289004 151676 289005 151740
rect 288939 151675 289005 151676
rect 288755 140452 288821 140453
rect 288755 140388 288756 140452
rect 288820 140388 288821 140452
rect 288755 140387 288821 140388
rect 288755 139500 288821 139501
rect 288755 139436 288756 139500
rect 288820 139436 288821 139500
rect 288755 139435 288821 139436
rect 288571 138548 288637 138549
rect 288571 138484 288572 138548
rect 288636 138484 288637 138548
rect 288571 138483 288637 138484
rect 288387 138276 288453 138277
rect 288387 138212 288388 138276
rect 288452 138212 288453 138276
rect 288387 138211 288453 138212
rect 287099 137868 287165 137869
rect 287099 137804 287100 137868
rect 287164 137804 287165 137868
rect 287099 137803 287165 137804
rect 285627 38044 285693 38045
rect 285627 37980 285628 38044
rect 285692 37980 285693 38044
rect 285627 37979 285693 37980
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 288758 19413 288818 139435
rect 288942 89045 289002 151675
rect 289794 147454 290414 182898
rect 290598 176221 290658 338131
rect 293514 331174 294134 366618
rect 297234 370894 297854 388167
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 294459 358460 294525 358461
rect 294459 358396 294460 358460
rect 294524 358396 294525 358460
rect 294459 358395 294525 358396
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 292619 252108 292685 252109
rect 292619 252044 292620 252108
rect 292684 252044 292685 252108
rect 292619 252043 292685 252044
rect 291331 245444 291397 245445
rect 291331 245380 291332 245444
rect 291396 245380 291397 245444
rect 291331 245379 291397 245380
rect 291147 244628 291213 244629
rect 291147 244564 291148 244628
rect 291212 244564 291213 244628
rect 291147 244563 291213 244564
rect 290779 241500 290845 241501
rect 290779 241436 290780 241500
rect 290844 241436 290845 241500
rect 290779 241435 290845 241436
rect 290595 176220 290661 176221
rect 290595 176156 290596 176220
rect 290660 176156 290661 176220
rect 290595 176155 290661 176156
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 290782 137733 290842 241435
rect 291150 138821 291210 244563
rect 291334 138957 291394 245379
rect 291515 243948 291581 243949
rect 291515 243884 291516 243948
rect 291580 243884 291581 243948
rect 291515 243883 291581 243884
rect 291518 139093 291578 243883
rect 292622 142085 292682 252043
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 294462 175405 294522 358395
rect 295931 337380 295997 337381
rect 295931 337316 295932 337380
rect 295996 337316 295997 337380
rect 295931 337315 295997 337316
rect 294459 175404 294525 175405
rect 294459 175340 294460 175404
rect 294524 175340 294525 175404
rect 294459 175339 294525 175340
rect 295934 157453 295994 337315
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 300954 374614 301574 388167
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 298691 333300 298757 333301
rect 298691 333236 298692 333300
rect 298756 333236 298757 333300
rect 298691 333235 298757 333236
rect 298694 306781 298754 333235
rect 298691 306780 298757 306781
rect 298691 306716 298692 306780
rect 298756 306716 298757 306780
rect 298691 306715 298757 306716
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 295931 157452 295997 157453
rect 295931 157388 295932 157452
rect 295996 157388 295997 157452
rect 295931 157387 295997 157388
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 292619 142084 292685 142085
rect 292619 142020 292620 142084
rect 292684 142020 292685 142084
rect 292619 142019 292685 142020
rect 291515 139092 291581 139093
rect 291515 139028 291516 139092
rect 291580 139028 291581 139092
rect 291515 139027 291581 139028
rect 291331 138956 291397 138957
rect 291331 138892 291332 138956
rect 291396 138892 291397 138956
rect 291331 138891 291397 138892
rect 291147 138820 291213 138821
rect 291147 138756 291148 138820
rect 291212 138756 291213 138820
rect 291147 138755 291213 138756
rect 290779 137732 290845 137733
rect 290779 137668 290780 137732
rect 290844 137668 290845 137732
rect 290779 137667 290845 137668
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 288939 89044 289005 89045
rect 288939 88980 288940 89044
rect 289004 88980 289005 89044
rect 288939 88979 289005 88980
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 288755 19412 288821 19413
rect 288755 19348 288756 19412
rect 288820 19348 288821 19412
rect 288755 19347 288821 19348
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 378334 305294 388167
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 304674 342334 305294 377778
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 304674 306334 305294 341778
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 304674 270334 305294 305778
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 304674 234334 305294 269778
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304674 198334 305294 233778
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 308394 382054 309014 388167
rect 308394 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 309014 382054
rect 308394 381734 309014 381818
rect 308394 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 309014 381734
rect 308394 346054 309014 381498
rect 308394 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 309014 346054
rect 308394 345734 309014 345818
rect 308394 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 309014 345734
rect 308394 310054 309014 345498
rect 308394 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 309014 310054
rect 308394 309734 309014 309818
rect 308394 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 309014 309734
rect 308394 274054 309014 309498
rect 308394 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 309014 274054
rect 308394 273734 309014 273818
rect 308394 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 309014 273734
rect 308394 238054 309014 273498
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 308394 202054 309014 237498
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 308394 166054 309014 201498
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 306971 152556 307037 152557
rect 306971 152492 306972 152556
rect 307036 152492 307037 152556
rect 306971 152491 307037 152492
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 90334 305294 125778
rect 306974 99517 307034 152491
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 306971 99516 307037 99517
rect 306971 99452 306972 99516
rect 307036 99452 307037 99516
rect 306971 99451 307037 99452
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 94054 309014 129498
rect 308394 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 309014 94054
rect 308394 93734 309014 93818
rect 308394 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 309014 93734
rect 308394 58054 309014 93498
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 385774 312734 388167
rect 312114 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 312734 385774
rect 312114 385454 312734 385538
rect 312114 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 312734 385454
rect 312114 349774 312734 385218
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 312114 313774 312734 349218
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 312114 277774 312734 313218
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 312114 241774 312734 277218
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 312114 97774 312734 133218
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 353494 316454 388167
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 315834 317494 316454 352938
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 315834 281494 316454 316938
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 315834 245494 316454 280938
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 363454 326414 388167
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 367174 330134 388167
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 370894 333854 388167
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 374614 337574 388167
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 378334 341294 388167
rect 340674 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 341294 378334
rect 340674 378014 341294 378098
rect 340674 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 341294 378014
rect 340674 342334 341294 377778
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 306334 341294 341778
rect 340674 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 341294 306334
rect 340674 306014 341294 306098
rect 340674 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 341294 306014
rect 340674 270334 341294 305778
rect 340674 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 341294 270334
rect 340674 270014 341294 270098
rect 340674 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 341294 270014
rect 340674 234334 341294 269778
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 344394 382054 345014 388167
rect 344394 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 345014 382054
rect 344394 381734 345014 381818
rect 344394 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 345014 381734
rect 344394 346054 345014 381498
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 344394 310054 345014 345498
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 344394 274054 345014 309498
rect 348114 385774 348734 388167
rect 348114 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 348734 385774
rect 348114 385454 348734 385538
rect 348114 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 348734 385454
rect 348114 349774 348734 385218
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 345611 276724 345677 276725
rect 345611 276660 345612 276724
rect 345676 276660 345677 276724
rect 345611 276659 345677 276660
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 344394 238054 345014 273498
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 342851 195260 342917 195261
rect 342851 195196 342852 195260
rect 342916 195196 342917 195260
rect 342851 195195 342917 195196
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 342854 155005 342914 195195
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 342851 155004 342917 155005
rect 342851 154940 342852 155004
rect 342916 154940 342917 155004
rect 342851 154939 342917 154940
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 130054 345014 165498
rect 345614 156637 345674 276659
rect 348114 241774 348734 277218
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 345611 156636 345677 156637
rect 345611 156572 345612 156636
rect 345676 156572 345677 156636
rect 345611 156571 345677 156572
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 133774 348734 169218
rect 351834 353494 352454 388167
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351834 245494 352454 280938
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351131 153372 351197 153373
rect 351131 153308 351132 153372
rect 351196 153308 351197 153372
rect 351131 153307 351197 153308
rect 351134 139365 351194 153307
rect 351131 139364 351197 139365
rect 351131 139300 351132 139364
rect 351196 139300 351197 139364
rect 351131 139299 351197 139300
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 363454 362414 388167
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 367174 366134 388167
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 370894 369854 388167
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 374614 373574 388167
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 378334 377294 388167
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 382054 381014 388167
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 385774 384734 388167
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 353494 388454 388167
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 363454 398414 388167
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 367174 402134 388167
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 370894 405854 388167
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 374614 409574 388167
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 378334 413294 388167
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 382054 417014 388167
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 385774 420734 388167
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 313774 420734 349218
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 133774 420734 169218
rect 420114 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 420734 133774
rect 420114 133454 420734 133538
rect 420114 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 420734 133454
rect 420114 97774 420734 133218
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 353494 424454 388167
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 423834 317494 424454 352938
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 423834 137494 424454 172938
rect 423834 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 424454 137494
rect 423834 137174 424454 137258
rect 423834 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 424454 137174
rect 423834 101494 424454 136938
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 363454 434414 388167
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 367174 438134 388167
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 370894 441854 388167
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 374614 445574 388167
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 378334 449294 388167
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 306334 449294 341778
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 382054 453014 388167
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 452394 310054 453014 345498
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 385774 456734 388167
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 353494 460454 388167
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 363454 470414 388167
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 367174 474134 388167
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 370894 477854 388167
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 374614 481574 410058
rect 481774 403069 481834 516835
rect 481958 512413 482018 543355
rect 482139 538116 482205 538117
rect 482139 538052 482140 538116
rect 482204 538052 482205 538116
rect 482139 538051 482205 538052
rect 482142 515949 482202 538051
rect 482323 523156 482389 523157
rect 482323 523092 482324 523156
rect 482388 523092 482389 523156
rect 482323 523091 482389 523092
rect 482326 516765 482386 523091
rect 482323 516764 482389 516765
rect 482323 516700 482324 516764
rect 482388 516700 482389 516764
rect 482323 516699 482389 516700
rect 482139 515948 482205 515949
rect 482139 515884 482140 515948
rect 482204 515884 482205 515948
rect 482139 515883 482205 515884
rect 481955 512412 482021 512413
rect 481955 512348 481956 512412
rect 482020 512348 482021 512412
rect 481955 512347 482021 512348
rect 483062 512005 483122 700435
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484347 634676 484413 634677
rect 484347 634612 484348 634676
rect 484412 634612 484413 634676
rect 484347 634611 484413 634612
rect 483243 526692 483309 526693
rect 483243 526628 483244 526692
rect 483308 526628 483309 526692
rect 483243 526627 483309 526628
rect 483059 512004 483125 512005
rect 483059 511940 483060 512004
rect 483124 511940 483125 512004
rect 483059 511939 483125 511940
rect 483246 420749 483306 526627
rect 483427 519076 483493 519077
rect 483427 519012 483428 519076
rect 483492 519012 483493 519076
rect 483427 519011 483493 519012
rect 483430 450669 483490 519011
rect 484350 456381 484410 634611
rect 484674 630334 485294 665778
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 487659 641204 487725 641205
rect 487659 641140 487660 641204
rect 487724 641140 487725 641204
rect 487659 641139 487725 641140
rect 486187 639028 486253 639029
rect 486187 638964 486188 639028
rect 486252 638964 486253 639028
rect 486187 638963 486253 638964
rect 485819 637124 485885 637125
rect 485819 637060 485820 637124
rect 485884 637060 485885 637124
rect 485819 637059 485885 637060
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 486334 485294 521778
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484347 456380 484413 456381
rect 484347 456316 484348 456380
rect 484412 456316 484413 456380
rect 484347 456315 484413 456316
rect 483427 450668 483493 450669
rect 483427 450604 483428 450668
rect 483492 450604 483493 450668
rect 483427 450603 483493 450604
rect 484674 450334 485294 485778
rect 485822 455837 485882 637059
rect 486003 633452 486069 633453
rect 486003 633388 486004 633452
rect 486068 633388 486069 633452
rect 486003 633387 486069 633388
rect 485819 455836 485885 455837
rect 485819 455772 485820 455836
rect 485884 455772 485885 455836
rect 485819 455771 485885 455772
rect 486006 454069 486066 633387
rect 486190 465901 486250 638963
rect 487107 637668 487173 637669
rect 487107 637604 487108 637668
rect 487172 637604 487173 637668
rect 487107 637603 487173 637604
rect 486371 545188 486437 545189
rect 486371 545124 486372 545188
rect 486436 545124 486437 545188
rect 486371 545123 486437 545124
rect 486187 465900 486253 465901
rect 486187 465836 486188 465900
rect 486252 465836 486253 465900
rect 486187 465835 486253 465836
rect 486003 454068 486069 454069
rect 486003 454004 486004 454068
rect 486068 454004 486069 454068
rect 486003 454003 486069 454004
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 483243 420748 483309 420749
rect 483243 420684 483244 420748
rect 483308 420684 483309 420748
rect 483243 420683 483309 420684
rect 483611 420204 483677 420205
rect 483611 420140 483612 420204
rect 483676 420140 483677 420204
rect 483611 420139 483677 420140
rect 481771 403068 481837 403069
rect 481771 403004 481772 403068
rect 481836 403004 481837 403068
rect 481771 403003 481837 403004
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 483614 307597 483674 420139
rect 484674 414334 485294 449778
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 484674 378334 485294 413778
rect 486374 400077 486434 545123
rect 487110 460189 487170 637603
rect 487291 559060 487357 559061
rect 487291 558996 487292 559060
rect 487356 558996 487357 559060
rect 487291 558995 487357 558996
rect 487107 460188 487173 460189
rect 487107 460124 487108 460188
rect 487172 460124 487173 460188
rect 487107 460123 487173 460124
rect 487294 450125 487354 558995
rect 487475 547636 487541 547637
rect 487475 547572 487476 547636
rect 487540 547572 487541 547636
rect 487475 547571 487541 547572
rect 487478 487389 487538 547571
rect 487662 495549 487722 641139
rect 488394 634054 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 489867 654260 489933 654261
rect 489867 654196 489868 654260
rect 489932 654196 489933 654260
rect 489867 654195 489933 654196
rect 489870 653850 489930 654195
rect 489686 653790 489930 653850
rect 489499 641748 489565 641749
rect 489499 641684 489500 641748
rect 489564 641684 489565 641748
rect 489499 641683 489565 641684
rect 489315 637668 489381 637669
rect 489315 637604 489316 637668
rect 489380 637604 489381 637668
rect 489315 637603 489381 637604
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 487659 495548 487725 495549
rect 487659 495484 487660 495548
rect 487724 495484 487725 495548
rect 487659 495483 487725 495484
rect 488394 490054 489014 525498
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 487475 487388 487541 487389
rect 487475 487324 487476 487388
rect 487540 487324 487541 487388
rect 487475 487323 487541 487324
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 487291 450124 487357 450125
rect 487291 450060 487292 450124
rect 487356 450060 487357 450124
rect 487291 450059 487357 450060
rect 488394 418054 489014 453498
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 486371 400076 486437 400077
rect 486371 400012 486372 400076
rect 486436 400012 486437 400076
rect 486371 400011 486437 400012
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 484674 342334 485294 377778
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 483611 307596 483677 307597
rect 483611 307532 483612 307596
rect 483676 307532 483677 307596
rect 483611 307531 483677 307532
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 306334 485294 341778
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 234334 485294 269778
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 484674 198334 485294 233778
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 382054 489014 417498
rect 489318 394909 489378 637603
rect 489502 459101 489562 641683
rect 489499 459100 489565 459101
rect 489499 459036 489500 459100
rect 489564 459036 489565 459100
rect 489499 459035 489565 459036
rect 489315 394908 489381 394909
rect 489315 394844 489316 394908
rect 489380 394844 489381 394908
rect 489315 394843 489381 394844
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 488394 346054 489014 381498
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 488394 310054 489014 345498
rect 489686 339010 489746 653790
rect 492114 637774 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 654737 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 654737 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 654956 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 654737 513854 658338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 654737 517574 662058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 654737 521294 665778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 654956 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 654737 528734 673218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 654737 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 494208 651454 494528 651486
rect 494208 651218 494250 651454
rect 494486 651218 494528 651454
rect 494208 651134 494528 651218
rect 494208 650898 494250 651134
rect 494486 650898 494528 651134
rect 494208 650866 494528 650898
rect 524928 651454 525248 651486
rect 524928 651218 524970 651454
rect 525206 651218 525248 651454
rect 524928 651134 525248 651218
rect 524928 650898 524970 651134
rect 525206 650898 525248 651134
rect 524928 650866 525248 650898
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 601774 492734 637218
rect 541019 636308 541085 636309
rect 541019 636244 541020 636308
rect 541084 636244 541085 636308
rect 541019 636243 541085 636244
rect 539547 629508 539613 629509
rect 539547 629444 539548 629508
rect 539612 629444 539613 629508
rect 539547 629443 539613 629444
rect 509568 619174 509888 619206
rect 509568 618938 509610 619174
rect 509846 618938 509888 619174
rect 509568 618854 509888 618938
rect 509568 618618 509610 618854
rect 509846 618618 509888 618854
rect 509568 618586 509888 618618
rect 494208 615454 494528 615486
rect 494208 615218 494250 615454
rect 494486 615218 494528 615454
rect 494208 615134 494528 615218
rect 494208 614898 494250 615134
rect 494486 614898 494528 615134
rect 494208 614866 494528 614898
rect 524928 615454 525248 615486
rect 524928 615218 524970 615454
rect 525206 615218 525248 615454
rect 524928 615134 525248 615218
rect 524928 614898 524970 615134
rect 525206 614898 525248 615134
rect 524928 614866 525248 614898
rect 539363 607748 539429 607749
rect 539363 607684 539364 607748
rect 539428 607684 539429 607748
rect 539363 607683 539429 607684
rect 538259 601900 538325 601901
rect 538259 601836 538260 601900
rect 538324 601836 538325 601900
rect 538259 601835 538325 601836
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 490419 598228 490485 598229
rect 490419 598164 490420 598228
rect 490484 598164 490485 598228
rect 490419 598163 490485 598164
rect 490051 520028 490117 520029
rect 490051 519964 490052 520028
rect 490116 519964 490117 520028
rect 490051 519963 490117 519964
rect 490054 492693 490114 519963
rect 490235 519620 490301 519621
rect 490235 519556 490236 519620
rect 490300 519556 490301 519620
rect 490235 519555 490301 519556
rect 490238 497589 490298 519555
rect 490422 508605 490482 598163
rect 492114 565774 492734 601218
rect 537339 600540 537405 600541
rect 537339 600476 537340 600540
rect 537404 600476 537405 600540
rect 537339 600475 537405 600476
rect 492995 598228 493061 598229
rect 492995 598164 492996 598228
rect 493060 598164 493061 598228
rect 492995 598163 493061 598164
rect 494099 598228 494165 598229
rect 494099 598164 494100 598228
rect 494164 598164 494165 598228
rect 494099 598163 494165 598164
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 491339 519348 491405 519349
rect 491339 519284 491340 519348
rect 491404 519284 491405 519348
rect 491339 519283 491405 519284
rect 490419 508604 490485 508605
rect 490419 508540 490420 508604
rect 490484 508540 490485 508604
rect 490419 508539 490485 508540
rect 490235 497588 490301 497589
rect 490235 497524 490236 497588
rect 490300 497524 490301 497588
rect 490235 497523 490301 497524
rect 490051 492692 490117 492693
rect 490051 492628 490052 492692
rect 490116 492628 490117 492692
rect 490051 492627 490117 492628
rect 491342 488885 491402 519283
rect 491523 518260 491589 518261
rect 491523 518196 491524 518260
rect 491588 518196 491589 518260
rect 491523 518195 491589 518196
rect 491526 497045 491586 518195
rect 491523 497044 491589 497045
rect 491523 496980 491524 497044
rect 491588 496980 491589 497044
rect 491523 496979 491589 496980
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 491339 488884 491405 488885
rect 491339 488820 491340 488884
rect 491404 488820 491405 488884
rect 491339 488819 491405 488820
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 349774 492734 385218
rect 492998 374781 493058 598163
rect 493179 526012 493245 526013
rect 493179 525948 493180 526012
rect 493244 525948 493245 526012
rect 493179 525947 493245 525948
rect 493182 482901 493242 525947
rect 493363 518124 493429 518125
rect 493363 518060 493364 518124
rect 493428 518060 493429 518124
rect 493363 518059 493429 518060
rect 493366 495957 493426 518059
rect 493363 495956 493429 495957
rect 493363 495892 493364 495956
rect 493428 495892 493429 495956
rect 493363 495891 493429 495892
rect 493179 482900 493245 482901
rect 493179 482836 493180 482900
rect 493244 482836 493245 482900
rect 493179 482835 493245 482836
rect 492995 374780 493061 374781
rect 492995 374716 492996 374780
rect 493060 374716 493061 374780
rect 492995 374715 493061 374716
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 489686 338950 490114 339010
rect 490054 338741 490114 338950
rect 490051 338740 490117 338741
rect 490051 338676 490052 338740
rect 490116 338676 490117 338740
rect 490051 338675 490117 338676
rect 490054 335370 490114 338675
rect 490054 335310 490482 335370
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 238054 489014 273498
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 488394 202054 489014 237498
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 488394 166054 489014 201498
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 490422 46341 490482 335310
rect 492114 313774 492734 349218
rect 494102 345813 494162 598163
rect 495834 569494 496454 600207
rect 496859 598228 496925 598229
rect 496859 598164 496860 598228
rect 496924 598164 496925 598228
rect 496859 598163 496925 598164
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 494283 555388 494349 555389
rect 494283 555324 494284 555388
rect 494348 555324 494349 555388
rect 494283 555323 494349 555324
rect 494286 439381 494346 555323
rect 494467 540156 494533 540157
rect 494467 540092 494468 540156
rect 494532 540092 494533 540156
rect 494467 540091 494533 540092
rect 494470 507925 494530 540091
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495387 533220 495453 533221
rect 495387 533156 495388 533220
rect 495452 533156 495453 533220
rect 495387 533155 495453 533156
rect 495834 533174 496454 533258
rect 495390 520165 495450 533155
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495571 522476 495637 522477
rect 495571 522412 495572 522476
rect 495636 522412 495637 522476
rect 495571 522411 495637 522412
rect 495387 520164 495453 520165
rect 495387 520100 495388 520164
rect 495452 520100 495453 520164
rect 495387 520099 495453 520100
rect 494651 519212 494717 519213
rect 494651 519148 494652 519212
rect 494716 519148 494717 519212
rect 494651 519147 494717 519148
rect 494467 507924 494533 507925
rect 494467 507860 494468 507924
rect 494532 507860 494533 507924
rect 494467 507859 494533 507860
rect 494654 495413 494714 519147
rect 495203 518940 495269 518941
rect 495203 518876 495204 518940
rect 495268 518910 495269 518940
rect 495268 518876 495450 518910
rect 495203 518875 495450 518876
rect 495206 518850 495450 518875
rect 494651 495412 494717 495413
rect 494651 495348 494652 495412
rect 494716 495348 494717 495412
rect 494651 495347 494717 495348
rect 495390 489973 495450 518850
rect 495574 509013 495634 522411
rect 495571 509012 495637 509013
rect 495571 508948 495572 509012
rect 495636 508948 495637 509012
rect 495571 508947 495637 508948
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495387 489972 495453 489973
rect 495387 489908 495388 489972
rect 495452 489908 495453 489972
rect 495387 489907 495453 489908
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 494283 439380 494349 439381
rect 494283 439316 494284 439380
rect 494348 439316 494349 439380
rect 494283 439315 494349 439316
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 353494 496454 388938
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 494099 345812 494165 345813
rect 494099 345748 494100 345812
rect 494164 345748 494165 345812
rect 494099 345747 494165 345748
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 241774 492734 277218
rect 492114 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 492734 241774
rect 492114 241454 492734 241538
rect 492114 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 492734 241454
rect 492114 205774 492734 241218
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 492114 169774 492734 205218
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 133774 492734 169218
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 492114 97774 492734 133218
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 490419 46340 490485 46341
rect 490419 46276 490420 46340
rect 490484 46276 490485 46340
rect 490419 46275 490485 46276
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 317494 496454 352938
rect 496862 350029 496922 598163
rect 501459 596868 501525 596869
rect 501459 596804 501460 596868
rect 501524 596804 501525 596868
rect 501459 596803 501525 596804
rect 498515 559876 498581 559877
rect 498515 559812 498516 559876
rect 498580 559812 498581 559876
rect 498515 559811 498581 559812
rect 498331 553076 498397 553077
rect 498331 553012 498332 553076
rect 498396 553012 498397 553076
rect 498331 553011 498397 553012
rect 498147 531860 498213 531861
rect 498147 531796 498148 531860
rect 498212 531796 498213 531860
rect 498147 531795 498213 531796
rect 497043 525740 497109 525741
rect 497043 525676 497044 525740
rect 497108 525676 497109 525740
rect 497043 525675 497109 525676
rect 497046 494325 497106 525675
rect 497227 518668 497293 518669
rect 497227 518604 497228 518668
rect 497292 518604 497293 518668
rect 497227 518603 497293 518604
rect 497230 498133 497290 518603
rect 497227 498132 497293 498133
rect 497227 498068 497228 498132
rect 497292 498068 497293 498132
rect 497227 498067 497293 498068
rect 497043 494324 497109 494325
rect 497043 494260 497044 494324
rect 497108 494260 497109 494324
rect 497043 494259 497109 494260
rect 498150 415989 498210 531795
rect 498334 489429 498394 553011
rect 498518 504117 498578 559811
rect 501275 557836 501341 557837
rect 501275 557772 501276 557836
rect 501340 557772 501341 557836
rect 501275 557771 501341 557772
rect 501091 554436 501157 554437
rect 501091 554372 501092 554436
rect 501156 554372 501157 554436
rect 501091 554371 501157 554372
rect 499803 554300 499869 554301
rect 499803 554236 499804 554300
rect 499868 554236 499869 554300
rect 499803 554235 499869 554236
rect 499619 554028 499685 554029
rect 499619 553964 499620 554028
rect 499684 553964 499685 554028
rect 499619 553963 499685 553964
rect 498699 545596 498765 545597
rect 498699 545532 498700 545596
rect 498764 545532 498765 545596
rect 498699 545531 498765 545532
rect 498515 504116 498581 504117
rect 498515 504052 498516 504116
rect 498580 504052 498581 504116
rect 498515 504051 498581 504052
rect 498702 493781 498762 545531
rect 498699 493780 498765 493781
rect 498699 493716 498700 493780
rect 498764 493716 498765 493780
rect 498699 493715 498765 493716
rect 498331 489428 498397 489429
rect 498331 489364 498332 489428
rect 498396 489364 498397 489428
rect 498331 489363 498397 489364
rect 499622 443189 499682 553963
rect 499806 488341 499866 554235
rect 500907 550356 500973 550357
rect 500907 550292 500908 550356
rect 500972 550292 500973 550356
rect 500907 550291 500973 550292
rect 500171 548996 500237 548997
rect 500171 548932 500172 548996
rect 500236 548932 500237 548996
rect 500171 548931 500237 548932
rect 499987 524924 500053 524925
rect 499987 524860 499988 524924
rect 500052 524860 500053 524924
rect 499987 524859 500053 524860
rect 499803 488340 499869 488341
rect 499803 488276 499804 488340
rect 499868 488276 499869 488340
rect 499803 488275 499869 488276
rect 499990 483989 500050 524859
rect 500174 507381 500234 548931
rect 500171 507380 500237 507381
rect 500171 507316 500172 507380
rect 500236 507316 500237 507380
rect 500171 507315 500237 507316
rect 500910 493237 500970 550291
rect 501094 498677 501154 554371
rect 501278 505205 501338 557771
rect 501275 505204 501341 505205
rect 501275 505140 501276 505204
rect 501340 505140 501341 505204
rect 501275 505139 501341 505140
rect 501091 498676 501157 498677
rect 501091 498612 501092 498676
rect 501156 498612 501157 498676
rect 501091 498611 501157 498612
rect 500907 493236 500973 493237
rect 500907 493172 500908 493236
rect 500972 493172 500973 493236
rect 500907 493171 500973 493172
rect 499987 483988 500053 483989
rect 499987 483924 499988 483988
rect 500052 483924 500053 483988
rect 499987 483923 500053 483924
rect 499619 443188 499685 443189
rect 499619 443124 499620 443188
rect 499684 443124 499685 443188
rect 499619 443123 499685 443124
rect 498147 415988 498213 415989
rect 498147 415924 498148 415988
rect 498212 415924 498213 415988
rect 498147 415923 498213 415924
rect 496859 350028 496925 350029
rect 496859 349964 496860 350028
rect 496924 349964 496925 350028
rect 496859 349963 496925 349964
rect 501462 325549 501522 596803
rect 505794 579454 506414 600207
rect 508451 595508 508517 595509
rect 508451 595444 508452 595508
rect 508516 595444 508517 595508
rect 508451 595443 508517 595444
rect 506979 594012 507045 594013
rect 506979 593948 506980 594012
rect 507044 593948 507045 594012
rect 506979 593947 507045 593948
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 502747 555116 502813 555117
rect 502747 555052 502748 555116
rect 502812 555052 502813 555116
rect 502747 555051 502813 555052
rect 502379 548860 502445 548861
rect 502379 548796 502380 548860
rect 502444 548796 502445 548860
rect 502379 548795 502445 548796
rect 502382 491061 502442 548795
rect 502563 547500 502629 547501
rect 502563 547436 502564 547500
rect 502628 547436 502629 547500
rect 502563 547435 502629 547436
rect 502566 492149 502626 547435
rect 502750 502485 502810 555051
rect 505139 549132 505205 549133
rect 505139 549068 505140 549132
rect 505204 549068 505205 549132
rect 505139 549067 505205 549068
rect 502931 532404 502997 532405
rect 502931 532340 502932 532404
rect 502996 532340 502997 532404
rect 502931 532339 502997 532340
rect 502934 504661 502994 532339
rect 503667 526284 503733 526285
rect 503667 526220 503668 526284
rect 503732 526220 503733 526284
rect 503667 526219 503733 526220
rect 502931 504660 502997 504661
rect 502931 504596 502932 504660
rect 502996 504596 502997 504660
rect 502931 504595 502997 504596
rect 502747 502484 502813 502485
rect 502747 502420 502748 502484
rect 502812 502420 502813 502484
rect 502747 502419 502813 502420
rect 502563 492148 502629 492149
rect 502563 492084 502564 492148
rect 502628 492084 502629 492148
rect 502563 492083 502629 492084
rect 502379 491060 502445 491061
rect 502379 490996 502380 491060
rect 502444 490996 502445 491060
rect 502379 490995 502445 490996
rect 503670 484533 503730 526219
rect 503851 518532 503917 518533
rect 503851 518468 503852 518532
rect 503916 518468 503917 518532
rect 503851 518467 503917 518468
rect 503854 496501 503914 518467
rect 503851 496500 503917 496501
rect 503851 496436 503852 496500
rect 503916 496436 503917 496500
rect 503851 496435 503917 496436
rect 503667 484532 503733 484533
rect 503667 484468 503668 484532
rect 503732 484468 503733 484532
rect 503667 484467 503733 484468
rect 505142 483445 505202 549067
rect 505794 543454 506414 578898
rect 506611 544372 506677 544373
rect 506611 544308 506612 544372
rect 506676 544308 506677 544372
rect 506611 544307 506677 544308
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505139 483444 505205 483445
rect 505139 483380 505140 483444
rect 505204 483380 505205 483444
rect 505139 483379 505205 483380
rect 505794 471454 506414 506898
rect 506614 501941 506674 544307
rect 506611 501940 506677 501941
rect 506611 501876 506612 501940
rect 506676 501876 506677 501940
rect 506611 501875 506677 501876
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 501459 325548 501525 325549
rect 501459 325484 501460 325548
rect 501524 325484 501525 325548
rect 501459 325483 501525 325484
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 245494 496454 280938
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 495834 209494 496454 244938
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 495834 173494 496454 208938
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 495834 137494 496454 172938
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 495834 101494 496454 136938
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 495834 65494 496454 100938
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 291454 506414 326898
rect 506982 304333 507042 593947
rect 507899 525604 507965 525605
rect 507899 525540 507900 525604
rect 507964 525540 507965 525604
rect 507899 525539 507965 525540
rect 507902 485077 507962 525539
rect 507899 485076 507965 485077
rect 507899 485012 507900 485076
rect 507964 485012 507965 485076
rect 507899 485011 507965 485012
rect 506979 304332 507045 304333
rect 506979 304268 506980 304332
rect 507044 304268 507045 304332
rect 506979 304267 507045 304268
rect 508454 303517 508514 595443
rect 509514 583174 510134 599988
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 513234 586894 513854 600207
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 510843 558380 510909 558381
rect 510843 558316 510844 558380
rect 510908 558316 510909 558380
rect 510843 558315 510909 558316
rect 510659 552804 510725 552805
rect 510659 552740 510660 552804
rect 510724 552740 510725 552804
rect 510659 552739 510725 552740
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 510662 485621 510722 552739
rect 510659 485620 510725 485621
rect 510659 485556 510660 485620
rect 510724 485556 510725 485620
rect 510659 485555 510725 485556
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 510846 441557 510906 558315
rect 511027 558244 511093 558245
rect 511027 558180 511028 558244
rect 511092 558180 511093 558244
rect 511027 558179 511093 558180
rect 511030 442101 511090 558179
rect 512131 552668 512197 552669
rect 512131 552604 512132 552668
rect 512196 552604 512197 552668
rect 512131 552603 512197 552604
rect 511211 546140 511277 546141
rect 511211 546076 511212 546140
rect 511276 546076 511277 546140
rect 511211 546075 511277 546076
rect 511214 499590 511274 546075
rect 511214 499530 511458 499590
rect 511398 486709 511458 499530
rect 511395 486708 511461 486709
rect 511395 486644 511396 486708
rect 511460 486644 511461 486708
rect 511395 486643 511461 486644
rect 512134 486165 512194 552603
rect 513234 550894 513854 586338
rect 516954 590614 517574 600207
rect 520674 594334 521294 600207
rect 526299 599996 526365 599997
rect 522251 599724 522317 599725
rect 522251 599660 522252 599724
rect 522316 599660 522317 599724
rect 522251 599659 522317 599660
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 518019 592652 518085 592653
rect 518019 592588 518020 592652
rect 518084 592588 518085 592652
rect 518019 592587 518085 592588
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 514155 560012 514221 560013
rect 514155 559948 514156 560012
rect 514220 559948 514221 560012
rect 514155 559947 514221 559948
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 512131 486164 512197 486165
rect 512131 486100 512132 486164
rect 512196 486100 512197 486164
rect 512131 486099 512197 486100
rect 511211 485892 511277 485893
rect 511211 485828 511212 485892
rect 511276 485828 511277 485892
rect 511211 485827 511277 485828
rect 511027 442100 511093 442101
rect 511027 442036 511028 442100
rect 511092 442036 511093 442100
rect 511027 442035 511093 442036
rect 510843 441556 510909 441557
rect 510843 441492 510844 441556
rect 510908 441492 510909 441556
rect 510843 441491 510909 441492
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 508451 303516 508517 303517
rect 508451 303452 508452 303516
rect 508516 303452 508517 303516
rect 508451 303451 508517 303452
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 295174 510134 330618
rect 511214 323917 511274 485827
rect 513234 478894 513854 514338
rect 514158 487797 514218 559947
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 514155 487796 514221 487797
rect 514155 487732 514156 487796
rect 514220 487732 514221 487796
rect 514155 487731 514221 487732
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 511211 323916 511277 323917
rect 511211 323852 511212 323916
rect 511276 323852 511277 323916
rect 511211 323851 511277 323852
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 518022 305149 518082 592587
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 522254 309229 522314 599659
rect 522435 599588 522501 599589
rect 522435 599524 522436 599588
rect 522500 599524 522501 599588
rect 522435 599523 522501 599524
rect 522438 317389 522498 599523
rect 524394 598054 525014 599988
rect 526299 599932 526300 599996
rect 526364 599932 526365 599996
rect 526299 599931 526365 599932
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 522435 317388 522501 317389
rect 522435 317324 522436 317388
rect 522500 317324 522501 317388
rect 522435 317323 522501 317324
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 522251 309228 522317 309229
rect 522251 309164 522252 309228
rect 522316 309164 522317 309228
rect 522251 309163 522317 309164
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 518019 305148 518085 305149
rect 518019 305084 518020 305148
rect 518084 305084 518085 305148
rect 518019 305083 518085 305084
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 274054 525014 309498
rect 526302 300253 526362 599931
rect 528114 565774 528734 600207
rect 530531 598228 530597 598229
rect 530531 598164 530532 598228
rect 530596 598164 530597 598228
rect 530531 598163 530597 598164
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 530534 327181 530594 598163
rect 531834 569494 532454 600207
rect 534579 600132 534645 600133
rect 534579 600068 534580 600132
rect 534644 600068 534645 600132
rect 534579 600067 534645 600068
rect 533291 599180 533357 599181
rect 533291 599116 533292 599180
rect 533356 599116 533357 599180
rect 533291 599115 533357 599116
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 530531 327180 530597 327181
rect 530531 327116 530532 327180
rect 530596 327116 530597 327180
rect 530531 327115 530597 327116
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 526299 300252 526365 300253
rect 526299 300188 526300 300252
rect 526364 300188 526365 300252
rect 526299 300187 526365 300188
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 317494 532454 352938
rect 533294 326365 533354 599115
rect 533291 326364 533357 326365
rect 533291 326300 533292 326364
rect 533356 326300 533357 326364
rect 533291 326299 533357 326300
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 534582 301069 534642 600067
rect 536051 598364 536117 598365
rect 536051 598300 536052 598364
rect 536116 598300 536117 598364
rect 536051 598299 536117 598300
rect 536054 328813 536114 598299
rect 536051 328812 536117 328813
rect 536051 328748 536052 328812
rect 536116 328748 536117 328812
rect 536051 328747 536117 328748
rect 537342 301885 537402 600475
rect 537523 599452 537589 599453
rect 537523 599388 537524 599452
rect 537588 599388 537589 599452
rect 537523 599387 537589 599388
rect 537526 308413 537586 599387
rect 538262 324733 538322 601835
rect 538443 601764 538509 601765
rect 538443 601700 538444 601764
rect 538508 601700 538509 601764
rect 538443 601699 538509 601700
rect 538446 327997 538506 601699
rect 538443 327996 538509 327997
rect 538443 327932 538444 327996
rect 538508 327932 538509 327996
rect 538443 327931 538509 327932
rect 538259 324732 538325 324733
rect 538259 324668 538260 324732
rect 538324 324668 538325 324732
rect 538259 324667 538325 324668
rect 539366 311133 539426 607683
rect 539550 315757 539610 629443
rect 539731 626788 539797 626789
rect 539731 626724 539732 626788
rect 539796 626724 539797 626788
rect 539731 626723 539797 626724
rect 539547 315756 539613 315757
rect 539547 315692 539548 315756
rect 539612 315692 539613 315756
rect 539547 315691 539613 315692
rect 539734 314125 539794 626723
rect 539915 624068 539981 624069
rect 539915 624004 539916 624068
rect 539980 624004 539981 624068
rect 539915 624003 539981 624004
rect 539731 314124 539797 314125
rect 539731 314060 539732 314124
rect 539796 314060 539797 314124
rect 539731 314059 539797 314060
rect 539918 312493 539978 624003
rect 540099 603668 540165 603669
rect 540099 603604 540100 603668
rect 540164 603604 540165 603668
rect 540099 603603 540165 603604
rect 540102 599997 540162 603603
rect 540099 599996 540165 599997
rect 540099 599932 540100 599996
rect 540164 599932 540165 599996
rect 540099 599931 540165 599932
rect 541022 319837 541082 636243
rect 541203 619988 541269 619989
rect 541203 619924 541204 619988
rect 541268 619924 541269 619988
rect 541203 619923 541269 619924
rect 541206 381581 541266 619923
rect 541794 615454 542414 650898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 543779 633588 543845 633589
rect 543779 633524 543780 633588
rect 543844 633524 543845 633588
rect 543779 633523 543845 633524
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 543227 610468 543293 610469
rect 543227 610404 543228 610468
rect 543292 610404 543293 610468
rect 543227 610403 543293 610404
rect 542859 609108 542925 609109
rect 542859 609044 542860 609108
rect 542924 609044 542925 609108
rect 542859 609043 542925 609044
rect 542675 606388 542741 606389
rect 542675 606324 542676 606388
rect 542740 606324 542741 606388
rect 542675 606323 542741 606324
rect 542678 600541 542738 606323
rect 542675 600540 542741 600541
rect 542675 600476 542676 600540
rect 542740 600476 542741 600540
rect 542675 600475 542741 600476
rect 542675 600268 542741 600269
rect 542675 600204 542676 600268
rect 542740 600204 542741 600268
rect 542675 600203 542741 600204
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541203 381580 541269 381581
rect 541203 381516 541204 381580
rect 541268 381516 541269 381580
rect 541203 381515 541269 381516
rect 541387 381036 541453 381037
rect 541387 380972 541388 381036
rect 541452 380972 541453 381036
rect 541387 380971 541453 380972
rect 541390 320653 541450 380971
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 542678 336021 542738 600203
rect 542862 595509 542922 609043
rect 543043 601084 543109 601085
rect 543043 601020 543044 601084
rect 543108 601020 543109 601084
rect 543043 601019 543109 601020
rect 542859 595508 542925 595509
rect 542859 595444 542860 595508
rect 542924 595444 542925 595508
rect 542859 595443 542925 595444
rect 543046 592653 543106 601019
rect 543230 594013 543290 610403
rect 543595 594828 543661 594829
rect 543595 594764 543596 594828
rect 543660 594764 543661 594828
rect 543595 594763 543661 594764
rect 543227 594012 543293 594013
rect 543227 593948 543228 594012
rect 543292 593948 543293 594012
rect 543227 593947 543293 593948
rect 543411 593468 543477 593469
rect 543411 593404 543412 593468
rect 543476 593404 543477 593468
rect 543411 593403 543477 593404
rect 543043 592652 543109 592653
rect 543043 592588 543044 592652
rect 543108 592588 543109 592652
rect 543043 592587 543109 592588
rect 543414 420205 543474 593403
rect 543411 420204 543477 420205
rect 543411 420140 543412 420204
rect 543476 420140 543477 420204
rect 543411 420139 543477 420140
rect 542675 336020 542741 336021
rect 542675 335956 542676 336020
rect 542740 335956 542741 336020
rect 542675 335955 542741 335956
rect 543598 333301 543658 594763
rect 543595 333300 543661 333301
rect 543595 333236 543596 333300
rect 543660 333236 543661 333300
rect 543595 333235 543661 333236
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541387 320652 541453 320653
rect 541387 320588 541388 320652
rect 541452 320588 541453 320652
rect 541387 320587 541453 320588
rect 541019 319836 541085 319837
rect 541019 319772 541020 319836
rect 541084 319772 541085 319836
rect 541019 319771 541085 319772
rect 539915 312492 539981 312493
rect 539915 312428 539916 312492
rect 539980 312428 539981 312492
rect 539915 312427 539981 312428
rect 539363 311132 539429 311133
rect 539363 311068 539364 311132
rect 539428 311068 539429 311132
rect 539363 311067 539429 311068
rect 537523 308412 537589 308413
rect 537523 308348 537524 308412
rect 537588 308348 537589 308412
rect 537523 308347 537589 308348
rect 537339 301884 537405 301885
rect 537339 301820 537340 301884
rect 537404 301820 537405 301884
rect 537339 301819 537405 301820
rect 534579 301068 534645 301069
rect 534579 301004 534580 301068
rect 534644 301004 534645 301068
rect 534579 301003 534645 301004
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 291454 542414 326898
rect 543782 318205 543842 633523
rect 545067 632228 545133 632229
rect 545067 632164 545068 632228
rect 545132 632164 545133 632228
rect 545067 632163 545133 632164
rect 543963 618628 544029 618629
rect 543963 618564 543964 618628
rect 544028 618564 544029 618628
rect 543963 618563 544029 618564
rect 543966 599725 544026 618563
rect 543963 599724 544029 599725
rect 543963 599660 543964 599724
rect 544028 599660 544029 599724
rect 543963 599659 544029 599660
rect 545070 599589 545130 632163
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545251 617268 545317 617269
rect 545251 617204 545252 617268
rect 545316 617204 545317 617268
rect 545251 617203 545317 617204
rect 545067 599588 545133 599589
rect 545067 599524 545068 599588
rect 545132 599524 545133 599588
rect 545067 599523 545133 599524
rect 545254 599453 545314 617203
rect 545251 599452 545317 599453
rect 545251 599388 545252 599452
rect 545316 599388 545317 599452
rect 545251 599387 545317 599388
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 555371 683908 555437 683909
rect 555371 683844 555372 683908
rect 555436 683844 555437 683908
rect 555371 683843 555437 683844
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 551139 630868 551205 630869
rect 551139 630804 551140 630868
rect 551204 630804 551205 630868
rect 551139 630803 551205 630804
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 548379 577692 548445 577693
rect 548379 577628 548380 577692
rect 548444 577628 548445 577692
rect 548379 577627 548445 577628
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 547091 524516 547157 524517
rect 547091 524452 547092 524516
rect 547156 524452 547157 524516
rect 547091 524451 547157 524452
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 544331 471476 544397 471477
rect 544331 471412 544332 471476
rect 544396 471412 544397 471476
rect 544331 471411 544397 471412
rect 543779 318204 543845 318205
rect 543779 318140 543780 318204
rect 543844 318140 543845 318204
rect 543779 318139 543845 318140
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 544334 159085 544394 471411
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 544331 159084 544397 159085
rect 544331 159020 544332 159084
rect 544396 159020 544397 159084
rect 544331 159019 544397 159020
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 151174 546134 186618
rect 547094 159901 547154 524451
rect 548382 160717 548442 577627
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 548379 160716 548445 160717
rect 548379 160652 548380 160716
rect 548444 160652 548445 160716
rect 548379 160651 548445 160652
rect 547091 159900 547157 159901
rect 547091 159836 547092 159900
rect 547156 159836 547157 159900
rect 547091 159835 547157 159836
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 154894 549854 190338
rect 551142 161533 551202 630803
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 551139 161532 551205 161533
rect 551139 161468 551140 161532
rect 551204 161468 551205 161532
rect 551139 161467 551205 161468
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 552954 158614 553574 194058
rect 555374 162349 555434 683843
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 558131 418300 558197 418301
rect 558131 418236 558132 418300
rect 558196 418236 558197 418300
rect 558131 418235 558197 418236
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 555371 162348 555437 162349
rect 555371 162284 555372 162348
rect 555436 162284 555437 162348
rect 555371 162283 555437 162284
rect 556674 162334 557294 197778
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 551139 150924 551205 150925
rect 551139 150860 551140 150924
rect 551204 150860 551205 150924
rect 551139 150859 551205 150860
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 551142 19821 551202 150859
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 551139 19820 551205 19821
rect 551139 19756 551140 19820
rect 551204 19756 551205 19820
rect 551139 19755 551205 19756
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 558134 158269 558194 418235
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 558131 158268 558197 158269
rect 558131 158204 558132 158268
rect 558196 158204 558197 158268
rect 558131 158203 558197 158204
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 580211 484668 580277 484669
rect 580211 484604 580212 484668
rect 580276 484604 580277 484668
rect 580211 484603 580277 484604
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 580214 349757 580274 484603
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 580395 365124 580461 365125
rect 580395 365060 580396 365124
rect 580460 365060 580461 365124
rect 580395 365059 580461 365060
rect 580211 349756 580277 349757
rect 580211 349692 580212 349756
rect 580276 349692 580277 349756
rect 580211 349691 580277 349692
rect 580398 337381 580458 365059
rect 580395 337380 580461 337381
rect 580395 337316 580396 337380
rect 580460 337316 580461 337380
rect 580395 337315 580461 337316
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 580211 312084 580277 312085
rect 580211 312020 580212 312084
rect 580276 312020 580277 312084
rect 580211 312019 580277 312020
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 580214 276725 580274 312019
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 580211 276724 580277 276725
rect 580211 276660 580212 276724
rect 580276 276660 580277 276724
rect 580211 276659 580277 276660
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 580211 219060 580277 219061
rect 580211 218996 580212 219060
rect 580276 218996 580277 219060
rect 580211 218995 580277 218996
rect 577794 183454 578414 218898
rect 580214 195261 580274 218995
rect 580211 195260 580277 195261
rect 580211 195196 580212 195260
rect 580276 195196 580277 195260
rect 580211 195195 580277 195196
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 580211 89044 580277 89045
rect 580211 88980 580212 89044
rect 580276 88980 580277 89044
rect 580211 88979 580277 88980
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 580214 59669 580274 88979
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 580211 59668 580277 59669
rect 580211 59604 580212 59668
rect 580276 59604 580277 59668
rect 580211 59603 580277 59604
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 79610 618938 79846 619174
rect 79610 618618 79846 618854
rect 110330 618938 110566 619174
rect 110330 618618 110566 618854
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 125690 615218 125926 615454
rect 125690 614898 125926 615134
rect 135866 605258 136102 605494
rect 136186 605258 136422 605494
rect 135866 604938 136102 605174
rect 136186 604938 136422 605174
rect 79610 582938 79846 583174
rect 79610 582618 79846 582854
rect 110330 582938 110566 583174
rect 110330 582618 110566 582854
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 125690 579218 125926 579454
rect 125690 578898 125926 579134
rect 135866 569258 136102 569494
rect 136186 569258 136422 569494
rect 135866 568938 136102 569174
rect 136186 568938 136422 569174
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 64250 471218 64486 471454
rect 64250 470898 64486 471134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 54250 255218 54486 255454
rect 54250 254898 54486 255134
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 64250 435218 64486 435454
rect 64250 434898 64486 435134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 64250 399218 64486 399454
rect 64250 398898 64486 399134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 79610 510938 79846 511174
rect 79610 510618 79846 510854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 79610 474938 79846 475174
rect 79610 474618 79846 474854
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 79610 438938 79846 439174
rect 79610 438618 79846 438854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 79610 402938 79846 403174
rect 79610 402618 79846 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 88706 558098 88942 558334
rect 89026 558098 89262 558334
rect 88706 557778 88942 558014
rect 89026 557778 89262 558014
rect 88706 522098 88942 522334
rect 89026 522098 89262 522334
rect 88706 521778 88942 522014
rect 89026 521778 89262 522014
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 92426 525818 92662 526054
rect 92746 525818 92982 526054
rect 92426 525498 92662 525734
rect 92746 525498 92982 525734
rect 96146 529538 96382 529774
rect 96466 529538 96702 529774
rect 96146 529218 96382 529454
rect 96466 529218 96702 529454
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 92426 489818 92662 490054
rect 92746 489818 92982 490054
rect 92426 489498 92662 489734
rect 92746 489498 92982 489734
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 94970 471218 95206 471454
rect 94970 470898 95206 471134
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 94970 435218 95206 435454
rect 94970 434898 95206 435134
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 94970 399218 95206 399454
rect 94970 398898 95206 399134
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 92426 309818 92662 310054
rect 92746 309818 92982 310054
rect 92426 309498 92662 309734
rect 92746 309498 92982 309734
rect 92426 273818 92662 274054
rect 92746 273818 92982 274054
rect 92426 273498 92662 273734
rect 92746 273498 92982 273734
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 99866 533258 100102 533494
rect 100186 533258 100422 533494
rect 99866 532938 100102 533174
rect 100186 532938 100422 533174
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 110330 510938 110566 511174
rect 110330 510618 110566 510854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 110330 474938 110566 475174
rect 110330 474618 110566 474854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 110330 438938 110566 439174
rect 110330 438618 110566 438854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 110330 402938 110566 403174
rect 110330 402618 110566 402854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 99866 281258 100102 281494
rect 100186 281258 100422 281494
rect 99866 280938 100102 281174
rect 100186 280938 100422 281174
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 84970 255218 85206 255454
rect 84970 254898 85206 255134
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 54250 219218 54486 219454
rect 54250 218898 54486 219134
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 69610 222938 69846 223174
rect 69610 222618 69846 222854
rect 100330 222938 100566 223174
rect 100330 222618 100566 222854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 84970 219218 85206 219454
rect 84970 218898 85206 219134
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 55080 75218 55316 75454
rect 55080 74898 55316 75134
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 59174 78938 59410 79174
rect 59174 78618 59410 78854
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 63268 75218 63504 75454
rect 63268 74898 63504 75134
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 67362 78938 67598 79174
rect 67362 78618 67598 78854
rect 71456 75218 71692 75454
rect 71456 74898 71692 75134
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 75550 78938 75786 79174
rect 75550 78618 75786 78854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 79644 75218 79880 75454
rect 79644 74898 79880 75134
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 83738 78938 83974 79174
rect 83738 78618 83974 78854
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 88706 126098 88942 126334
rect 89026 126098 89262 126334
rect 88706 125778 88942 126014
rect 89026 125778 89262 126014
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 165818 92662 166054
rect 92746 165818 92982 166054
rect 92426 165498 92662 165734
rect 92746 165498 92982 165734
rect 92426 129818 92662 130054
rect 92746 129818 92982 130054
rect 92426 129498 92662 129734
rect 92746 129498 92982 129734
rect 92426 93818 92662 94054
rect 92746 93818 92982 94054
rect 92426 93498 92662 93734
rect 92746 93498 92982 93734
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 169538 96382 169774
rect 96466 169538 96702 169774
rect 96146 169218 96382 169454
rect 96466 169218 96702 169454
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 96146 97538 96382 97774
rect 96466 97538 96702 97774
rect 96146 97218 96382 97454
rect 96466 97218 96702 97454
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 173258 100102 173494
rect 100186 173258 100422 173494
rect 99866 172938 100102 173174
rect 100186 172938 100422 173174
rect 99866 137258 100102 137494
rect 100186 137258 100422 137494
rect 99866 136938 100102 137174
rect 100186 136938 100422 137174
rect 99866 101258 100102 101494
rect 100186 101258 100422 101494
rect 99866 100938 100102 101174
rect 100186 100938 100422 101174
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 124706 558098 124942 558334
rect 125026 558098 125262 558334
rect 124706 557778 124942 558014
rect 125026 557778 125262 558014
rect 124706 522098 124942 522334
rect 125026 522098 125262 522334
rect 124706 521778 124942 522014
rect 125026 521778 125262 522014
rect 135866 533258 136102 533494
rect 136186 533258 136422 533494
rect 135866 532938 136102 533174
rect 136186 532938 136422 533174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 199610 618938 199846 619174
rect 199610 618618 199846 618854
rect 230330 618938 230566 619174
rect 230330 618618 230566 618854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 184250 615218 184486 615454
rect 184250 614898 184486 615134
rect 214970 615218 215206 615454
rect 214970 614898 215206 615134
rect 245690 615218 245926 615454
rect 245690 614898 245926 615134
rect 199610 582938 199846 583174
rect 199610 582618 199846 582854
rect 230330 582938 230566 583174
rect 230330 582618 230566 582854
rect 184250 579218 184486 579454
rect 184250 578898 184486 579134
rect 214970 579218 215206 579454
rect 214970 578898 215206 579134
rect 245690 579218 245926 579454
rect 245690 578898 245926 579134
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 268706 594098 268942 594334
rect 269026 594098 269262 594334
rect 268706 593778 268942 594014
rect 269026 593778 269262 594014
rect 268706 558098 268942 558334
rect 269026 558098 269262 558334
rect 268706 557778 268942 558014
rect 269026 557778 269262 558014
rect 268706 522098 268942 522334
rect 269026 522098 269262 522334
rect 268706 521778 268942 522014
rect 269026 521778 269262 522014
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 272426 597818 272662 598054
rect 272746 597818 272982 598054
rect 272426 597498 272662 597734
rect 272746 597498 272982 597734
rect 272426 561818 272662 562054
rect 272746 561818 272982 562054
rect 272426 561498 272662 561734
rect 272746 561498 272982 561734
rect 276146 601538 276382 601774
rect 276466 601538 276702 601774
rect 276146 601218 276382 601454
rect 276466 601218 276702 601454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 279866 605258 280102 605494
rect 280186 605258 280422 605494
rect 279866 604938 280102 605174
rect 280186 604938 280422 605174
rect 276146 565538 276382 565774
rect 276466 565538 276702 565774
rect 276146 565218 276382 565454
rect 276466 565218 276702 565454
rect 272426 525818 272662 526054
rect 272746 525818 272982 526054
rect 272426 525498 272662 525734
rect 272746 525498 272982 525734
rect 279866 569258 280102 569494
rect 280186 569258 280422 569494
rect 279866 568938 280102 569174
rect 280186 568938 280422 569174
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 279866 533258 280102 533494
rect 280186 533258 280422 533494
rect 279866 532938 280102 533174
rect 280186 532938 280422 533174
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 319610 618938 319846 619174
rect 319610 618618 319846 618854
rect 350330 618938 350566 619174
rect 350330 618618 350566 618854
rect 304250 615218 304486 615454
rect 304250 614898 304486 615134
rect 334970 615218 335206 615454
rect 334970 614898 335206 615134
rect 365690 615218 365926 615454
rect 365690 614898 365926 615134
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 319610 582938 319846 583174
rect 319610 582618 319846 582854
rect 350330 582938 350566 583174
rect 350330 582618 350566 582854
rect 304250 579218 304486 579454
rect 304250 578898 304486 579134
rect 334970 579218 335206 579454
rect 334970 578898 335206 579134
rect 365690 579218 365926 579454
rect 365690 578898 365926 579134
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 304706 522098 304942 522334
rect 305026 522098 305262 522334
rect 304706 521778 304942 522014
rect 305026 521778 305262 522014
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 340706 522098 340942 522334
rect 341026 522098 341262 522334
rect 340706 521778 340942 522014
rect 341026 521778 341262 522014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 141050 510938 141286 511174
rect 141050 510618 141286 510854
rect 171770 510938 172006 511174
rect 171770 510618 172006 510854
rect 202490 510938 202726 511174
rect 202490 510618 202726 510854
rect 233210 510938 233446 511174
rect 233210 510618 233446 510854
rect 263930 510938 264166 511174
rect 263930 510618 264166 510854
rect 294650 510938 294886 511174
rect 294650 510618 294886 510854
rect 325370 510938 325606 511174
rect 325370 510618 325606 510854
rect 356090 510938 356326 511174
rect 356090 510618 356326 510854
rect 386810 510938 387046 511174
rect 386810 510618 387046 510854
rect 417530 510938 417766 511174
rect 417530 510618 417766 510854
rect 448250 510938 448486 511174
rect 448250 510618 448486 510854
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 310010 507218 310246 507454
rect 310010 506898 310246 507134
rect 340730 507218 340966 507454
rect 340730 506898 340966 507134
rect 371450 507218 371686 507454
rect 371450 506898 371686 507134
rect 402170 507218 402406 507454
rect 402170 506898 402406 507134
rect 432890 507218 433126 507454
rect 432890 506898 433126 507134
rect 463610 507218 463846 507454
rect 463610 506898 463846 507134
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 141050 474938 141286 475174
rect 141050 474618 141286 474854
rect 171770 474938 172006 475174
rect 171770 474618 172006 474854
rect 202490 474938 202726 475174
rect 202490 474618 202726 474854
rect 233210 474938 233446 475174
rect 233210 474618 233446 474854
rect 263930 474938 264166 475174
rect 263930 474618 264166 474854
rect 294650 474938 294886 475174
rect 294650 474618 294886 474854
rect 325370 474938 325606 475174
rect 325370 474618 325606 474854
rect 356090 474938 356326 475174
rect 356090 474618 356326 474854
rect 386810 474938 387046 475174
rect 386810 474618 387046 474854
rect 417530 474938 417766 475174
rect 417530 474618 417766 474854
rect 448250 474938 448486 475174
rect 448250 474618 448486 474854
rect 125690 471218 125926 471454
rect 125690 470898 125926 471134
rect 156410 471218 156646 471454
rect 156410 470898 156646 471134
rect 187130 471218 187366 471454
rect 187130 470898 187366 471134
rect 217850 471218 218086 471454
rect 217850 470898 218086 471134
rect 248570 471218 248806 471454
rect 248570 470898 248806 471134
rect 279290 471218 279526 471454
rect 279290 470898 279526 471134
rect 310010 471218 310246 471454
rect 310010 470898 310246 471134
rect 340730 471218 340966 471454
rect 340730 470898 340966 471134
rect 371450 471218 371686 471454
rect 371450 470898 371686 471134
rect 402170 471218 402406 471454
rect 402170 470898 402406 471134
rect 432890 471218 433126 471454
rect 432890 470898 433126 471134
rect 463610 471218 463846 471454
rect 463610 470898 463846 471134
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 141050 438938 141286 439174
rect 141050 438618 141286 438854
rect 171770 438938 172006 439174
rect 171770 438618 172006 438854
rect 202490 438938 202726 439174
rect 202490 438618 202726 438854
rect 233210 438938 233446 439174
rect 233210 438618 233446 438854
rect 263930 438938 264166 439174
rect 263930 438618 264166 438854
rect 294650 438938 294886 439174
rect 294650 438618 294886 438854
rect 325370 438938 325606 439174
rect 325370 438618 325606 438854
rect 356090 438938 356326 439174
rect 356090 438618 356326 438854
rect 386810 438938 387046 439174
rect 386810 438618 387046 438854
rect 417530 438938 417766 439174
rect 417530 438618 417766 438854
rect 448250 438938 448486 439174
rect 448250 438618 448486 438854
rect 125690 435218 125926 435454
rect 125690 434898 125926 435134
rect 156410 435218 156646 435454
rect 156410 434898 156646 435134
rect 187130 435218 187366 435454
rect 187130 434898 187366 435134
rect 217850 435218 218086 435454
rect 217850 434898 218086 435134
rect 248570 435218 248806 435454
rect 248570 434898 248806 435134
rect 279290 435218 279526 435454
rect 279290 434898 279526 435134
rect 310010 435218 310246 435454
rect 310010 434898 310246 435134
rect 340730 435218 340966 435454
rect 340730 434898 340966 435134
rect 371450 435218 371686 435454
rect 371450 434898 371686 435134
rect 402170 435218 402406 435454
rect 402170 434898 402406 435134
rect 432890 435218 433126 435454
rect 432890 434898 433126 435134
rect 463610 435218 463846 435454
rect 463610 434898 463846 435134
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 141050 402938 141286 403174
rect 141050 402618 141286 402854
rect 171770 402938 172006 403174
rect 171770 402618 172006 402854
rect 202490 402938 202726 403174
rect 202490 402618 202726 402854
rect 233210 402938 233446 403174
rect 233210 402618 233446 402854
rect 263930 402938 264166 403174
rect 263930 402618 264166 402854
rect 294650 402938 294886 403174
rect 294650 402618 294886 402854
rect 325370 402938 325606 403174
rect 325370 402618 325606 402854
rect 356090 402938 356326 403174
rect 356090 402618 356326 402854
rect 386810 402938 387046 403174
rect 386810 402618 387046 402854
rect 417530 402938 417766 403174
rect 417530 402618 417766 402854
rect 448250 402938 448486 403174
rect 448250 402618 448486 402854
rect 125690 399218 125926 399454
rect 125690 398898 125926 399134
rect 156410 399218 156646 399454
rect 156410 398898 156646 399134
rect 187130 399218 187366 399454
rect 187130 398898 187366 399134
rect 217850 399218 218086 399454
rect 217850 398898 218086 399134
rect 248570 399218 248806 399454
rect 248570 398898 248806 399134
rect 279290 399218 279526 399454
rect 279290 398898 279526 399134
rect 310010 399218 310246 399454
rect 310010 398898 310246 399134
rect 340730 399218 340966 399454
rect 340730 398898 340966 399134
rect 371450 399218 371686 399454
rect 371450 398898 371686 399134
rect 402170 399218 402406 399454
rect 402170 398898 402406 399134
rect 432890 399218 433126 399454
rect 432890 398898 433126 399134
rect 463610 399218 463846 399454
rect 463610 398898 463846 399134
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 128426 129818 128662 130054
rect 128746 129818 128982 130054
rect 128426 129498 128662 129734
rect 128746 129498 128982 129734
rect 128426 93818 128662 94054
rect 128746 93818 128982 94054
rect 128426 93498 128662 93734
rect 128746 93498 128982 93734
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 240146 385538 240382 385774
rect 240466 385538 240702 385774
rect 240146 385218 240382 385454
rect 240466 385218 240702 385454
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 244250 327218 244486 327454
rect 244250 326898 244486 327134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 259610 330938 259846 331174
rect 259610 330618 259846 330854
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 268706 378098 268942 378334
rect 269026 378098 269262 378334
rect 268706 377778 268942 378014
rect 269026 377778 269262 378014
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 272426 381818 272662 382054
rect 272746 381818 272982 382054
rect 272426 381498 272662 381734
rect 272746 381498 272982 381734
rect 272426 345818 272662 346054
rect 272746 345818 272982 346054
rect 272426 345498 272662 345734
rect 272746 345498 272982 345734
rect 276146 385538 276382 385774
rect 276466 385538 276702 385774
rect 276146 385218 276382 385454
rect 276466 385218 276702 385454
rect 276146 349538 276382 349774
rect 276466 349538 276702 349774
rect 276146 349218 276382 349454
rect 276466 349218 276702 349454
rect 274970 327218 275206 327454
rect 274970 326898 275206 327134
rect 279866 353258 280102 353494
rect 280186 353258 280422 353494
rect 279866 352938 280102 353174
rect 280186 352938 280422 353174
rect 279866 317258 280102 317494
rect 280186 317258 280422 317494
rect 279866 316938 280102 317174
rect 280186 316938 280422 317174
rect 259610 294938 259846 295174
rect 259610 294618 259846 294854
rect 244250 291218 244486 291454
rect 244250 290898 244486 291134
rect 274970 291218 275206 291454
rect 274970 290898 275206 291134
rect 279866 281258 280102 281494
rect 280186 281258 280422 281494
rect 279866 280938 280102 281174
rect 280186 280938 280422 281174
rect 259610 258938 259846 259174
rect 259610 258618 259846 258854
rect 244250 255218 244486 255454
rect 244250 254898 244486 255134
rect 274970 255218 275206 255454
rect 274970 254898 275206 255134
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 259610 222938 259846 223174
rect 259610 222618 259846 222854
rect 244250 219218 244486 219454
rect 244250 218898 244486 219134
rect 274970 219218 275206 219454
rect 274970 218898 275206 219134
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 259610 186938 259846 187174
rect 259610 186618 259846 186854
rect 244250 183218 244486 183454
rect 244250 182898 244486 183134
rect 274970 183218 275206 183454
rect 274970 182898 275206 183134
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 259610 150938 259846 151174
rect 259610 150618 259846 150854
rect 244250 147218 244486 147454
rect 244250 146898 244486 147134
rect 274970 147218 275206 147454
rect 274970 146898 275206 147134
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 272426 93818 272662 94054
rect 272746 93818 272982 94054
rect 272426 93498 272662 93734
rect 272746 93498 272982 93734
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 308426 381818 308662 382054
rect 308746 381818 308982 382054
rect 308426 381498 308662 381734
rect 308746 381498 308982 381734
rect 308426 345818 308662 346054
rect 308746 345818 308982 346054
rect 308426 345498 308662 345734
rect 308746 345498 308982 345734
rect 308426 309818 308662 310054
rect 308746 309818 308982 310054
rect 308426 309498 308662 309734
rect 308746 309498 308982 309734
rect 308426 273818 308662 274054
rect 308746 273818 308982 274054
rect 308426 273498 308662 273734
rect 308746 273498 308982 273734
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 93818 308662 94054
rect 308746 93818 308982 94054
rect 308426 93498 308662 93734
rect 308746 93498 308982 93734
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 385538 312382 385774
rect 312466 385538 312702 385774
rect 312146 385218 312382 385454
rect 312466 385218 312702 385454
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 378098 340942 378334
rect 341026 378098 341262 378334
rect 340706 377778 340942 378014
rect 341026 377778 341262 378014
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 340706 306098 340942 306334
rect 341026 306098 341262 306334
rect 340706 305778 340942 306014
rect 341026 305778 341262 306014
rect 340706 270098 340942 270334
rect 341026 270098 341262 270334
rect 340706 269778 340942 270014
rect 341026 269778 341262 270014
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 344426 381818 344662 382054
rect 344746 381818 344982 382054
rect 344426 381498 344662 381734
rect 344746 381498 344982 381734
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 348146 385538 348382 385774
rect 348466 385538 348702 385774
rect 348146 385218 348382 385454
rect 348466 385218 348702 385454
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 420146 133538 420382 133774
rect 420466 133538 420702 133774
rect 420146 133218 420382 133454
rect 420466 133218 420702 133454
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 423866 137258 424102 137494
rect 424186 137258 424422 137494
rect 423866 136938 424102 137174
rect 424186 136938 424422 137174
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 494250 651218 494486 651454
rect 494250 650898 494486 651134
rect 524970 651218 525206 651454
rect 524970 650898 525206 651134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 509610 618938 509846 619174
rect 509610 618618 509846 618854
rect 494250 615218 494486 615454
rect 494250 614898 494486 615134
rect 524970 615218 525206 615454
rect 524970 614898 525206 615134
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 492146 241538 492382 241774
rect 492466 241538 492702 241774
rect 492146 241218 492382 241454
rect 492466 241218 492702 241454
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 494250 651454
rect 494486 651218 524970 651454
rect 525206 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 494250 651134
rect 494486 650898 524970 651134
rect 525206 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 79610 619174
rect 79846 618938 110330 619174
rect 110566 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 199610 619174
rect 199846 618938 230330 619174
rect 230566 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 319610 619174
rect 319846 618938 350330 619174
rect 350566 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509610 619174
rect 509846 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 79610 618854
rect 79846 618618 110330 618854
rect 110566 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 199610 618854
rect 199846 618618 230330 618854
rect 230566 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 319610 618854
rect 319846 618618 350330 618854
rect 350566 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509610 618854
rect 509846 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 125690 615454
rect 125926 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 184250 615454
rect 184486 615218 214970 615454
rect 215206 615218 245690 615454
rect 245926 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 304250 615454
rect 304486 615218 334970 615454
rect 335206 615218 365690 615454
rect 365926 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 494250 615454
rect 494486 615218 524970 615454
rect 525206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 125690 615134
rect 125926 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 184250 615134
rect 184486 614898 214970 615134
rect 215206 614898 245690 615134
rect 245926 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 304250 615134
rect 304486 614898 334970 615134
rect 335206 614898 365690 615134
rect 365926 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 494250 615134
rect 494486 614898 524970 615134
rect 525206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 79610 583174
rect 79846 582938 110330 583174
rect 110566 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 199610 583174
rect 199846 582938 230330 583174
rect 230566 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 319610 583174
rect 319846 582938 350330 583174
rect 350566 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 79610 582854
rect 79846 582618 110330 582854
rect 110566 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 199610 582854
rect 199846 582618 230330 582854
rect 230566 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 319610 582854
rect 319846 582618 350330 582854
rect 350566 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 125690 579454
rect 125926 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 184250 579454
rect 184486 579218 214970 579454
rect 215206 579218 245690 579454
rect 245926 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 304250 579454
rect 304486 579218 334970 579454
rect 335206 579218 365690 579454
rect 365926 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 125690 579134
rect 125926 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 184250 579134
rect 184486 578898 214970 579134
rect 215206 578898 245690 579134
rect 245926 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 304250 579134
rect 304486 578898 334970 579134
rect 335206 578898 365690 579134
rect 365926 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 79610 511174
rect 79846 510938 110330 511174
rect 110566 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 141050 511174
rect 141286 510938 171770 511174
rect 172006 510938 202490 511174
rect 202726 510938 233210 511174
rect 233446 510938 263930 511174
rect 264166 510938 294650 511174
rect 294886 510938 325370 511174
rect 325606 510938 356090 511174
rect 356326 510938 386810 511174
rect 387046 510938 417530 511174
rect 417766 510938 448250 511174
rect 448486 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 79610 510854
rect 79846 510618 110330 510854
rect 110566 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 141050 510854
rect 141286 510618 171770 510854
rect 172006 510618 202490 510854
rect 202726 510618 233210 510854
rect 233446 510618 263930 510854
rect 264166 510618 294650 510854
rect 294886 510618 325370 510854
rect 325606 510618 356090 510854
rect 356326 510618 386810 510854
rect 387046 510618 417530 510854
rect 417766 510618 448250 510854
rect 448486 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 310010 507454
rect 310246 507218 340730 507454
rect 340966 507218 371450 507454
rect 371686 507218 402170 507454
rect 402406 507218 432890 507454
rect 433126 507218 463610 507454
rect 463846 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 310010 507134
rect 310246 506898 340730 507134
rect 340966 506898 371450 507134
rect 371686 506898 402170 507134
rect 402406 506898 432890 507134
rect 433126 506898 463610 507134
rect 463846 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 79610 475174
rect 79846 474938 110330 475174
rect 110566 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 141050 475174
rect 141286 474938 171770 475174
rect 172006 474938 202490 475174
rect 202726 474938 233210 475174
rect 233446 474938 263930 475174
rect 264166 474938 294650 475174
rect 294886 474938 325370 475174
rect 325606 474938 356090 475174
rect 356326 474938 386810 475174
rect 387046 474938 417530 475174
rect 417766 474938 448250 475174
rect 448486 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 79610 474854
rect 79846 474618 110330 474854
rect 110566 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 141050 474854
rect 141286 474618 171770 474854
rect 172006 474618 202490 474854
rect 202726 474618 233210 474854
rect 233446 474618 263930 474854
rect 264166 474618 294650 474854
rect 294886 474618 325370 474854
rect 325606 474618 356090 474854
rect 356326 474618 386810 474854
rect 387046 474618 417530 474854
rect 417766 474618 448250 474854
rect 448486 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 64250 471454
rect 64486 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 94970 471454
rect 95206 471218 125690 471454
rect 125926 471218 156410 471454
rect 156646 471218 187130 471454
rect 187366 471218 217850 471454
rect 218086 471218 248570 471454
rect 248806 471218 279290 471454
rect 279526 471218 310010 471454
rect 310246 471218 340730 471454
rect 340966 471218 371450 471454
rect 371686 471218 402170 471454
rect 402406 471218 432890 471454
rect 433126 471218 463610 471454
rect 463846 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 64250 471134
rect 64486 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 94970 471134
rect 95206 470898 125690 471134
rect 125926 470898 156410 471134
rect 156646 470898 187130 471134
rect 187366 470898 217850 471134
rect 218086 470898 248570 471134
rect 248806 470898 279290 471134
rect 279526 470898 310010 471134
rect 310246 470898 340730 471134
rect 340966 470898 371450 471134
rect 371686 470898 402170 471134
rect 402406 470898 432890 471134
rect 433126 470898 463610 471134
rect 463846 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 79610 439174
rect 79846 438938 110330 439174
rect 110566 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 141050 439174
rect 141286 438938 171770 439174
rect 172006 438938 202490 439174
rect 202726 438938 233210 439174
rect 233446 438938 263930 439174
rect 264166 438938 294650 439174
rect 294886 438938 325370 439174
rect 325606 438938 356090 439174
rect 356326 438938 386810 439174
rect 387046 438938 417530 439174
rect 417766 438938 448250 439174
rect 448486 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 79610 438854
rect 79846 438618 110330 438854
rect 110566 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 141050 438854
rect 141286 438618 171770 438854
rect 172006 438618 202490 438854
rect 202726 438618 233210 438854
rect 233446 438618 263930 438854
rect 264166 438618 294650 438854
rect 294886 438618 325370 438854
rect 325606 438618 356090 438854
rect 356326 438618 386810 438854
rect 387046 438618 417530 438854
rect 417766 438618 448250 438854
rect 448486 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 64250 435454
rect 64486 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 94970 435454
rect 95206 435218 125690 435454
rect 125926 435218 156410 435454
rect 156646 435218 187130 435454
rect 187366 435218 217850 435454
rect 218086 435218 248570 435454
rect 248806 435218 279290 435454
rect 279526 435218 310010 435454
rect 310246 435218 340730 435454
rect 340966 435218 371450 435454
rect 371686 435218 402170 435454
rect 402406 435218 432890 435454
rect 433126 435218 463610 435454
rect 463846 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 64250 435134
rect 64486 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 94970 435134
rect 95206 434898 125690 435134
rect 125926 434898 156410 435134
rect 156646 434898 187130 435134
rect 187366 434898 217850 435134
rect 218086 434898 248570 435134
rect 248806 434898 279290 435134
rect 279526 434898 310010 435134
rect 310246 434898 340730 435134
rect 340966 434898 371450 435134
rect 371686 434898 402170 435134
rect 402406 434898 432890 435134
rect 433126 434898 463610 435134
rect 463846 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 79610 403174
rect 79846 402938 110330 403174
rect 110566 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 141050 403174
rect 141286 402938 171770 403174
rect 172006 402938 202490 403174
rect 202726 402938 233210 403174
rect 233446 402938 263930 403174
rect 264166 402938 294650 403174
rect 294886 402938 325370 403174
rect 325606 402938 356090 403174
rect 356326 402938 386810 403174
rect 387046 402938 417530 403174
rect 417766 402938 448250 403174
rect 448486 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 79610 402854
rect 79846 402618 110330 402854
rect 110566 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 141050 402854
rect 141286 402618 171770 402854
rect 172006 402618 202490 402854
rect 202726 402618 233210 402854
rect 233446 402618 263930 402854
rect 264166 402618 294650 402854
rect 294886 402618 325370 402854
rect 325606 402618 356090 402854
rect 356326 402618 386810 402854
rect 387046 402618 417530 402854
rect 417766 402618 448250 402854
rect 448486 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 64250 399454
rect 64486 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 94970 399454
rect 95206 399218 125690 399454
rect 125926 399218 156410 399454
rect 156646 399218 187130 399454
rect 187366 399218 217850 399454
rect 218086 399218 248570 399454
rect 248806 399218 279290 399454
rect 279526 399218 310010 399454
rect 310246 399218 340730 399454
rect 340966 399218 371450 399454
rect 371686 399218 402170 399454
rect 402406 399218 432890 399454
rect 433126 399218 463610 399454
rect 463846 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 64250 399134
rect 64486 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 94970 399134
rect 95206 398898 125690 399134
rect 125926 398898 156410 399134
rect 156646 398898 187130 399134
rect 187366 398898 217850 399134
rect 218086 398898 248570 399134
rect 248806 398898 279290 399134
rect 279526 398898 310010 399134
rect 310246 398898 340730 399134
rect 340966 398898 371450 399134
rect 371686 398898 402170 399134
rect 402406 398898 432890 399134
rect 433126 398898 463610 399134
rect 463846 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 259610 331174
rect 259846 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 259610 330854
rect 259846 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 244250 327454
rect 244486 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 274970 327454
rect 275206 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 244250 327134
rect 244486 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 274970 327134
rect 275206 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 259610 295174
rect 259846 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 259610 294854
rect 259846 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 244250 291454
rect 244486 291218 274970 291454
rect 275206 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 244250 291134
rect 244486 290898 274970 291134
rect 275206 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 259610 259174
rect 259846 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 259610 258854
rect 259846 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 54250 255454
rect 54486 255218 84970 255454
rect 85206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 244250 255454
rect 244486 255218 274970 255454
rect 275206 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 54250 255134
rect 54486 254898 84970 255134
rect 85206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 244250 255134
rect 244486 254898 274970 255134
rect 275206 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 69610 223174
rect 69846 222938 100330 223174
rect 100566 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 259610 223174
rect 259846 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 69610 222854
rect 69846 222618 100330 222854
rect 100566 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 259610 222854
rect 259846 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 54250 219454
rect 54486 219218 84970 219454
rect 85206 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 244250 219454
rect 244486 219218 274970 219454
rect 275206 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 54250 219134
rect 54486 218898 84970 219134
rect 85206 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 244250 219134
rect 244486 218898 274970 219134
rect 275206 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 259610 187174
rect 259846 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 259610 186854
rect 259846 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 244250 183454
rect 244486 183218 274970 183454
rect 275206 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 244250 183134
rect 244486 182898 274970 183134
rect 275206 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 259610 151174
rect 259846 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 259610 150854
rect 259846 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 244250 147454
rect 244486 147218 274970 147454
rect 275206 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 244250 147134
rect 244486 146898 274970 147134
rect 275206 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 59174 79174
rect 59410 78938 67362 79174
rect 67598 78938 75550 79174
rect 75786 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 83738 79174
rect 83974 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 59174 78854
rect 59410 78618 67362 78854
rect 67598 78618 75550 78854
rect 75786 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 83738 78854
rect 83974 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 55080 75454
rect 55316 75218 63268 75454
rect 63504 75218 71456 75454
rect 71692 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 79644 75454
rect 79880 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 55080 75134
rect 55316 74898 63268 75134
rect 63504 74898 71456 75134
rect 71692 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 79644 75134
rect 79880 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use ci2406_z80  ci2406_z80
timestamp 0
transform 1 0 50000 0 1 200000
box 0 0 60000 60000
use execution_unit  eu0
timestamp 0
transform 1 0 60000 0 1 560000
box 0 0 75000 75000
use execution_unit  eu1
timestamp 0
transform 1 0 180000 0 1 560000
box 0 0 75000 75000
use execution_unit  eu2
timestamp 0
transform 1 0 300000 0 1 560000
box 0 0 75000 75000
use multiplexer  multiplexer
timestamp 0
transform 1 0 240000 0 1 140000
box 0 0 40000 200000
use scrapcpu  scrapcpu
timestamp 0
transform 1 0 490000 0 1 600000
box 0 0 50000 55000
use unused_tie  unused_tie
timestamp 0
transform 1 0 50000 0 1 50000
box 0 0 35000 35000
use vliw  vliw
timestamp 0
transform 1 0 60000 0 1 390000
box 0 0 420000 128000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 198167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 260449 74414 558575 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 633097 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 198167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 260449 110414 389988 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 634540 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 519809 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 633097 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 633097 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 140887 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 318905 254414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 633097 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 519809 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 633097 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 633097 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 519809 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 519809 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 388167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 519809 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 600207 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 654737 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 198167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 260449 81854 558575 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 633097 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 558575 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 633097 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 519809 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 633097 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 633097 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 140887 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 318905 261854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 519809 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 519809 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 633097 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 633097 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 519809 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 519809 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 388167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 519809 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 600207 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 654737 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 198167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 260449 89294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 633097 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 633097 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 519809 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 519809 197294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 633097 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 519809 233294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 633097 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 140887 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 318905 269294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 519809 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 519809 305294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 633097 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 519809 341294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 633097 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 519809 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 519809 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 388167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 519809 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 600207 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 654737 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 198167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 260449 60734 558575 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 633097 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 198167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 260449 96734 558575 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 633097 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 633097 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 519809 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 633097 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 140887 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 318905 240734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 633097 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 140887 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 318905 276734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 519809 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 633097 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 633097 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 519809 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 519809 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 388167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 519809 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 600207 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 654737 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 198167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 260449 93014 558575 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 633097 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 633097 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 519809 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 633097 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 633097 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 140887 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 318905 273014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 519809 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 633097 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 633097 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 519809 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 519809 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 388167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 519809 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 599988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 654956 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 198167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 260449 64454 389988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 634540 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 198167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 260449 100454 558575 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 633097 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 519809 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 519809 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 633097 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 139988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 633097 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 519809 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 633097 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 633097 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 519809 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 519809 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 388167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 519809 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 600207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 654737 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 600207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 654737 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 198167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 260449 78134 558575 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 633097 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 558575 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 633097 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 519809 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 633097 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 633097 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 140887 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 318905 258134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 519809 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 519809 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 633097 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 634540 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 519809 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 519809 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 388167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 519809 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 599988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 654956 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 198167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 260449 85574 558575 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 633097 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 558575 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 633097 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 519809 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 633097 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 633097 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 140887 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 318905 265574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 519809 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 633097 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 633097 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 633097 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 519809 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 388167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 519809 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 600207 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 654737 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
