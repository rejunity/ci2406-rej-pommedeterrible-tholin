* NGSPICE file created from wrapped_as1802.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

.subckt wrapped_as1802 custom_settings[0] custom_settings[10] custom_settings[11]
+ custom_settings[12] custom_settings[13] custom_settings[14] custom_settings[15]
+ custom_settings[16] custom_settings[17] custom_settings[18] custom_settings[19]
+ custom_settings[1] custom_settings[20] custom_settings[21] custom_settings[22] custom_settings[23]
+ custom_settings[24] custom_settings[25] custom_settings[26] custom_settings[27]
+ custom_settings[28] custom_settings[29] custom_settings[2] custom_settings[3] custom_settings[4]
+ custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8] custom_settings[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
+ io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
XANTENNA__4563__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6209__A2 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4315__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6914_ _6932_/C _6910_/C _7020_/A vssd1 vssd1 vccd1 vccd1 _6914_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout162_A _7558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6845_ _6845_/A _6845_/B vssd1 vssd1 vccd1 vccd1 _6887_/A sky130_fd_sc_hd__nor2_1
XANTENNA__6917__B1 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6776_ _6822_/A _6774_/Y _6765_/X vssd1 vssd1 vccd1 vccd1 _6790_/S sky130_fd_sc_hd__a21o_4
X_3988_ _3988_/A _3988_/B _3988_/C vssd1 vssd1 vccd1 vccd1 _4015_/B sky130_fd_sc_hd__and3_2
X_5727_ _5727_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__or2_1
XFILLER_0_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5658_ _6581_/A _6518_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5658_/X sky130_fd_sc_hd__and3_1
XANTENNA__4251__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4609_ _4600_/Y _4603_/Y _5024_/S vssd1 vssd1 vccd1 vccd1 _4609_/X sky130_fd_sc_hd__mux2_1
X_5589_ _5854_/C _5589_/B _5589_/C vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold362 _5205_/X vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _7437_/Q vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
X_7328_ _7424_/CLK _7328_/D vssd1 vssd1 vccd1 vccd1 _7328_/Q sky130_fd_sc_hd__dfxtp_1
Xhold351 _7205_/X vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold384 _5227_/X vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _5271_/X vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _7354_/Q vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
X_7259_ _7541_/CLK _7259_/D vssd1 vssd1 vccd1 vccd1 _7259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5408__A0 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4845__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6384__B2 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3817__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer7 _5605_/X vssd1 vssd1 vccd1 vccd1 _5609_/B sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4242__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3924__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6300__A _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5350__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output56_A _4003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7587_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4870__A1 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5414__A3 _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4960_ input25/X _4959_/X _5031_/S vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__mux2_1
X_3911_ _7279_/Q _7594_/Q _7263_/Q _7487_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3912_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4891_ _6048_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4891_/Y sky130_fd_sc_hd__nand2_1
X_3842_ _3915_/A _3836_/X _7363_/Q vssd1 vssd1 vccd1 vccd1 _3842_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6630_ _6630_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6685_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3808__S0 _7360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6561_ _6611_/A _6561_/B vssd1 vssd1 vccd1 vccd1 _6603_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5512_ _5530_/A _5512_/B vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__and2_1
X_3773_ _6911_/A _4036_/A vssd1 vssd1 vccd1 vccd1 _3962_/C sky130_fd_sc_hd__or2_2
X_6492_ _6521_/A _6521_/D _6491_/X _6468_/Y vssd1 vssd1 vccd1 vccd1 _6496_/B sky130_fd_sc_hd__a211o_1
X_5443_ hold90/A _6683_/B vssd1 vssd1 vccd1 vccd1 _5460_/A sky130_fd_sc_hd__nor2_2
X_5374_ _4685_/X _5373_/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7471_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4233__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4325_ _4323_/X _4324_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4325_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7025__B _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7113_ _7102_/B _7111_/X _7112_/X _6220_/C vssd1 vssd1 vccd1 vccd1 _7113_/X sky130_fd_sc_hd__a31o_1
Xfanout116 _3664_/Y vssd1 vssd1 vccd1 vccd1 _3931_/S sky130_fd_sc_hd__buf_4
Xfanout127 hold663/X vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__buf_6
Xfanout138 _6827_/A vssd1 vssd1 vccd1 vccd1 _6710_/A sky130_fd_sc_hd__clkbuf_8
Xfanout105 _3684_/X vssd1 vssd1 vccd1 vccd1 _6413_/S sky130_fd_sc_hd__clkbuf_8
X_4256_ _4254_/X _4255_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7044_ _7078_/A _7044_/B _7044_/C _7044_/D vssd1 vssd1 vccd1 vccd1 _7044_/X sky130_fd_sc_hd__or4_1
Xfanout149 _6637_/A vssd1 vssd1 vccd1 vccd1 _5854_/C sky130_fd_sc_hd__buf_4
X_4187_ _4401_/S _4183_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4187_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4613__A1 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5496__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6828_ _6836_/B _6828_/B vssd1 vssd1 vccd1 vccd1 _6828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4377__B1 _4320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6759_ _6759_/A _6759_/B vssd1 vssd1 vccd1 vccd1 _6759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6118__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4224__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6120__A _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold170 _4965_/X vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _5161_/X vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _6171_/X vssd1 vssd1 vccd1 vccd1 _7519_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5170__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7097__S _7551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6109__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5345__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5089_/X _4973_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__mux2_1
X_4110_ _4107_/Y _4108_/X _4109_/X _3901_/B vssd1 vssd1 vccd1 vccd1 _4111_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _5977_/B _7554_/Q _3698_/A _6417_/B vssd1 vssd1 vccd1 vccd1 _6416_/A sky130_fd_sc_hd__a31o_1
XANTENNA__5080__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4843__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5992_ _6015_/B _6015_/C _4027_/Y _4021_/A vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4943_ _6066_/A _4917_/A _4942_/Y vssd1 vssd1 vccd1 vccd1 _4943_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3829__A _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6348__A1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4874_ _4902_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4875_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6613_ _6613_/A _6613_/B vssd1 vssd1 vccd1 vccd1 _6613_/Y sky130_fd_sc_hd__xnor2_1
X_7593_ _7593_/CLK _7593_/D vssd1 vssd1 vccd1 vccd1 _7593_/Q sky130_fd_sc_hd__dfxtp_1
X_3825_ _7268_/Q _7608_/Q _7600_/Q _7616_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3825_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5020__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6899__A2 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6544_ _6544_/A vssd1 vssd1 vccd1 vccd1 _6544_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout125_A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3756_ _6374_/A _6413_/S vssd1 vssd1 vccd1 vccd1 _6220_/B sky130_fd_sc_hd__nand2_4
X_6475_ _6532_/A _6476_/B _6474_/A vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__a21bo_1
X_5426_ _7497_/Q _6683_/B vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__or2_1
X_3687_ _5977_/B _7554_/Q vssd1 vssd1 vccd1 vccd1 _4007_/A sky130_fd_sc_hd__or2_4
XFILLER_0_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4531__A0 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6520__A1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5357_ _5357_/A _5393_/B _7193_/C vssd1 vssd1 vccd1 vccd1 _5374_/S sky130_fd_sc_hd__or3b_4
XANTENNA__6875__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5288_ hold209/X _4849_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _7428_/D sky130_fd_sc_hd__mux2_1
X_4308_ _4360_/B _4307_/X _4304_/Y vssd1 vssd1 vccd1 vccd1 _6062_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5087__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4239_ _5002_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6086__S _6086_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7027_ _6306_/B _7024_/X _6311_/A _6922_/B vssd1 vssd1 vccd1 vccd1 _7027_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4834__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4826__C _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5938__B _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4334__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3739__A _7556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4445__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5165__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4053__A2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4590_ hold620/X _4638_/C _4529_/S vssd1 vssd1 vccd1 vccd1 _4590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5075__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4513__A0 _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6260_ _6311_/A _6808_/B vssd1 vssd1 vccd1 vccd1 _6945_/B sky130_fd_sc_hd__nor2_1
X_5211_ hold323/X _5038_/X _5211_/S vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__mux2_1
X_6191_ _6191_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6191_/X sky130_fd_sc_hd__or2_1
X_5142_ _5376_/A _7176_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5157_/S sky130_fd_sc_hd__and3_4
XFILLER_0_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5069__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5073_ hold279/X _5015_/X _5075_/S vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4816__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4277__C1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4024_ _6375_/C _4279_/C vssd1 vssd1 vccd1 vccd1 _4263_/B sky130_fd_sc_hd__nand2_4
XANTENNA__6018__B1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5241__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4154__S _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ _6920_/A _3965_/D _4122_/C _6922_/A vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__a211o_1
X_4926_ _4208_/A _4924_/X _6096_/A vssd1 vssd1 vccd1 vccd1 _4926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4857_ _4974_/B _4266_/Y _4856_/Y _4123_/A vssd1 vssd1 vccd1 vccd1 _4857_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _7376_/Q _7304_/Q _7296_/Q _7288_/Q _7360_/Q _7361_/Q vssd1 vssd1 vccd1 vccd1
+ _3808_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7576_ _7587_/CLK _7576_/D vssd1 vssd1 vccd1 vccd1 _7576_/Q sky130_fd_sc_hd__dfxtp_1
X_4788_ _5393_/A _5393_/B _5159_/C vssd1 vssd1 vccd1 vccd1 _4806_/S sky130_fd_sc_hd__or3b_4
XFILLER_0_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6527_ _6575_/A _6569_/B _6569_/C _6563_/A _6505_/X vssd1 vssd1 vccd1 vccd1 _6531_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3739_ _7556_/Q _3739_/B vssd1 vssd1 vccd1 vccd1 _3742_/C sky130_fd_sc_hd__nor2_1
X_6458_ _6521_/B _6521_/C _6629_/A vssd1 vssd1 vccd1 vccd1 _6461_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ hold267/X _4719_/Y _5409_/S vssd1 vssd1 vccd1 vccd1 _5409_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6389_ input32/X _6388_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6389_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7049__A2 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4329__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4853__A _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5299__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4510__A3 _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6962__B _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5223__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6971__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5760_ _5769_/A _5760_/B vssd1 vssd1 vccd1 vccd1 _5761_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4360_/B _4711_/B vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3785__A1 _7543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3785__B2 _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5691_ _5691_/A vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__inv_2
X_7430_ _7430_/CLK _7430_/D vssd1 vssd1 vccd1 vccd1 _7430_/Q sky130_fd_sc_hd__dfxtp_1
X_4642_ _7482_/Q _7470_/Q _7462_/Q _7256_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4642_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4573_ _4573_/A vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__inv_2
XFILLER_0_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7361_ _7569_/CLK _7361_/D vssd1 vssd1 vccd1 vccd1 _7361_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7292_ _7372_/CLK _7292_/D vssd1 vssd1 vccd1 vccd1 _7292_/Q sky130_fd_sc_hd__dfxtp_1
X_6312_ _6235_/A _6911_/A _7098_/A _6311_/X vssd1 vssd1 vccd1 vccd1 _6333_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6243_ _6244_/A _6857_/A vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6174_ _3751_/Y _6172_/X _6173_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6174_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout192_A _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5125_ hold541/X _4990_/Y _5129_/S vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5056_ hold261/X _4996_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _7322_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6872__B _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ _4007_/A _4007_/B _6220_/B vssd1 vssd1 vccd1 vccd1 _4007_/X sky130_fd_sc_hd__or3_1
XFILLER_0_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6411__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5958_ _5958_/A _5958_/B vssd1 vssd1 vccd1 vccd1 _5958_/Y sky130_fd_sc_hd__nand2_1
X_4909_ _4351_/A _4351_/B _4986_/S vssd1 vssd1 vccd1 vccd1 _4909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3776__A1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7195__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5889_ _6581_/A _5918_/D _5888_/C vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7559_ _7579_/CLK _7559_/D vssd1 vssd1 vccd1 vccd1 _7559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5150__A0 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit8 split8/A vssd1 vssd1 vccd1 vccd1 split8/X sky130_fd_sc_hd__buf_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__buf_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4583__A _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5453__A1 _5452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5205__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6953__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3862__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7400_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4716__B1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6022__B _6022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5353__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__A _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__A1 _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5589__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer28 _5549_/B vssd1 vssd1 vccd1 vccd1 _5561_/A2 sky130_fd_sc_hd__clkbuf_1
X_6930_ _6290_/B _6290_/C _6872_/A vssd1 vssd1 vccd1 vccd1 _6931_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7197__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6861_ _6862_/B _6874_/C _6860_/X vssd1 vssd1 vccd1 vccd1 _6864_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5812_ _5811_/A _5803_/X _5811_/Y _6311_/A _5810_/X vssd1 vssd1 vccd1 vccd1 _5812_/X
+ sky130_fd_sc_hd__a221o_1
X_6792_ _6864_/A _6795_/B vssd1 vssd1 vccd1 vccd1 _6848_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6944__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6944__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5743_ _5747_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5763_/C sky130_fd_sc_hd__and2_1
XANTENNA__3853__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5674_ _5675_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6213__A _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7413_ _7413_/CLK _7413_/D vssd1 vssd1 vccd1 vccd1 _7413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4625_ _4625_/A _4625_/B _4625_/C vssd1 vssd1 vccd1 vccd1 _4625_/X sky130_fd_sc_hd__or3_1
XFILLER_0_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold511 _5347_/X vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
X_7344_ _7423_/CLK _7344_/D vssd1 vssd1 vccd1 vccd1 _7344_/Q sky130_fd_sc_hd__dfxtp_2
X_4556_ _6793_/A _4555_/X _4700_/B vssd1 vssd1 vccd1 vccd1 _4557_/B sky130_fd_sc_hd__mux2_1
Xhold500 _7523_/Q vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold522 _7415_/Q vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _5233_/X vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _5180_/X vssd1 vssd1 vccd1 vccd1 _7380_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4237__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout205_A _7340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5771__B _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold588 _7394_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _7315_/Q vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _7324_/Q vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _7422_/Q vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
X_7275_ _7379_/CLK _7275_/D vssd1 vssd1 vccd1 vccd1 _7275_/Q sky130_fd_sc_hd__dfxtp_1
X_4487_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4533_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7044__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6226_ input36/X _6225_/B _6225_/Y _6015_/A vssd1 vssd1 vccd1 vccd1 _7553_/D sky130_fd_sc_hd__o211a_1
Xhold599 _7259_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6157_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6157_/Y sky130_fd_sc_hd__nor2_1
X_5108_ _5107_/X _4973_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__mux2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6088_/A vssd1 vssd1 vccd1 vccd1 _6088_/Y sky130_fd_sc_hd__inv_2
X_5039_ hold566/X _5038_/X _5039_/S vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7188__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3997__B2 _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3844__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5665__C _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6163__A2 _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5173__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__A _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7112__A1 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7112__B2 _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput64 _7580_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_12
Xoutput53 _5918_/D vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
Xoutput75 _7524_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XANTENNA__6793__A _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7179__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5348__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5362__A0 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6154__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4410_ _4701_/B _4406_/X _4409_/X vssd1 vssd1 vccd1 vccd1 _4410_/X sky130_fd_sc_hd__o21ba_1
X_5390_ _5389_/X _4637_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7482_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_78_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _7436_/Q _7428_/Q _7412_/Q _7404_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4341_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5083__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7103__A1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4272_ _4407_/A _4879_/S _4272_/C vssd1 vssd1 vccd1 vccd1 _4272_/Y sky130_fd_sc_hd__nand3_1
X_7060_ _6882_/B split4/A vssd1 vssd1 vccd1 vccd1 _7060_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6011_ _6204_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _7502_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6209__A3 _3739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6208__A _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6913_ _6913_/A vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__inv_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout155_A _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6844_ _6844_/A _6844_/B vssd1 vssd1 vccd1 vccd1 _6845_/B sky130_fd_sc_hd__and2_1
XFILLER_0_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6775_ _6822_/A _6774_/Y _6765_/X vssd1 vssd1 vccd1 vccd1 _6775_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _5990_/A _6374_/B vssd1 vssd1 vccd1 vccd1 _6922_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ _6874_/A _6869_/A _6857_/A _6261_/A vssd1 vssd1 vccd1 vccd1 _5727_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4156__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6145__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5782__A _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5657_ _6683_/A _6742_/A _5640_/B _5639_/B vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4608_ _4658_/A _4606_/X _4607_/Y _4930_/S vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__o211a_1
X_5588_ _5589_/B _5589_/C vssd1 vssd1 vccd1 vccd1 _5612_/B sky130_fd_sc_hd__and2_1
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4398__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4251__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 _5307_/X vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
X_7327_ _7446_/CLK _7327_/D vssd1 vssd1 vccd1 vccd1 _7327_/Q sky130_fd_sc_hd__dfxtp_1
Xhold330 _4888_/X vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _7268_/Q vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _7604_/Q _4540_/B vssd1 vssd1 vccd1 vccd1 _4539_/Y sky130_fd_sc_hd__nand2_1
Xhold374 _7403_/Q vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _7277_/Q vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _7482_/Q vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _7274_/Q vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
X_7258_ _7541_/CLK hold71/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_2
X_6209_ _6922_/A _5990_/A _3739_/B _3763_/A vssd1 vssd1 vccd1 vccd1 _6209_/X sky130_fd_sc_hd__a31o_1
X_7189_ hold651/X _4679_/X _7191_/S vssd1 vssd1 vccd1 vccd1 _7189_/X sky130_fd_sc_hd__mux2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5022__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5957__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4861__A _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6908__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5168__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3817__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4072__S _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5592__B1 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__A0 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6136__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6788__A _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4800__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4242__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6300__B _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5895__A1 _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7097__A0 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output49_A _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3910_ _3934_/A _6120_/A vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__nand2_1
X_4890_ _4862_/A _6039_/A _6048_/A vssd1 vssd1 vccd1 vccd1 _4892_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _3839_/X _3840_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3841_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4386__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3808__S1 _7361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6560_ _6673_/A _6561_/B vssd1 vssd1 vccd1 vccd1 _6596_/B sky130_fd_sc_hd__and2_1
X_3772_ _3780_/B _7123_/C _3948_/A vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5511_ _6518_/A _5507_/A _5507_/B _5536_/A vssd1 vssd1 vccd1 vccd1 _5512_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6127__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6491_ _6468_/B _6506_/B _6468_/A vssd1 vssd1 vccd1 vccd1 _6491_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4710__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5442_ _5444_/B _5444_/C _5788_/D vssd1 vssd1 vccd1 vccd1 _5442_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5373_ hold301/X _4719_/Y _5373_/S vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4233__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4324_ _7398_/Q _7390_/Q _7366_/Q _7382_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4324_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7088__B1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7112_ _3716_/Y _7108_/Y _7110_/Y _6913_/A vssd1 vssd1 vccd1 vccd1 _7112_/X sky130_fd_sc_hd__o22a_1
Xfanout106 _5452_/A vssd1 vssd1 vccd1 vccd1 _6869_/A sky130_fd_sc_hd__buf_6
Xfanout117 _6142_/S vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__clkbuf_8
X_7043_ _7034_/X _7042_/X _7043_/S vssd1 vssd1 vccd1 vccd1 _7044_/D sky130_fd_sc_hd__mux2_1
Xfanout128 _7587_/Q vssd1 vssd1 vccd1 vccd1 _6683_/A sky130_fd_sc_hd__clkbuf_4
X_4255_ _7420_/Q _7352_/Q _7344_/Q _7324_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4255_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4946__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout139 _7579_/Q vssd1 vssd1 vccd1 vccd1 _6827_/A sky130_fd_sc_hd__buf_6
X_4186_ _4184_/X _4185_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4186_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6827_ _6827_/A _6891_/A vssd1 vssd1 vccd1 vccd1 _6828_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6758_ _6759_/A _6759_/B split7/A vssd1 vssd1 vccd1 vccd1 _6758_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4129__A1 _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6689_ _6659_/Y _6684_/X _6686_/X _5788_/D vssd1 vssd1 vccd1 vccd1 _6728_/B sky130_fd_sc_hd__o211ai_1
X_5709_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5711_/B sky130_fd_sc_hd__xor2_1
XANTENNA__5326__A0 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4224__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6120__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold171 _7308_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _6207_/X vssd1 vssd1 vccd1 vccd1 _6208_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7079__B1 _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 _7304_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _7295_/Q vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5014__C1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4530__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6311__A _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5361__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3670__A _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ _4122_/D _4033_/X _6023_/S _4067_/C vssd1 vssd1 vccd1 vccd1 _4046_/C sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6981__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5991_ _5990_/A _6415_/A _6415_/B _4029_/Y _4267_/D vssd1 vssd1 vccd1 vccd1 _5991_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3803__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4942_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873_ _4873_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__nor2_1
X_6612_ _6673_/A _6612_/B vssd1 vssd1 vccd1 vccd1 _6617_/B sky130_fd_sc_hd__nor2_1
X_7592_ _7592_/CLK _7592_/D vssd1 vssd1 vccd1 vccd1 _7592_/Q sky130_fd_sc_hd__dfxtp_1
X_3824_ _7372_/Q _7300_/Q _7292_/Q _7284_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3824_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3755_ _6417_/B _4021_/A vssd1 vssd1 vccd1 vccd1 _4267_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6543_ _6484_/B _7090_/B _6542_/X _6534_/Y vssd1 vssd1 vccd1 vccd1 _6544_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3845__A _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6474_ _6474_/A _6486_/A vssd1 vssd1 vccd1 vccd1 _6480_/A sky130_fd_sc_hd__or2_1
X_3686_ _5977_/B _7554_/Q vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__nor2_2
X_5425_ _6683_/B _5818_/B _5438_/A _6875_/A hold78/A vssd1 vssd1 vccd1 vccd1 _5432_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout118_A _6160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5356_ _4685_/X _5355_/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7463_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5287_ hold208/X _4864_/X _5301_/S vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__mux2_1
X_4307_ _4306_/X _4305_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5271__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4238_ _4238_/A vssd1 vssd1 vccd1 vccd1 _5002_/B sky130_fd_sc_hd__inv_2
X_7026_ _6962_/A _6911_/A _7098_/A _7025_/X vssd1 vssd1 vccd1 vccd1 _7044_/B sky130_fd_sc_hd__o211a_1
XANTENNA__6284__A1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6284__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4169_ _7351_/Q _5037_/B vssd1 vssd1 vccd1 vccd1 _4170_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7198__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4047__A0 hold66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3942__A_N _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3739__B _3739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4445__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3755__A _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7544__CLK _7544_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4289__C _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5970__A _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5181__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7597_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_3_5__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6306__A _6338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6983__C1 _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5356__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3665__A _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4761__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5210_ _4996_/X hold589/X _5212_/S vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6190_ hold88/X hold42/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__mux2_1
X_5141_ _5357_/A _5321_/B _7175_/B vssd1 vssd1 vccd1 vccd1 _5158_/S sky130_fd_sc_hd__or3b_4
XANTENNA__5091__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5072_ _5071_/X _4973_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__mux2_1
X_4023_ _6329_/A _4140_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__and3_2
XANTENNA__4372__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4435__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5974_ _6922_/A _5977_/B _5974_/C _5974_/D vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__or4_1
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4925_ _4873_/A _4199_/B _4208_/A vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4856_ _6808_/B _4123_/B _4698_/A _4855_/Y vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__o211ai_1
X_3807_ _7480_/Q _7468_/Q _7460_/Q _7254_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3807_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7575_ _7587_/CLK _7575_/D vssd1 vssd1 vccd1 vccd1 _7575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4787_ _4747_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _5159_/C sky130_fd_sc_hd__and2b_2
X_6526_ _6563_/A _6570_/A vssd1 vssd1 vccd1 vccd1 _6557_/B sky130_fd_sc_hd__nor2_1
X_3738_ input39/X _7559_/Q vssd1 vssd1 vccd1 vccd1 _3739_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3669_ _6802_/B vssd1 vssd1 vccd1 vccd1 _3669_/Y sky130_fd_sc_hd__inv_2
X_6457_ _6629_/A _6521_/B _6521_/C vssd1 vssd1 vccd1 vccd1 _6461_/A sky130_fd_sc_hd__and3_1
X_5408_ _4637_/X _5407_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7490_/D sky130_fd_sc_hd__mux2_1
X_6388_ _6872_/A _6383_/Y _6387_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6388_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5339_ _5357_/A _5393_/B _7175_/B vssd1 vssd1 vccd1 vccd1 _5356_/S sky130_fd_sc_hd__or3b_4
X_7009_ _7009_/A _7009_/B _7009_/C vssd1 vssd1 vccd1 vccd1 _7009_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4853__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6126__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4991__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4743__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5176__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3929__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4709_/X _4708_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__mux2_1
X_5690_ _5665_/X _5677_/A _6516_/A _5788_/D vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__o211a_1
X_4641_ _7282_/Q _7597_/Q _7266_/Q _7490_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4641_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4734__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5086__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4572_ _4572_/A _4625_/A vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_40_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7360_ _7624_/CLK _7360_/D vssd1 vssd1 vccd1 vccd1 _7360_/Q sky130_fd_sc_hd__dfxtp_4
X_7291_ _7379_/CLK _7291_/D vssd1 vssd1 vccd1 vccd1 _7291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6311_ _6311_/A _7230_/A vssd1 vssd1 vccd1 vccd1 _6311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6242_ _7025_/A _6673_/A vssd1 vssd1 vccd1 vccd1 _6242_/X sky130_fd_sc_hd__or2_1
XANTENNA__4593__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6173_ _6173_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__or2_1
X_5124_ _5123_/X _4947_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _7356_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout185_A _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5055_ hold260/X _5015_/X _5057_/S vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4345__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4006_ _4004_/A _4004_/B _3666_/Y _4005_/X vssd1 vssd1 vccd1 vccd1 _4006_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5957_ _6235_/A _6827_/A vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__nand2_2
XANTENNA__4973__A1 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4908_ _4908_/A _4982_/A vssd1 vssd1 vccd1 vccd1 _4908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3776__A2 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _6581_/A _5918_/D _5888_/C vssd1 vssd1 vccd1 vccd1 _5913_/B sky130_fd_sc_hd__and3_1
XFILLER_0_105_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839_ hold493/X _4629_/X _4843_/S vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7558_ _7599_/CLK _7558_/D vssd1 vssd1 vccd1 vccd1 _7558_/Q sky130_fd_sc_hd__dfxtp_4
X_7489_ _7489_/CLK _7489_/D vssd1 vssd1 vccd1 vccd1 _7489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6509_ _6467_/B _6509_/B _6521_/A vssd1 vssd1 vccd1 vccd1 _6513_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xsplit9 split9/A vssd1 vssd1 vccd1 vccd1 split9/X sky130_fd_sc_hd__buf_4
XANTENNA__4336__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4803__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6953__A2 hold610/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3943__A _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_wb_clk_i _7544_/CLK vssd1 vssd1 vccd1 vccd1 _7534_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__A2 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4327__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer29 split1/A vssd1 vssd1 vccd1 vccd1 _5555_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6860_ _6860_/A _6860_/B vssd1 vssd1 vccd1 vccd1 _6860_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5811_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5811_/Y sky130_fd_sc_hd__nor2_2
X_6791_ _6795_/B vssd1 vssd1 vccd1 vccd1 _6791_/Y sky130_fd_sc_hd__inv_2
X_5742_ _5758_/A _5742_/B vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5673_ _5701_/B _5673_/B vssd1 vssd1 vccd1 vccd1 _5675_/B sky130_fd_sc_hd__nor2_1
X_7412_ _7430_/CLK _7412_/D vssd1 vssd1 vccd1 vccd1 _7412_/Q sky130_fd_sc_hd__dfxtp_1
X_4624_ _4624_/A _4624_/B vssd1 vssd1 vccd1 vccd1 _4625_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5380__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4555_ _4554_/Y _4552_/Y _4701_/B vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__mux2_1
X_7343_ _7569_/CLK _7343_/D vssd1 vssd1 vccd1 vccd1 _7343_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold501 _6183_/X vssd1 vssd1 vccd1 vccd1 _7523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _7251_/Q vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _7460_/Q vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _7464_/Q vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _7408_/Q vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5771__C _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold578 _7300_/Q vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 _5039_/X vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _5061_/X vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ _7306_/CLK _7274_/D vssd1 vssd1 vccd1 vccd1 _7274_/Q sky130_fd_sc_hd__dfxtp_1
X_4486_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__or2_1
Xhold589 _5209_/X vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4566__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6225_ _6225_/A _6225_/B vssd1 vssd1 vccd1 vccd1 _6225_/Y sky130_fd_sc_hd__nand2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _3702_/Y _4649_/Y _6155_/X _6022_/B _6157_/B vssd1 vssd1 vccd1 vccd1 _6156_/X
+ sky130_fd_sc_hd__o221a_1
X_5107_ hold629/X _4990_/Y _5111_/S vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__mux2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _5026_/B _6089_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6088_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5038_ _4529_/S _4170_/B _5037_/X _5036_/X vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__o31a_4
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3997__A2 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5199__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6989_ _6989_/A _6989_/B vssd1 vssd1 vccd1 vccd1 _6989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6123__B _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5665__D _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5371__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput65 _7581_/Q vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_12
XANTENNA__5123__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 _6532_/A vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput76 _7525_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XFILLER_0_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6387__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5364__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3673__A _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ _4474_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4271_ _4271_/A _5027_/A vssd1 vssd1 vccd1 vccd1 _4272_/C sky130_fd_sc_hd__nand2_1
X_6010_ _6191_/B _6190_/S _3758_/Y vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__6195__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6090__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6912_ _3712_/B _7123_/C _6313_/X _6911_/Y vssd1 vssd1 vccd1 vccd1 _6913_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6843_ _6844_/A _6844_/B vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6774_ _6823_/B _6831_/B vssd1 vssd1 vccd1 vccd1 _6774_/Y sky130_fd_sc_hd__nor2_2
X_3986_ _5988_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _6374_/B sky130_fd_sc_hd__or2_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5725_ _6802_/A _6799_/A vssd1 vssd1 vccd1 vccd1 _7009_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5656_ _6581_/A _6518_/A vssd1 vssd1 vccd1 vccd1 _5659_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5353__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4607_ _6673_/A _4658_/A vssd1 vssd1 vccd1 vccd1 _4607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5782__B _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold320 _7316_/Q vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5274__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5587_ _6710_/A _5591_/B _5587_/C _5587_/D vssd1 vssd1 vccd1 vccd1 _5589_/C sky130_fd_sc_hd__or4_4
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold331 _7310_/Q vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _4753_/X vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _7287_/Q vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ _4685_/A _4538_/B vssd1 vssd1 vccd1 vccd1 _4538_/X sky130_fd_sc_hd__or2_4
X_7326_ _7453_/CLK _7326_/D vssd1 vssd1 vccd1 vccd1 _7326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold375 _5229_/X vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _7276_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
X_7257_ _7596_/CLK _7257_/D vssd1 vssd1 vccd1 vccd1 _7257_/Q sky130_fd_sc_hd__dfxtp_1
Xhold364 _7490_/Q vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _7374_/Q _7302_/Q _7294_/Q _7286_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4469_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5105__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold397 _7396_/Q vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _6218_/A _6208_/B vssd1 vssd1 vccd1 vccd1 _7538_/D sky130_fd_sc_hd__nand2_1
X_7188_ _7187_/X _4589_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7605_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4845__C _4846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6139_ _6139_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6139_/Y sky130_fd_sc_hd__nor2_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6081__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5813__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5957__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6908__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5592__A1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5184__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4589__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5895__A2 _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7097__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4528__S _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6072__A2 _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5359__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3668__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _7424_/Q _7356_/Q _7348_/Q _7328_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3840_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6044__A _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3771_ _3780_/B _7123_/C _3948_/A vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5510_ _7494_/Q _6808_/B vssd1 vssd1 vccd1 vccd1 _5536_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6490_ _6754_/A _6532_/B vssd1 vssd1 vccd1 vccd1 _6490_/X sky130_fd_sc_hd__and2_1
XANTENNA__5094__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4499__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5335__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5441_ _6875_/A _5441_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__and2_1
X_5372_ _4637_/X _5371_/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7470_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6210__C _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4323_ _7438_/Q _7430_/Q _7414_/Q _7406_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4323_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7111_ _6910_/A _6309_/B _7109_/X _3775_/Y _6738_/A vssd1 vssd1 vccd1 vccd1 _7111_/X
+ sky130_fd_sc_hd__o32a_1
Xfanout129 _6962_/A vssd1 vssd1 vccd1 vccd1 _6690_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7042_ _5879_/A _7038_/X _7039_/Y _7041_/Y _6989_/A vssd1 vssd1 vccd1 vccd1 _7042_/X
+ sky130_fd_sc_hd__a32o_1
Xfanout107 _5504_/A vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__buf_8
Xfanout118 _6160_/S vssd1 vssd1 vccd1 vccd1 _6142_/S sky130_fd_sc_hd__buf_8
X_4254_ _7316_/Q _7332_/Q _7308_/Q _7444_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4254_/X sky130_fd_sc_hd__mux4_1
X_4185_ _7421_/Q _7353_/Q _7345_/Q _7325_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4185_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6063__A2 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4074__A1 hold524/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5269__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6826_ _6827_/A _6891_/A vssd1 vssd1 vccd1 vccd1 _6836_/B sky130_fd_sc_hd__or2_1
XFILLER_0_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6757_ _6675_/X _6751_/B _6706_/X _6668_/X vssd1 vssd1 vccd1 vccd1 _6759_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4901__S _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5708_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5834_/A sky130_fd_sc_hd__nand2_1
X_3969_ _6920_/A _4267_/C vssd1 vssd1 vccd1 vccd1 _5974_/D sky130_fd_sc_hd__nand2_1
X_6688_ _6659_/Y _6685_/Y _6682_/X _6629_/A vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5639_ _5639_/A _5639_/B vssd1 vssd1 vccd1 vccd1 _5640_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7309_ _7446_/CLK _7309_/D vssd1 vssd1 vccd1 vccd1 _7309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold150 _6007_/Y vssd1 vssd1 vccd1 vccd1 _7500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _7521_/Q vssd1 vssd1 vccd1 vccd1 _6176_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _4865_/X vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _7303_/Q vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _4815_/X vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout80_A _4144_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold644_A _7590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6054__A2 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5179__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7003__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7003__B2 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4811__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6799__A _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5317__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6311__B _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4112__A _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output61_A hold70/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6045__A2 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7242__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5990_ _5990_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6925_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5089__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3803__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4941_ _4971_/B _4941_/B vssd1 vssd1 vccd1 vccd1 _4946_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4872_ _7344_/Q _4872_/B vssd1 vssd1 vccd1 vccd1 _4872_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3823_ _3821_/X _3822_/X _3915_/A vssd1 vssd1 vccd1 vccd1 _3823_/X sky130_fd_sc_hd__mux2_1
X_6611_ _6611_/A _6611_/B vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__nor2_1
X_7591_ _7592_/CLK _7591_/D vssd1 vssd1 vccd1 vccd1 _7591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4721__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7446_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6542_ _6535_/A _6534_/B _7090_/B vssd1 vssd1 vccd1 vccd1 _6542_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3754_ _6216_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__or2_1
XANTENNA__5308__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6473_ _6485_/B _6485_/C _6485_/D _6485_/A vssd1 vssd1 vccd1 vccd1 _6486_/A sky130_fd_sc_hd__a31oi_1
X_3685_ _3759_/A _3685_/B vssd1 vssd1 vccd1 vccd1 _3685_/Y sky130_fd_sc_hd__nand2_1
X_5424_ _6875_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _5428_/B sky130_fd_sc_hd__or2_4
XANTENNA__4022__A _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5355_ hold461/X _4719_/Y _5355_/S vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3861__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5286_ _7151_/B _7194_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5301_/S sky130_fd_sc_hd__and3_4
X_4306_ _7424_/Q _7356_/Q _7348_/Q _7328_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4306_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4237_ _4689_/A _4235_/X _4236_/Y _4232_/Y vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__a2bb2o_2
X_7025_ _7025_/A _7230_/A vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__or2_1
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_4168_ _7350_/Q _4997_/B vssd1 vssd1 vccd1 vccd1 _5037_/B sky130_fd_sc_hd__or2_2
XFILLER_0_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6036__A2 _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5788__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5244__A0 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4099_ _6066_/A _4917_/A vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__or2_1
XANTENNA__4047__A1 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6809_ _6809_/A vssd1 vssd1 vccd1 vccd1 _6865_/B sky130_fd_sc_hd__inv_2
XANTENNA__4631__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3755__B _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7224__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4806__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6983__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4107__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4994__C1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3892__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3946__A _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5372__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5140_ input34/X _6225_/B _5139_/Y _6373_/A vssd1 vssd1 vccd1 vccd1 _7363_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ hold564/X _4990_/Y _5075_/S vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4277__A1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4022_ _5990_/A _4039_/C vssd1 vssd1 vccd1 vccd1 _4290_/D sky130_fd_sc_hd__nand2_4
XFILLER_0_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4372__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7215__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5973_ _3656_/A wire79/X _5972_/X _6218_/A vssd1 vssd1 vccd1 vccd1 _5973_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4924_ _4955_/A _4974_/B _4923_/Y vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3883__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4855_ _4999_/B _4269_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4855_/Y sky130_fd_sc_hd__o21ai_1
X_4786_ _4785_/X _4685_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7283_/D sky130_fd_sc_hd__mux2_1
X_3806_ _3931_/S _3806_/B vssd1 vssd1 vccd1 vccd1 _3806_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4451__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7574_ _7587_/CLK _7574_/D vssd1 vssd1 vccd1 vccd1 _7574_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__6232__A _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6525_ _6575_/A _6569_/B _6569_/C vssd1 vssd1 vccd1 vccd1 _6570_/A sky130_fd_sc_hd__a21o_1
X_3737_ _7473_/Q _4267_/C _3970_/B hold56/X _3693_/Y vssd1 vssd1 vccd1 vccd1 hold57/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3668_ _4689_/A vssd1 vssd1 vccd1 vccd1 _3668_/Y sky130_fd_sc_hd__inv_8
X_6456_ _5571_/X _6430_/A _5626_/X _5604_/A vssd1 vssd1 vccd1 vccd1 _6521_/C sky130_fd_sc_hd__o211ai_2
X_5407_ hold364/X _4679_/X _5409_/S vssd1 vssd1 vccd1 vccd1 _5407_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5282__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6387_ hold128/X _6415_/A _6356_/B hold524/X vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__a22o_1
X_5338_ _5022_/X hold552/X _5338_/S vssd1 vssd1 vccd1 vccd1 _7451_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5269_ hold487/X _4864_/X _5283_/S vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4268__A1 _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7008_ _7009_/B _7008_/B vssd1 vssd1 vccd1 vccd1 _7008_/X sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__7206__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3779__B1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3766__A _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5192__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3929__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5208__A0 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6956__B1 _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5367__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4481__A2_N _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _4638_/X _4639_/Y _4529_/S vssd1 vssd1 vccd1 vccd1 _4640_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3676__A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4571_ _4672_/B _6135_/B vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6310_ _6236_/A _6309_/Y _6234_/Y vssd1 vssd1 vccd1 vccd1 _6310_/Y sky130_fd_sc_hd__a21oi_1
X_7290_ _7306_/CLK _7290_/D vssd1 vssd1 vccd1 vccd1 _7290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6241_ _6273_/A _6673_/A vssd1 vssd1 vccd1 vccd1 _7092_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4300__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6172_ hold72/X hold50/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5695__B1 _6338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4593__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5123_ hold210/X _4964_/X _5129_/S vssd1 vssd1 vccd1 vccd1 _5123_/X sky130_fd_sc_hd__mux2_1
X_5054_ _5053_/X _4973_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4345__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4005_ _7542_/Q input20/X _3666_/A _4004_/Y _7540_/Q vssd1 vssd1 vccd1 vccd1 _4005_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout178_A _7453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3856__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _5956_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5960_/A sky130_fd_sc_hd__and2_1
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4907_ _5008_/A _4901_/X _4906_/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__a211o_1
X_5887_ _5887_/A _5913_/A vssd1 vssd1 vccd1 vccd1 _5888_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4838_ _4837_/X _4538_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7304_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5277__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4281__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4769_ _7211_/B _7150_/B _5375_/C vssd1 vssd1 vccd1 vccd1 _4786_/S sky130_fd_sc_hd__and3_4
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7557_ _7557_/CLK _7557_/D vssd1 vssd1 vccd1 vccd1 _7557_/Q sky130_fd_sc_hd__dfxtp_4
X_7488_ _7598_/CLK _7488_/D vssd1 vssd1 vccd1 vccd1 _7488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6508_ _6508_/A _6508_/B vssd1 vssd1 vccd1 vccd1 _6508_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6439_ _6438_/X _6437_/Y _6463_/S _5580_/B vssd1 vssd1 vccd1 vccd1 _6476_/B sky130_fd_sc_hd__o2bb2a_2
XANTENNA__4489__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4336__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5989__A1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6938__B1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3847__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5187__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4091__S _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3943__B _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7451_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4327__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer19 split1/A vssd1 vssd1 vccd1 vccd1 _5541_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5886__A _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5810_ _5810_/A _5810_/B _5810_/C _5810_/D vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__or4_4
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6790_ _6732_/B _6789_/Y _6790_/S vssd1 vssd1 vccd1 vccd1 _6795_/B sky130_fd_sc_hd__mux2_4
XANTENNA__6481__S _6481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _5758_/A _5742_/B vssd1 vssd1 vccd1 vccd1 _5747_/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7411_ _7443_/CLK _7411_/D vssd1 vssd1 vccd1 vccd1 _7411_/Q sky130_fd_sc_hd__dfxtp_1
X_5672_ _6738_/A _6673_/A _5669_/Y _5701_/A vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__o22a_1
X_4623_ _4672_/B _6144_/B vssd1 vssd1 vccd1 vccd1 _4624_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 _7366_/Q vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
X_4554_ _4554_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4554_/Y sky130_fd_sc_hd__xnor2_1
X_7342_ _7569_/CLK _7342_/D vssd1 vssd1 vccd1 vccd1 _7342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold535 _7411_/Q vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _5241_/X vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
X_7273_ _7621_/CLK _7273_/D vssd1 vssd1 vccd1 vccd1 _7273_/Q sky130_fd_sc_hd__dfxtp_1
Xhold524 _7569_/Q vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4949__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4485_ _4443_/X hold497/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7252_/D sky130_fd_sc_hd__mux2_1
Xhold546 _5359_/X vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _4829_/X vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _7334_/Q vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _7359_/Q vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ input35/X _6225_/B _6223_/Y _6373_/A vssd1 vssd1 vccd1 vccd1 _7552_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4030__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5771__D _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4566__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6025_/Y _6152_/Y _6154_/X vssd1 vssd1 vccd1 vccd1 _6155_/X sky130_fd_sc_hd__o21a_1
X_5106_ _5105_/X _4947_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _7348_/D sky130_fd_sc_hd__mux2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6085_/X hold40/X _6086_/S vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__mux2_1
X_5037_ _5037_/A _5037_/B vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__and2_1
XFILLER_0_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6396__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _6988_/A _6988_/B vssd1 vssd1 vccd1 vccd1 _6988_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5939_ _7123_/A _6827_/A vssd1 vssd1 vccd1 vccd1 _5940_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7609_ _7617_/CLK _7609_/D vssd1 vssd1 vccd1 vccd1 _7609_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4254__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3763__B _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput66 hold94/A vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_12
Xoutput55 _6710_/A vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4882__A1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4634__A1 _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4814__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3938__B _6084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6387__B2 hold524/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4115__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4270_ _5024_/S _4271_/A vssd1 vssd1 vccd1 vccd1 _4270_/X sky130_fd_sc_hd__or2_1
XANTENNA__5380__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6911_ _6911_/A _6911_/B vssd1 vssd1 vccd1 vccd1 _6911_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6842_ _6784_/B _6841_/X _6891_/B vssd1 vssd1 vccd1 vccd1 _6844_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5050__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3985_ _5980_/B _4081_/A _3985_/C _3980_/X vssd1 vssd1 vccd1 vccd1 _3985_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_9_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6773_ _6773_/A _6773_/B vssd1 vssd1 vccd1 vccd1 _6831_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4025__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5724_ _6808_/A _5788_/B _6864_/A _6793_/A vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__and4_1
XFILLER_0_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5655_ _5739_/A _5739_/B vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4606_ _4603_/Y _4605_/X _4701_/B vssd1 vssd1 vccd1 vccd1 _4606_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5782__C _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6240__A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold310 _5051_/X vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
X_7325_ _7453_/CLK _7325_/D vssd1 vssd1 vccd1 vccd1 _7325_/Q sky130_fd_sc_hd__dfxtp_1
X_5586_ _6840_/A _5586_/A2 _5534_/A vssd1 vssd1 vccd1 vccd1 _5589_/B sky130_fd_sc_hd__a21o_1
Xhold332 _7336_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _5043_/X vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _4797_/X vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _3922_/X _4106_/X _4536_/Y _4535_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _4538_/B
+ sky130_fd_sc_hd__o32a_1
Xhold387 _4771_/X vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _7483_/Q vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
X_7256_ _7481_/CLK _7256_/D vssd1 vssd1 vccd1 vccd1 _7256_/Q sky130_fd_sc_hd__dfxtp_1
X_4468_ _4467_/X _4667_/B vssd1 vssd1 vccd1 vccd1 _4468_/Y sky130_fd_sc_hd__nand2b_1
Xhold354 _7444_/Q vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _7358_/Q vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold398 _5215_/X vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
X_7187_ hold620/X _4629_/X _7191_/S vssd1 vssd1 vccd1 vccd1 _7187_/X sky130_fd_sc_hd__mux2_1
X_6207_ _3644_/Y _3645_/Y _6207_/S vssd1 vssd1 vccd1 vccd1 _6207_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5290__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4399_ _7373_/Q _7301_/Q _7293_/Q _7285_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4399_/X sky130_fd_sc_hd__mux4_1
X_6138_ _3702_/Y _4553_/B _6137_/X _6375_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6138_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6069_ _4977_/B _6071_/B _6911_/A vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6908__A3 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4809__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4855__A1 _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4544__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4466__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3770_ _3770_/A _3770_/B vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__or2_1
XFILLER_0_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _5444_/B _5444_/C vssd1 vssd1 vccd1 vccd1 _5441_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5371_ hold305/X _4679_/X _5373_/S vssd1 vssd1 vccd1 vccd1 _5371_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _4474_/A _6053_/B vssd1 vssd1 vccd1 vccd1 _4353_/B sky130_fd_sc_hd__nand2_1
X_7110_ _7110_/A _7110_/B vssd1 vssd1 vccd1 vccd1 _7110_/Y sky130_fd_sc_hd__xnor2_1
X_4253_ _4401_/S _4253_/B vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__or2_1
XANTENNA__5099__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 _3670_/Y vssd1 vssd1 vccd1 vccd1 _6875_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7041_ _7041_/A _7041_/B vssd1 vssd1 vccd1 vccd1 _7041_/Y sky130_fd_sc_hd__nor2_1
Xfanout119 _7090_/A vssd1 vssd1 vccd1 vccd1 _7043_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4184_ _7317_/Q _7333_/Q _7309_/Q _7445_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4184_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5271__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6235__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5023__A1 _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6825_ _6771_/B _6775_/Y _6824_/X vssd1 vssd1 vccd1 vccd1 _6891_/A sky130_fd_sc_hd__a21oi_1
X_6756_ _6756_/A _6756_/B vssd1 vssd1 vccd1 vccd1 _6759_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ _6345_/A _5990_/A _6331_/A _3967_/X vssd1 vssd1 vccd1 vccd1 _7473_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _5821_/B _5707_/B vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3899_ _3939_/A _6093_/A vssd1 vssd1 vccd1 vccd1 _3937_/A sky130_fd_sc_hd__nand2_1
X_6687_ _6659_/Y _6685_/Y _6682_/X vssd1 vssd1 vccd1 vccd1 _6687_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5638_ _6690_/A _6802_/A _6637_/A _6702_/A vssd1 vssd1 vccd1 vccd1 _5639_/B sky130_fd_sc_hd__and4_1
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5569_ _6431_/A _5570_/C vssd1 vssd1 vccd1 vccd1 _5571_/B sky130_fd_sc_hd__or2_1
X_7308_ _7448_/CLK _7308_/D vssd1 vssd1 vccd1 vccd1 _7308_/Q sky130_fd_sc_hd__dfxtp_1
Xhold151 _7535_/Q vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _7566_/Q vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _6177_/X vssd1 vssd1 vccd1 vccd1 _7521_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _7338_/Q vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _7612_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _4835_/X vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4837__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7239_ hold111/X hold60/X _7241_/S vssd1 vssd1 vccd1 vccd1 _7239_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5262__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold637_A _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6039__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4687__S0 _7452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5253__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _6066_/A _4940_/B vssd1 vssd1 vccd1 vccd1 _4941_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4461__C1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4871_ _4083_/X _4869_/X _4870_/Y vssd1 vssd1 vccd1 vccd1 _4871_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA_split26_A _6445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3822_ _7476_/Q _7464_/Q _7456_/Q _7250_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3822_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6610_ _6568_/B _6607_/X split9/X vssd1 vssd1 vccd1 vccd1 _6611_/B sky130_fd_sc_hd__mux2_1
X_7590_ _7590_/CLK _7590_/D vssd1 vssd1 vccd1 vccd1 _7590_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5894__A _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6348__A4 _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6541_ _6583_/B _6583_/C vssd1 vssd1 vccd1 vccd1 _7090_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _6216_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _6207_/S sky130_fd_sc_hd__nor2_8
XFILLER_0_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6472_ _6507_/B _6466_/B _6506_/B _6498_/B _6468_/A vssd1 vssd1 vccd1 vccd1 _6485_/D
+ sky130_fd_sc_hd__a2111o_1
X_3684_ _3759_/A _3685_/B vssd1 vssd1 vccd1 vccd1 _3684_/X sky130_fd_sc_hd__and2_1
X_5423_ _6875_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__nor2_1
X_5354_ _4637_/X _5353_/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7462_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _7320_/Q _7336_/Q _7312_/Q _7448_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4305_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5285_ _7150_/B _7193_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5302_/S sky130_fd_sc_hd__and3_4
XANTENNA__4819__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4236_ _4401_/S _4230_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4236_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7024_ _7040_/A _7040_/B _6989_/B _6910_/A vssd1 vssd1 vccd1 vccd1 _7024_/X sky130_fd_sc_hd__a31o_1
X_4167_ _7348_/Q _7349_/Q _4948_/B vssd1 vssd1 vccd1 vccd1 _4997_/B sky130_fd_sc_hd__or3_1
X_4098_ _6057_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6992__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6992__B2 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6808_ _6808_/A _6808_/B vssd1 vssd1 vccd1 vccd1 _6809_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold120_A _7543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6739_ _6875_/A _6739_/B vssd1 vssd1 vccd1 vccd1 _6740_/B sky130_fd_sc_hd__or2_4
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5180__A0 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4359__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__B _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4669__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5786__A2 _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6983__B2 _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3892__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4822__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7608_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout90 _4290_/X vssd1 vssd1 vccd1 vccd1 _4672_/B sky130_fd_sc_hd__buf_4
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7160__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5070_ hold253/X _4947_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _7328_/D sky130_fd_sc_hd__mux2_1
X_4021_ _4021_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4279_/C sky130_fd_sc_hd__nor2_8
XANTENNA__5226__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _6516_/A _5811_/Y _5970_/X _5971_/Y _5810_/X vssd1 vssd1 vccd1 vccd1 _5972_/X
+ sky130_fd_sc_hd__a221o_1
X_4923_ _4902_/B _4900_/B _4209_/B vssd1 vssd1 vccd1 vccd1 _4923_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4732__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3883__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4854_ _4953_/B _4853_/Y _4930_/S vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_7_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6513__A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _7280_/Q _7595_/Q _7264_/Q _7488_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3806_/B sky130_fd_sc_hd__mux4_1
X_4785_ hold379/X _4719_/Y _4785_/S vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__mux2_1
X_7573_ _7577_/CLK _7573_/D vssd1 vssd1 vccd1 vccd1 _7573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6524_ _6871_/A _6524_/B vssd1 vssd1 vccd1 vccd1 _6569_/C sky130_fd_sc_hd__xnor2_1
X_3736_ _6015_/A _4009_/A _4039_/A vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__and3_1
X_3667_ _4688_/S vssd1 vssd1 vccd1 vccd1 _3667_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4968__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6455_ _5621_/Y _5622_/X _5626_/X _5608_/A vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__a31o_1
X_5406_ _4589_/X hold436/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7489_/D sky130_fd_sc_hd__mux2_1
X_6386_ _6385_/X hold637/X _6414_/S vssd1 vssd1 vccd1 vccd1 _6386_/X sky130_fd_sc_hd__mux2_1
X_5337_ hold551/X _5038_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5337_/X sky130_fd_sc_hd__mux2_1
X_5268_ _7212_/C _5376_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5283_/S sky130_fd_sc_hd__and3_4
X_4219_ _4955_/A _4219_/B vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__nand2_1
X_7007_ _6253_/Y _6977_/B _6264_/A vssd1 vssd1 vccd1 vccd1 _7008_/B sky130_fd_sc_hd__a21oi_1
X_5199_ hold537/X _4887_/X _5211_/S vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5217__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3779__A1 _7559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3951__A1 _7546_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3782__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3703__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4817__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6405__A0 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4118__A _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _4672_/B _6135_/B vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5144__A0 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5383__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6240_ _7025_/A _6673_/A vssd1 vssd1 vccd1 vccd1 _6240_/X sky130_fd_sc_hd__and2_1
XFILLER_0_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5695__A1 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6171_ _3751_/Y _6169_/X _6170_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6171_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5122_ _5121_/X _4921_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _7355_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5447__A1 _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5053_ hold250/X _4990_/Y _5057_/S vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5412__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _4004_/A _4004_/B vssd1 vssd1 vccd1 vccd1 _4004_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6947__A1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5955_ _5955_/A _5955_/B _5955_/C _5955_/D vssd1 vssd1 vccd1 vccd1 _5955_/X sky130_fd_sc_hd__or4_1
XANTENNA__3856__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4906_ _4976_/B _4904_/X _4905_/Y _4930_/S vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6243__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5886_ _6273_/A _6683_/A _6771_/A _6773_/A vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__and4_1
X_4837_ hold193/X _4580_/X _4843_/S vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4281__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4768_ _4767_/X _4685_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7275_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7556_ _7557_/CLK _7556_/D vssd1 vssd1 vccd1 vccd1 _7556_/Q sky130_fd_sc_hd__dfxtp_4
X_7487_ _7487_/CLK _7487_/D vssd1 vssd1 vccd1 vccd1 _7487_/Q sky130_fd_sc_hd__dfxtp_1
X_4699_ _4699_/A _4699_/B vssd1 vssd1 vccd1 vccd1 _4699_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4698__A _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6389__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7124__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6507_ _6461_/A _6507_/B vssd1 vssd1 vccd1 vccd1 _6508_/B sky130_fd_sc_hd__nand2b_1
X_3719_ _4037_/A _5805_/A _6421_/B vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__and3_4
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6438_ _6437_/A _6437_/B _6463_/S vssd1 vssd1 vccd1 vccd1 _6438_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4489__A2 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5686__A1 _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6369_ _6373_/A _6369_/B vssd1 vssd1 vccd1 vccd1 _7565_/D sky130_fd_sc_hd__and2_1
XANTENNA__3792__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__clkbuf_2
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__buf_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3777__A _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3847__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6153__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5374__A0 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7115__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3943__C _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4885__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A1 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6328__A _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7150__C _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4652__A2 _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7599_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6929__A1 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5378__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4790__B _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5886__B _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5740_ _5740_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5742_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7410_ _7443_/CLK _7410_/D vssd1 vssd1 vccd1 vccd1 _7410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5671_ _5701_/A _6718_/A _6802_/A _5671_/D vssd1 vssd1 vccd1 vccd1 _5701_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4622_ _4672_/B _6144_/B vssd1 vssd1 vccd1 vccd1 _4624_/A sky130_fd_sc_hd__and2_1
XFILLER_0_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6583__A_N _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7341_ _7453_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 _7341_/Q sky130_fd_sc_hd__dfxtp_4
X_4553_ _4554_/A _4553_/B vssd1 vssd1 vccd1 vccd1 _4553_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7106__A1 _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 _5247_/X vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 _5147_/X vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ hold496/X _4483_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__mux2_1
X_7272_ _7306_/CLK _7272_/D vssd1 vssd1 vccd1 vccd1 _7272_/Q sky130_fd_sc_hd__dfxtp_1
Xhold525 _4074_/X vssd1 vssd1 vccd1 vccd1 _7453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _7474_/Q vssd1 vssd1 vccd1 vccd1 _4001_/D sky130_fd_sc_hd__buf_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold547 _7371_/Q vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _5129_/X vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _7570_/Q vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__clkbuf_2
X_6223_ _6223_/A _6225_/B vssd1 vssd1 vccd1 vccd1 _6223_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5668__A1 _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4030__B _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _7606_/Q _6153_/A _6153_/Y _3975_/X vssd1 vssd1 vccd1 vccd1 _6154_/X sky130_fd_sc_hd__a211o_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout190_A _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5105_ _4948_/A _4964_/X _5111_/S vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__mux2_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6427_/B _6083_/X _6084_/Y _5002_/B _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6085_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6238__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5036_ _4162_/B _5031_/X _5035_/X _4989_/A vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4628__C1 _4144_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5288__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6987_ _6935_/A _6926_/Y _6985_/Y _6986_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7585_/D
+ sky130_fd_sc_hd__o221a_1
X_5938_ _6235_/A _6844_/A vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5356__A0 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5869_ _5869_/A _5869_/B _5869_/C vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__nand3_1
X_7608_ _7608_/CLK _7608_/D vssd1 vssd1 vccd1 vccd1 _7608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4254__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6420__B _6427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7539_ _7541_/CLK _7539_/D vssd1 vssd1 vccd1 vccd1 _7539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4221__A _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3843__A1_N _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput45 _7540_/Q vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_12
Xoutput67 _7556_/Q vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_12
Xoutput56 _4003_/X vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
XANTENNA__6148__A _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4634__A2 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4190__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3842__B1 _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5198__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4115__B _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4830__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6611__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4858__C1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_4_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5822__A1 _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4181__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6910_ _6910_/A _6932_/C _6910_/C vssd1 vssd1 vccd1 vccd1 _6910_/X sky130_fd_sc_hd__and3_1
XANTENNA__5822__B2 _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6841_ _6841_/A _6841_/B vssd1 vssd1 vccd1 vccd1 _6841_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5035__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6772_ _6822_/B vssd1 vssd1 vccd1 vccd1 _6823_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3984_ _6225_/A _4044_/A vssd1 vssd1 vccd1 vccd1 _4031_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_45_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5723_ _5723_/A _5723_/B vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__and2_1
XANTENNA__4740__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5338__A0 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5654_ _5654_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5739_/B sky130_fd_sc_hd__and2_1
XFILLER_0_60_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4605_ _4698_/A _4698_/B _4604_/Y vssd1 vssd1 vccd1 vccd1 _4605_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5782__D _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6240__B _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5889__A1 _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold311 _7593_/Q vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 _5057_/X vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
X_7324_ _7453_/CLK _7324_/D vssd1 vssd1 vccd1 vccd1 _7324_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4561__A1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5585_ _5585_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5587_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold344 _7263_/Q vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _5087_/X vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 _7379_/Q vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ _6139_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _4536_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout203_A _7340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4467_ _4465_/X _4466_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4467_/X sky130_fd_sc_hd__mux2_1
X_7255_ _7618_/CLK _7255_/D vssd1 vssd1 vccd1 vccd1 _7255_/Q sky130_fd_sc_hd__dfxtp_1
Xhold355 _5323_/X vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _7325_/Q vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3880__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold366 _7619_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4976__A _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold399 _7436_/Q vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_4398_ _4689_/A _4398_/B vssd1 vssd1 vccd1 vccd1 _4398_/X sky130_fd_sc_hd__and2_1
Xhold388 _7352_/Q vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
X_7186_ _7185_/X _4538_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7604_/D sky130_fd_sc_hd__mux2_1
X_6206_ _7244_/A _6206_/B vssd1 vssd1 vccd1 vccd1 _7537_/D sky130_fd_sc_hd__or2_1
X_6137_ _6025_/Y _6134_/Y _6136_/X vssd1 vssd1 vccd1 vccd1 _6137_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4864__A2 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6068_ _6067_/X hold44/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__mux2_1
XANTENNA__4172__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5019_ _5019_/A _5019_/B vssd1 vssd1 vccd1 vccd1 _5019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_as1802_214 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_214/HI io_out[25] sky130_fd_sc_hd__conb_1
XFILLER_0_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7201__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4466__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4791__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3965__A _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5370_ _4589_/X hold190/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7469_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5391__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4321_ _4474_/A _6053_/B vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__and2_1
X_4252_ _7396_/Q _7388_/Q _7364_/Q _7380_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4253_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7040_ _7040_/A _7040_/B _7040_/C vssd1 vssd1 vccd1 vccd1 _7041_/B sky130_fd_sc_hd__and3_1
Xfanout109 _3670_/Y vssd1 vssd1 vccd1 vccd1 _6629_/A sky130_fd_sc_hd__buf_2
X_4183_ _7437_/Q _7429_/Q _7413_/Q _7405_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4183_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4735__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6516__A _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6235__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout153_A _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6824_ _6832_/A _6831_/C _6824_/C vssd1 vssd1 vccd1 vccd1 _6824_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6755_ _6773_/A _6773_/B _6831_/A vssd1 vssd1 vccd1 vccd1 _6755_/Y sky130_fd_sc_hd__o21ai_1
X_3967_ _5978_/A _3693_/Y _3966_/X _6920_/A vssd1 vssd1 vccd1 vccd1 _3967_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4782__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6251__A _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5706_ _6691_/A _6673_/A _5703_/Y _5821_/A vssd1 vssd1 vccd1 vccd1 _5707_/B sky130_fd_sc_hd__o22a_1
X_3898_ _3665_/Y _3897_/X _3894_/X vssd1 vssd1 vccd1 vccd1 _6093_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6686_ split18/X _6648_/X _6658_/X _6630_/A vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5637_ _6738_/A _6857_/A _7040_/A vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__o21a_1
XANTENNA__6523__A2 _6481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5568_ _6710_/A _5568_/B vssd1 vssd1 vccd1 vccd1 _5570_/C sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_7307_ _7378_/CLK _7307_/D vssd1 vssd1 vccd1 vccd1 _7307_/Q sky130_fd_sc_hd__dfxtp_1
X_4519_ _7375_/Q _7303_/Q _7295_/Q _7287_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4519_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold152 _6201_/X vssd1 vssd1 vccd1 vccd1 _6202_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6397__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 _6370_/X vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _7567_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _7337_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _5091_/X vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ _4049_/X hold213/X _7241_/S vssd1 vssd1 vccd1 vccd1 _7238_/X sky130_fd_sc_hd__mux2_1
X_5499_ _5499_/A _5499_/B vssd1 vssd1 vccd1 vccd1 _5500_/C sky130_fd_sc_hd__xor2_1
Xhold174 _7520_/Q vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _7434_/Q vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
X_7169_ _7169_/A _7169_/B _7169_/C vssd1 vssd1 vccd1 vccd1 _7233_/B sky130_fd_sc_hd__or3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7236__B1 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__B _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5014__A2 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4773__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4687__S1 _7453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _4083_/X _4869_/X _5022_/A vssd1 vssd1 vccd1 vccd1 _4870_/Y sky130_fd_sc_hd__a21oi_1
X_3821_ _7276_/Q _7591_/Q _7260_/Q _7484_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3821_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5894__B _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5386__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4764__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6071__A _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6540_ _6656_/A _6540_/B _6540_/C vssd1 vssd1 vccd1 vccd1 _6583_/C sky130_fd_sc_hd__and3_1
XFILLER_0_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3752_ _3759_/A _6216_/B vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__nor2_1
X_6471_ _6568_/A _6471_/B vssd1 vssd1 vccd1 vccd1 _6498_/B sky130_fd_sc_hd__xnor2_1
X_3683_ _3683_/A _6216_/C vssd1 vssd1 vccd1 vccd1 _3685_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5422_ _5788_/D _5415_/Y _5418_/Y _5417_/B vssd1 vssd1 vccd1 vccd1 _5422_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_0_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5353_ hold468/X _4679_/X _5355_/S vssd1 vssd1 vccd1 vccd1 _5353_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4304_ _4303_/X _4360_/B vssd1 vssd1 vccd1 vccd1 _4304_/Y sky130_fd_sc_hd__nand2b_1
X_5284_ hold492/X _5022_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _7427_/D sky130_fd_sc_hd__mux2_1
X_4235_ _4233_/X _4234_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__mux2_1
X_7023_ _7023_/A _7023_/B _7023_/C vssd1 vssd1 vccd1 vccd1 _7023_/X sky130_fd_sc_hd__and3_1
XANTENNA__7630__A _7630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4166_ _7347_/Q _4166_/B vssd1 vssd1 vccd1 vccd1 _4948_/B sky130_fd_sc_hd__or2_2
X_4097_ _6048_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__or2_1
XANTENNA__5788__C _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6807_ _6807_/A _6807_/B vssd1 vssd1 vccd1 vccd1 _6865_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5296__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4755__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4999_ _5026_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4999_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6738_ _6738_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6796_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6669_ _6771_/A _6669_/B vssd1 vssd1 vccd1 vccd1 _6747_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4669__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6983__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A1 _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5995__A _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4746__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout80 _4144_/Y vssd1 vssd1 vccd1 vccd1 _4162_/B sky130_fd_sc_hd__clkbuf_8
Xfanout91 _6162_/A vssd1 vssd1 vccd1 vccd1 _6356_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7145__C1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7449_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5171__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4357__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4020_ _6374_/A _4846_/A vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _5970_/A _5413_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5971_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4922_ _4955_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4853_ _6142_/S _4999_/B vssd1 vssd1 vccd1 vccd1 _4853_/Y sky130_fd_sc_hd__nand2_1
X_4784_ _4783_/X _4637_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7282_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4737__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3804_ _7363_/Q _3802_/X _3803_/Y _3798_/Y vssd1 vssd1 vccd1 vccd1 _6148_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5934__B1 _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7572_ _7577_/CLK _7572_/D vssd1 vssd1 vccd1 vccd1 _7572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6523_ _6507_/B _6481_/S _6522_/Y _6521_/X vssd1 vssd1 vccd1 vccd1 _6524_/B sky130_fd_sc_hd__a31o_1
X_3735_ _4021_/A _6417_/A vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6454_ _6637_/A _6454_/B vssd1 vssd1 vccd1 vccd1 _6468_/A sky130_fd_sc_hd__xnor2_2
X_5405_ hold435/X _4629_/X _5409_/S vssd1 vssd1 vccd1 vccd1 _5405_/X sky130_fd_sc_hd__mux2_1
X_3666_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5162__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4596__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6385_ input31/X _6384_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5336_ _4996_/X hold431/X _5338_/S vssd1 vssd1 vccd1 vccd1 _7450_/D sky130_fd_sc_hd__mux2_1
X_5267_ _7211_/C _5375_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5284_/S sky130_fd_sc_hd__and3_4
X_4218_ _4955_/B vssd1 vssd1 vccd1 vccd1 _4219_/B sky130_fd_sc_hd__inv_2
X_7006_ _7070_/A _7040_/A _6991_/X _7098_/A vssd1 vssd1 vccd1 vccd1 _7012_/C sky130_fd_sc_hd__a2bb2o_1
X_5198_ _4849_/X hold527/X _5212_/S vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4195__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4149_ _4964_/S _4728_/B vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4520__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6423__B _6427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3951__A2 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5153__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6102__B1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4833__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5392__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6892__A1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5695__A2 _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6170_ _6170_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6170_/X sky130_fd_sc_hd__or2_1
X_5121_ hold583/X _4937_/Y _5129_/S vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__mux2_1
X_5052_ hold310/X _4947_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _7320_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4309__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4003_ _7542_/Q input19/X hold52/A vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__a21o_2
XANTENNA__5412__B _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4743__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5954_ hold101/X wire79/X _5952_/Y _5953_/X _6218_/A vssd1 vssd1 vccd1 vccd1 _5954_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6524__A _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4905_ _6799_/A _4905_/B vssd1 vssd1 vccd1 vccd1 _4905_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6243__B _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5885_ _6273_/A _6771_/A _6840_/A _6630_/A vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__o2bb2a_1
X_4836_ hold195/X _4492_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7303_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7624_ _7624_/CLK hold59/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5383__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7555_ _7579_/CLK _7555_/D vssd1 vssd1 vccd1 vccd1 _7555_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767_ hold495/X _4719_/Y _4767_/S vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6506_ _6506_/A _6506_/B vssd1 vssd1 vccd1 vccd1 _6508_/A sky130_fd_sc_hd__or2_1
X_7486_ _7593_/CLK _7486_/D vssd1 vssd1 vccd1 vccd1 _7486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4698_ _4698_/A _4698_/B _4698_/C vssd1 vssd1 vccd1 vccd1 _4699_/B sky130_fd_sc_hd__or3_1
X_3718_ _6326_/B _6421_/B vssd1 vssd1 vccd1 vccd1 _3962_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3649_ hold64/X vssd1 vssd1 vccd1 vccd1 _3649_/Y sky130_fd_sc_hd__inv_2
X_6437_ _6437_/A _6437_/B vssd1 vssd1 vccd1 vccd1 _6437_/Y sky130_fd_sc_hd__nand2_1
X_6368_ hold60/X hold142/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6368_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5686__A2 _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5319_ hold186/X _5038_/X _5319_/S vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3792__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6635__A1 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7090__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6299_ _6297_/X _6298_/Y _7551_/Q _3716_/Y _6233_/Y vssd1 vssd1 vccd1 vccd1 _6314_/A
+ sky130_fd_sc_hd__a2111oi_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__buf_1
XANTENNA__6635__B2 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold180_A _7519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6399__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6434__A _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5610__A2 _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7115__A2 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5126__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7204__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7544_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5232__B _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3687__B _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7592_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _6808_/A _5788_/B _6771_/A _6773_/A vssd1 vssd1 vccd1 vccd1 _5701_/A sky130_fd_sc_hd__and4_1
XFILLER_0_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5365__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4621_ _4667_/B _4616_/X _4620_/X vssd1 vssd1 vccd1 vccd1 _6144_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__3907__S _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7340_ _7454_/CLK _7340_/D vssd1 vssd1 vccd1 vccd1 _7340_/Q sky130_fd_sc_hd__dfxtp_4
X_4552_ _4601_/B _4552_/B vssd1 vssd1 vccd1 vccd1 _4552_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7106__A2 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold504 _5148_/X vssd1 vssd1 vccd1 vccd1 _7366_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 _7388_/Q vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5117__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4483_ _4444_/Y _4482_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4483_/X sky130_fd_sc_hd__mux2_8
X_7271_ _7379_/CLK _7271_/D vssd1 vssd1 vccd1 vccd1 _7271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold515 _3995_/X vssd1 vssd1 vccd1 vccd1 _4002_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold548 _5157_/X vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 _7389_/Q vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _4077_/X vssd1 vssd1 vccd1 vccd1 _7454_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6222_ _3643_/Y _6220_/X _6221_/Y vssd1 vssd1 vccd1 vccd1 _6222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4738__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6153_/A _6153_/B vssd1 vssd1 vccd1 vccd1 _6153_/Y sky130_fd_sc_hd__nor2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5423__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6519__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5104_ _5103_/X _4921_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _7347_/D sky130_fd_sc_hd__mux2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6084_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6084_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6238__B _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5035_ _5034_/B _5032_/X _5033_/Y _5034_/Y _4963_/S vssd1 vssd1 vccd1 vccd1 _5035_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout183_A _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3878__A _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7042__A1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6986_ input33/X _4021_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _6986_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7042__B2 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4800__A0 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5937_ hold90/X wire79/X _5936_/X _6218_/A vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__o211a_1
XFILLER_0_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7607_ _7623_/CLK _7607_/D vssd1 vssd1 vccd1 vccd1 _7607_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _5869_/A _5869_/B _5869_/C vssd1 vssd1 vccd1 vccd1 _5904_/A sky130_fd_sc_hd__a21o_1
XANTENNA__4188__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4819_ hold246/X _4629_/X _4823_/S vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5799_ _5798_/A _5798_/Y _5800_/B _5747_/X vssd1 vssd1 vccd1 vccd1 _5800_/C sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7538_ _7538_/CLK _7538_/D vssd1 vssd1 vccd1 vccd1 _7538_/Q sky130_fd_sc_hd__dfxtp_1
X_7469_ _7489_/CLK _7469_/D vssd1 vssd1 vccd1 vccd1 _7469_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5108__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput57 _7558_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
Xoutput46 _7559_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
XANTENNA_fanout96_A _6022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput68 _7630_/X vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__buf_12
XFILLER_0_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6148__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4190__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3842__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5347__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7006__A1_N _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4705__S0 _7340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5389__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4181__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7024__A1 _7040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6840_ _6840_/A _6840_/B vssd1 vssd1 vccd1 vccd1 _7129_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__5586__A1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6771_ _6771_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6822_/B sky130_fd_sc_hd__xnor2_1
X_3983_ _3983_/A _4007_/A vssd1 vssd1 vccd1 vccd1 _4030_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5722_ _5843_/B _5720_/X _5688_/A _5689_/X vssd1 vssd1 vccd1 vccd1 _5723_/B sky130_fd_sc_hd__a211o_1
XANTENNA__6802__A _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5653_ _5736_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4322__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4604_ _4553_/B _4552_/B _4600_/Y vssd1 vssd1 vccd1 vccd1 _4604_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5418__A _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5584_ _5584_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5587_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5889__A2 _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 _7471_/Q vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
X_7323_ _7434_/CLK _7323_/D vssd1 vssd1 vccd1 vccd1 _7323_/Q sky130_fd_sc_hd__dfxtp_1
X_4535_ _6244_/A _4440_/A _4440_/Y _4534_/X vssd1 vssd1 vccd1 vccd1 _4535_/X sky130_fd_sc_hd__o22a_1
Xhold312 _7156_/X vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7395_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _7414_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6299__C1 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7254_ _7483_/CLK _7254_/D vssd1 vssd1 vccd1 vccd1 _7254_/Q sky130_fd_sc_hd__dfxtp_1
X_4466_ _7478_/Q _7466_/Q _7458_/Q _7252_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4466_/X sky130_fd_sc_hd__mux4_1
Xhold356 _7382_/Q vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _4737_/X vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _5063_/X vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _7219_/X vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
X_4397_ _4395_/X _4396_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4398_/B sky130_fd_sc_hd__mux2_1
Xhold389 _5115_/X vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_7185_ hold650/X _4580_/X _7191_/S vssd1 vssd1 vccd1 vccd1 _7185_/X sky130_fd_sc_hd__mux2_1
X_6205_ _5996_/A hold62/X _6207_/S vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6136_ _7604_/Q _6153_/A _6135_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6136_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4522__A_N _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6067_ _6922_/A _6065_/X _6066_/Y _4219_/B _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6067_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4077__A1 hold558/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4172__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5018_ _6093_/A _5018_/B vssd1 vssd1 vccd1 vccd1 _5019_/B sky130_fd_sc_hd__and2_1
XFILLER_0_68_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7015__A1 _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_as1802_215 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_215/HI io_out[26] sky130_fd_sc_hd__conb_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6969_ split4/X _6969_/B vssd1 vssd1 vccd1 vccd1 _6969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5329__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4232__A _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5510__B _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7006__B2 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4126__B _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4841__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3965__B _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3981__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4320_ _4320_/A _6053_/B vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__or2_1
XFILLER_0_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4251_ _7436_/Q _7428_/Q _7412_/Q _7404_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4251_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4182_ _4688_/S _4182_/B vssd1 vssd1 vccd1 vccd1 _4182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7245__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4059__A1 hold601/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5559__A1 _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6823_ _6823_/A _6823_/B vssd1 vssd1 vccd1 vccd1 _6824_/C sky130_fd_sc_hd__nand2_1
XANTENNA__4036__B _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout146_A _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6754_ _6754_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6831_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6532__A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3966_ _4267_/C _3970_/B _5974_/C _3965_/X vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6685_ _6685_/A _6685_/B vssd1 vssd1 vccd1 vccd1 _6685_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6251__B _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5705_ _5821_/A _6716_/A _6690_/A _5705_/D vssd1 vssd1 vccd1 vccd1 _5821_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3897_ _3895_/X _3896_/X _3931_/S vssd1 vssd1 vccd1 vccd1 _3897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5636_ _6690_/A _6637_/A vssd1 vssd1 vccd1 vccd1 _7040_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5567_ _5566_/B _5579_/S _6656_/A vssd1 vssd1 vccd1 vccd1 _5568_/B sky130_fd_sc_hd__o21a_1
X_4518_ _4516_/X _4517_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__mux2_1
X_7306_ _7306_/CLK _7306_/D vssd1 vssd1 vccd1 vccd1 _7306_/Q sky130_fd_sc_hd__dfxtp_1
X_5498_ _5498_/A vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__inv_2
Xhold142 _7565_/Q vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _6372_/X vssd1 vssd1 vccd1 vccd1 _6373_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _7543_/Q vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _7532_/Q vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _7443_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _5090_/X vssd1 vssd1 vccd1 vccd1 _7337_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _7374_/Q _7302_/Q _7294_/Q _7286_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4449_/X sky130_fd_sc_hd__mux4_1
X_7237_ _7236_/X hold58/X _7237_/S vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__mux2_1
Xhold175 _6174_/X vssd1 vssd1 vccd1 vccd1 _7520_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _5299_/X vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
X_7168_ _7168_/A _7168_/B _7168_/C _6416_/B vssd1 vssd1 vccd1 vccd1 _7169_/C sky130_fd_sc_hd__or4b_1
X_6119_ _6328_/A _4453_/Y _6118_/X _6375_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6119_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4926__S _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7070_/A _5958_/A _7096_/Y _3716_/Y _4037_/X vssd1 vssd1 vccd1 vccd1 _7102_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3769__C _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6426__B _6427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7172__B1 _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4568__A_N _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4897__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7227__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__A0 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3895__S0 _7360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4137__A _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5410__A0 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3820_ _7363_/Q _3818_/X _3819_/Y _3814_/Y vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3976__A _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3695__B _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3751_ _3759_/A _6216_/C vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6470_ _6568_/A _6471_/B _6453_/X vssd1 vssd1 vccd1 vccd1 _6485_/C sky130_fd_sc_hd__a21o_1
X_3682_ hold70/X vssd1 vssd1 vccd1 vccd1 _3682_/Y sky130_fd_sc_hd__inv_2
X_5421_ _5424_/B vssd1 vssd1 vccd1 vccd1 _5421_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5352_ _4589_/X hold573/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7461_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4600__A _4601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4303_ _4301_/X _4302_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4303_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5415__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5283_ hold491/X _5038_/X _5283_/S vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7022_ _7040_/B _7022_/B vssd1 vssd1 vccd1 vccd1 _7023_/C sky130_fd_sc_hd__nand2_1
X_4234_ _7426_/Q _7358_/Q _7350_/Q _7330_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4234_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4746__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7218__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4165_ _7344_/Q _7345_/Q _7346_/Q vssd1 vssd1 vccd1 vccd1 _4166_/B sky130_fd_sc_hd__or3_2
X_4096_ _4862_/A _6039_/A vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__or2_1
XANTENNA__5788__D _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4452__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ _6775_/Y _6802_/Y _6803_/X _5788_/D vssd1 vssd1 vccd1 vccd1 _6806_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3796__A1_N _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4998_ _5037_/B _4997_/Y _4964_/S vssd1 vssd1 vccd1 vccd1 _4998_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6737_ _6875_/A _6739_/B vssd1 vssd1 vccd1 vccd1 _6737_/X sky130_fd_sc_hd__and2_1
X_3949_ _4036_/A _6911_/B vssd1 vssd1 vccd1 vccd1 _3949_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6668_ _6771_/A _6669_/B vssd1 vssd1 vccd1 vccd1 _6668_/X sky130_fd_sc_hd__and2_1
X_6599_ _6710_/A _6652_/A vssd1 vssd1 vccd1 vccd1 _6600_/B sky130_fd_sc_hd__nand2_1
XANTENNA_hold106_A _7581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5619_ _5620_/B _5620_/C vssd1 vssd1 vccd1 vccd1 _6442_/B sky130_fd_sc_hd__or2_1
XANTENNA__6201__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7209__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout92 _6162_/A vssd1 vssd1 vccd1 vccd1 _6153_/A sky130_fd_sc_hd__buf_4
XFILLER_0_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout81 _4143_/X vssd1 vssd1 vccd1 vccd1 _4963_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__4404__B _4407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7145__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6900__A _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3958__A_N _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7207__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3801__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7581_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4357__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6066__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5885__A1_N _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3868__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4434__A1 _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ _5970_/A _5970_/B _5970_/C _5970_/D vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__or4_1
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4921_ _5022_/A _4921_/B vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__or2_4
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5397__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4852_ _6142_/S _4999_/B vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__or2_2
X_3803_ _3915_/A _3799_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _3803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4293__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4783_ hold475/X _4679_/X _4785_/S vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7571_ _7624_/CLK _7571_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6522_ _6522_/A _6522_/B vssd1 vssd1 vccd1 vccd1 _6522_/Y sky130_fd_sc_hd__nand2_1
X_3734_ _3988_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _6417_/A sky130_fd_sc_hd__nand2_1
X_3665_ _7363_/Q vssd1 vssd1 vccd1 vccd1 _3665_/Y sky130_fd_sc_hd__inv_2
X_6453_ _6637_/A _6454_/B vssd1 vssd1 vccd1 vccd1 _6453_/X sky130_fd_sc_hd__or2_1
X_5404_ _4538_/X _5403_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7488_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4596__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6384_ _6383_/A _6382_/X _6383_/Y _6311_/A vssd1 vssd1 vccd1 vccd1 _6384_/X sky130_fd_sc_hd__a22o_1
X_5335_ hold430/X _5015_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5335_/X sky130_fd_sc_hd__mux2_1
X_5266_ hold289/X _5022_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _7419_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _4689_/A _4215_/X _4216_/Y _4212_/Y vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7005_ _6265_/B _7009_/B _7004_/Y vssd1 vssd1 vccd1 vccd1 _7012_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__6257__A _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5197_ hold526/X _4864_/X _5211_/S vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__mux2_1
X_4148_ _7530_/Q _4145_/X _4162_/B vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__mux2_2
X_4079_ _4039_/C _4062_/Y _4078_/Y input16/X _7244_/A vssd1 vssd1 vccd1 vccd1 _4079_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4520__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4505__A _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4284__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7127__B1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold592_A hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_8_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6102__A1 _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4386__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7047__B1_N _7046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5916__A1 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6630__A _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5120_ _5119_/X _4897_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _7354_/D sky130_fd_sc_hd__mux2_1
X_5051_ hold309/X _4964_/X _5057_/S vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4104__B1 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ _4002_/A _4002_/B _4002_/C _4002_/D vssd1 vssd1 vccd1 vccd1 _4002_/X sky130_fd_sc_hd__or4_1
XFILLER_0_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5080__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5953_ _6628_/A _5811_/Y _5810_/X vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__a21o_1
X_4904_ _5001_/A _4900_/Y _4903_/X vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__o21a_1
X_5884_ _6273_/A _5918_/D _5859_/A _5861_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__a31o_1
X_4835_ hold194/X _4529_/X _4843_/S vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__mux2_1
X_7623_ _7623_/CLK _7623_/D vssd1 vssd1 vccd1 vccd1 _7623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4766_ _4765_/X _4637_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7274_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3918__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7554_ _7579_/CLK _7554_/D vssd1 vssd1 vccd1 vccd1 _7554_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6505_ _6529_/B _6505_/B _6505_/C _6505_/D vssd1 vssd1 vccd1 vccd1 _6505_/X sky130_fd_sc_hd__or4_4
X_3717_ _6326_/B _6421_/B vssd1 vssd1 vccd1 vccd1 _7123_/B sky130_fd_sc_hd__and2_1
X_7485_ _7485_/CLK _7485_/D vssd1 vssd1 vccd1 vccd1 _7485_/Q sky130_fd_sc_hd__dfxtp_1
X_4697_ _6096_/A _4701_/C _4696_/X vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4698__C _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6868__C1 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3648_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3648_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6436_ _6442_/A _6442_/B _5575_/X vssd1 vssd1 vccd1 vccd1 _6437_/B sky130_fd_sc_hd__o21a_1
X_6367_ _6373_/A _6367_/B vssd1 vssd1 vccd1 vccd1 _7564_/D sky130_fd_sc_hd__and2_1
X_5318_ hold233/X _4996_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _7442_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6298_ _6298_/A _6827_/A vssd1 vssd1 vccd1 vccd1 _6298_/Y sky130_fd_sc_hd__nand2_1
X_5249_ _7150_/B _7175_/B _5303_/C vssd1 vssd1 vccd1 vccd1 _5266_/S sky130_fd_sc_hd__and3_4
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7569_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5322__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__buf_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4934__S _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6399__B2 hold213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5071__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6450__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4582__A0 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6087__A0 _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5232__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4844__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6625__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7220__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4496__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4667_/B _4620_/B vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6562__A1 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4551_ _4601_/A _4879_/S vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_13_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold505 _7410_/Q vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _5197_/X vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
X_7270_ _7621_/CLK _7270_/D vssd1 vssd1 vccd1 vccd1 _7270_/Q sky130_fd_sc_hd__dfxtp_1
X_4482_ _4464_/X _4481_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__mux2_1
Xhold516 _4002_/X vssd1 vssd1 vccd1 vccd1 _7472_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold549 _7280_/Q vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _5199_/X vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6221_ _6922_/B _6220_/X _6015_/A vssd1 vssd1 vccd1 vccd1 _6221_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4420__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6152_ _6152_/A vssd1 vssd1 vccd1 vccd1 _6152_/Y sky130_fd_sc_hd__inv_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5704__A _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5103_ hold639/X _4937_/Y _5111_/S vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6078__A0 _4238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6519__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4628__A1 _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6328_/A _5002_/B _6082_/X _6375_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6083_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5142__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5034_ _6093_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _5034_/Y sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4754__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_A _7454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5053__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6985_ _6967_/X _6984_/Y _4723_/A vssd1 vssd1 vccd1 vccd1 _6985_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5936_ _6244_/A _5811_/Y _5934_/Y _5935_/Y _5810_/X vssd1 vssd1 vccd1 vccd1 _5936_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A _7544_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3894__A _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7606_ _7623_/CLK _7606_/D vssd1 vssd1 vccd1 vccd1 _7606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5867_ _5898_/B _5867_/B vssd1 vssd1 vccd1 vccd1 _5869_/C sky130_fd_sc_hd__or2_1
XFILLER_0_106_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4818_ _4817_/X _4538_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7296_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5798_ _5798_/A _7073_/A _5798_/C vssd1 vssd1 vccd1 vccd1 _5798_/Y sky130_fd_sc_hd__nand3_2
X_4749_ _7211_/B _7211_/C _5375_/C vssd1 vssd1 vccd1 vccd1 _4768_/S sky130_fd_sc_hd__and3_4
X_7537_ _7537_/CLK _7537_/D vssd1 vssd1 vccd1 vccd1 _7537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7468_ _7483_/CLK _7468_/D vssd1 vssd1 vccd1 vccd1 _7468_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6305__A1 _7040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6419_ _6419_/A _6419_/B _7168_/C _6417_/X vssd1 vssd1 vccd1 vccd1 _6427_/A sky130_fd_sc_hd__or4b_4
X_7399_ _7430_/CLK _7399_/D vssd1 vssd1 vccd1 vccd1 _7399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3833__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput58 _4006_/X vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput47 _7526_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
Xoutput69 _7631_/X vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__buf_12
XANTENNA__6069__A0 _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout89_A _4290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4108__A2_N _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5292__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6445__A _6445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5044__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4839__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7215__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4858__A1 _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5524__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4705__S1 _7341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5283__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5035__A1 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4469__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3982_ _6225_/A _5988_/A _3992_/C vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__or3_1
X_6770_ _6789_/A _6766_/Y _6767_/Y _6768_/X vssd1 vssd1 vccd1 vccd1 _6822_/A sky130_fd_sc_hd__a211o_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4794__A0 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5721_ _5688_/A _5689_/X _5843_/B _5720_/X vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__o211ai_2
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6802__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5652_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5739_/A sky130_fd_sc_hd__xnor2_1
X_4603_ _4553_/Y _4601_/C _4602_/X vssd1 vssd1 vccd1 vccd1 _4603_/Y sky130_fd_sc_hd__a21boi_1
X_5583_ _5533_/Y _5583_/B vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__and2b_1
Xhold302 _7488_/Q vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4641__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7322_ _7450_/CLK _7322_/D vssd1 vssd1 vccd1 vccd1 _7322_/Q sky130_fd_sc_hd__dfxtp_1
X_4534_ _4632_/C _4534_/B vssd1 vssd1 vccd1 vccd1 _4534_/X sky130_fd_sc_hd__and2_1
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold324 _5211_/X vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _5255_/X vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _7281_/Q vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6299__B1 _7551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 _7398_/Q vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _7278_/Q _7593_/Q _7262_/Q _7486_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4465_/X sky130_fd_sc_hd__mux4_1
Xhold357 _5183_/X vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _7369_/Q vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
X_7253_ _7481_/CLK _7253_/D vssd1 vssd1 vccd1 vccd1 _7253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold379 _7283_/Q vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
X_4396_ _7477_/Q _7465_/Q _7457_/Q _7251_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4396_/X sky130_fd_sc_hd__mux4_1
X_7184_ hold627/X _4492_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7184_/X sky130_fd_sc_hd__mux2_1
X_6204_ _6204_/A _6204_/B vssd1 vssd1 vccd1 vccd1 _7536_/D sky130_fd_sc_hd__or2_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6135_ _6153_/A _6135_/B vssd1 vssd1 vccd1 vccd1 _6135_/Y sky130_fd_sc_hd__nor2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6066_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6066_/Y sky130_fd_sc_hd__nor2_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4484__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5017_ hold424/X _4996_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _7314_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5274__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3889__A _6084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_as1802_216 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_216/HI io_out[27] sky130_fd_sc_hd__conb_1
XFILLER_0_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6968_ _6968_/A _6968_/B vssd1 vssd1 vccd1 vccd1 _6969_/B sky130_fd_sc_hd__xnor2_1
X_6899_ _7101_/A _3716_/Y _6287_/B vssd1 vssd1 vccd1 vccd1 _6899_/Y sky130_fd_sc_hd__a21oi_1
X_5919_ _6298_/A _6673_/A _5916_/Y _5941_/A vssd1 vssd1 vccd1 vccd1 _5920_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5265__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5017__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4407__B _4407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5973__C1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6114__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3965__C _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7190__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4250_ _4271_/A _5027_/A vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4181_ _7397_/Q _7389_/Q _7365_/Q _7381_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4182_/B sky130_fd_sc_hd__mux4_1
XANTENNA__5256__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6822_ _6822_/A _6822_/B vssd1 vssd1 vccd1 vccd1 _6831_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6753_ split7/X _6751_/Y _6752_/X vssd1 vssd1 vccd1 vccd1 _6771_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3965_ _6345_/A _5990_/A _6375_/A _3965_/D vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__and4_1
X_3896_ _7427_/Q _7359_/Q _7351_/Q _7331_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3896_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6684_ _6685_/A _6685_/B vssd1 vssd1 vccd1 vccd1 _6684_/X sky130_fd_sc_hd__and2_1
X_5704_ _6802_/A _6808_/A _6771_/A _6773_/A vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__and4_1
XFILLER_0_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _6683_/A _6742_/A vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5192__A0 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4614__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7181__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 _4052_/X vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5566_ _6710_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__and2_1
X_4517_ _7479_/Q _7467_/Q _7459_/Q _7253_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4517_/X sky130_fd_sc_hd__mux4_1
X_7305_ _7620_/CLK _7305_/D vssd1 vssd1 vccd1 vccd1 _7305_/Q sky130_fd_sc_hd__dfxtp_1
X_5497_ _5497_/A _5854_/C vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__and2_4
Xhold132 _7562_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _6368_/X vssd1 vssd1 vccd1 vccd1 _6369_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _6222_/Y vssd1 vssd1 vccd1 vccd1 _7543_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4689_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4448_/X sky130_fd_sc_hd__and2_1
Xhold176 _7331_/Q vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _7616_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _6195_/X vssd1 vssd1 vccd1 vccd1 _6196_/B sky130_fd_sc_hd__dlygate4sd3_1
X_7236_ _7234_/Y _7235_/X _7236_/B1 vssd1 vssd1 vccd1 vccd1 _7236_/X sky130_fd_sc_hd__o21a_1
Xhold187 _5319_/X vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _7339_/Q vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_7167_ _7166_/X _4685_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7598_/D sky130_fd_sc_hd__mux2_1
X_4379_ _6071_/B _6062_/B _4474_/A vssd1 vssd1 vccd1 vccd1 _5011_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5247__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6118_ _6025_/Y _6115_/Y _6117_/X vssd1 vssd1 vccd1 vccd1 _6118_/X sky130_fd_sc_hd__o21a_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7098_/A _7098_/B vssd1 vssd1 vccd1 vccd1 _7102_/B sky130_fd_sc_hd__nand2_1
X_6049_ _6417_/B _6047_/X _6048_/Y _4902_/B _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6049_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6995__A1 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3769__D _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5802__A _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6986__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3895__S1 _7361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3976__B _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _3759_/A _6216_/C vssd1 vssd1 vccd1 vccd1 _6191_/B sky130_fd_sc_hd__and2_2
XFILLER_0_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7163__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681_ _3681_/A vssd1 vssd1 vccd1 vccd1 _7547_/D sky130_fd_sc_hd__inv_2
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5420_ _6683_/B _5955_/B _5955_/D hold78/A vssd1 vssd1 vccd1 vccd1 _5424_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5351_ hold572/X _4629_/X _5355_/S vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__mux2_1
X_4302_ _7400_/Q _7392_/Q _7368_/Q _7384_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4302_/X sky130_fd_sc_hd__mux4_1
X_5282_ _5281_/X _4996_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _7426_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4233_ _7322_/Q _7338_/Q _7314_/Q _7450_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4233_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7021_ _7040_/B _7022_/B vssd1 vssd1 vccd1 vccd1 _7023_/B sky130_fd_sc_hd__or2_1
XANTENNA__3931__S _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6808__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5229__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4164_ _5376_/A _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _4720_/S sky130_fd_sc_hd__and3_4
XFILLER_0_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4095_ _5357_/A _5393_/A _5393_/B vssd1 vssd1 vccd1 vccd1 _4721_/S sky130_fd_sc_hd__or3_4
XFILLER_0_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4762__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5937__C1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6805_ _6790_/S _6802_/Y _6801_/Y _5788_/D vssd1 vssd1 vccd1 vccd1 _6811_/A sky130_fd_sc_hd__a211o_1
XANTENNA__5401__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4997_ _7350_/Q _4997_/B vssd1 vssd1 vccd1 vccd1 _4997_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6736_ _6690_/A _6690_/X split7/A vssd1 vssd1 vccd1 vccd1 _6739_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3948_ _3948_/A _7070_/A vssd1 vssd1 vccd1 vccd1 _3954_/A sky130_fd_sc_hd__nor2_1
XANTENNA__7154__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3879_ _6066_/A _6057_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _4971_/B sky130_fd_sc_hd__and3_1
X_6667_ _6611_/B _6666_/Y _6709_/S vssd1 vssd1 vccd1 vccd1 _6669_/B sky130_fd_sc_hd__mux2_2
X_6598_ _6597_/B _6603_/A _6603_/B _6596_/X _6555_/Y vssd1 vssd1 vccd1 vccd1 _6651_/A
+ sky130_fd_sc_hd__a311o_1
XANTENNA__6901__A1 _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5618_ _5615_/A _5615_/B _5617_/X _5616_/X _5612_/X vssd1 vssd1 vccd1 vccd1 _5622_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5549_ _5577_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5606__B _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3841__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7219_ hold366/X _4529_/X _7227_/S vssd1 vssd1 vccd1 vccd1 _7219_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6718__A _6718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4238__A _4238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5060__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6453__A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout82 _4116_/Y vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__buf_4
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7145__A1 _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7145__B2 _6166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6900__B _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout93 _4034_/Y vssd1 vssd1 vccd1 vccd1 _6162_/A sky130_fd_sc_hd__buf_4
XANTENNA__5156__A0 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4701__A _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3801__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7223__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6628__A _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7617_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output52_A _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3987__A _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4582__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3868__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _4940_/B _4106_/X _4915_/Y _4919_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _4921_/B
+ sky130_fd_sc_hd__o32a_1
X_4851_ _7176_/B _5322_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5039_/S sky130_fd_sc_hd__and3_4
X_3802_ _3800_/X _3801_/X _3931_/S vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4293__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4782_ hold314/X _4589_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7281_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7570_ _7570_/CLK _7570_/D vssd1 vssd1 vccd1 vccd1 _7570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7194__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6521_ _6521_/A _6521_/B _6521_/C _6521_/D vssd1 vssd1 vccd1 vccd1 _6521_/X sky130_fd_sc_hd__and4_1
X_3733_ _3733_/A _3733_/B _3983_/A vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__or3_1
X_3664_ _3915_/A vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__inv_2
X_6452_ _5595_/X _6451_/Y _6463_/S vssd1 vssd1 vccd1 vccd1 _6454_/B sky130_fd_sc_hd__mux2_1
X_5403_ hold302/X _4580_/X _5409_/S vssd1 vssd1 vccd1 vccd1 _5403_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5426__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6383_ _6383_/A _6383_/B vssd1 vssd1 vccd1 vccd1 _6383_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_100_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5334_ _4973_/X _5333_/X _5338_/S vssd1 vssd1 vccd1 vccd1 _5334_/X sky130_fd_sc_hd__mux2_1
X_5265_ hold288/X _5038_/X _5265_/S vssd1 vssd1 vccd1 vccd1 _5265_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4757__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5196_ _5376_/A _7194_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5211_/S sky130_fd_sc_hd__and3_4
X_4216_ _4401_/S _4210_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4216_/Y sky130_fd_sc_hd__a21oi_1
X_7004_ _6265_/B _7009_/B _7020_/A vssd1 vssd1 vccd1 vccd1 _7004_/Y sky130_fd_sc_hd__o21ai_1
X_4147_ _6220_/C _4290_/D _6023_/S vssd1 vssd1 vccd1 vccd1 _4147_/X sky130_fd_sc_hd__or3_2
XANTENNA__6257__B _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ _6869_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _4078_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6273__A _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4284__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6719_ _6719_/A _6719_/B vssd1 vssd1 vccd1 vccd1 _6719_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7043__S _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7063__B1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4118__D _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6911__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5916__A2 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6630__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7218__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4431__A _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6122__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4352__A1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5050_ _5049_/X _4921_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _7319_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4104__A1 _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _3965_/D _6375_/A _5990_/A _4001_/D vssd1 vssd1 vccd1 vccd1 _4002_/D sky130_fd_sc_hd__and4b_1
XFILLER_0_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6093__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _5952_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5952_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6801__B1 _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5201__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4903_ _4209_/A _4698_/A _4902_/Y _4901_/X _4263_/B vssd1 vssd1 vccd1 vccd1 _4903_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5368__A0 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5883_ hold508/X wire79/X _5881_/Y _5882_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _5883_/X
+ sky130_fd_sc_hd__o221a_1
X_4834_ hold273/X _4443_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7302_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7622_ _7623_/CLK _7622_/D vssd1 vssd1 vccd1 vccd1 _7622_/Q sky130_fd_sc_hd__dfxtp_1
X_4765_ hold363/X _4679_/X _4767_/S vssd1 vssd1 vccd1 vccd1 _4765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3918__A1 _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7553_ _7579_/CLK _7553_/D vssd1 vssd1 vccd1 vccd1 _7553_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6032__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6504_ _6505_/C _6505_/D vssd1 vssd1 vccd1 vccd1 _6504_/Y sky130_fd_sc_hd__nor2_1
X_3716_ _4036_/A _3716_/B vssd1 vssd1 vccd1 vccd1 _3716_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_fanout121_A _7590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7484_ _7592_/CLK _7484_/D vssd1 vssd1 vccd1 vccd1 _7484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4696_ _6142_/S _4694_/A _4930_/S vssd1 vssd1 vccd1 vccd1 _4696_/X sky130_fd_sc_hd__a21o_1
X_3647_ hold80/X vssd1 vssd1 vccd1 vccd1 _3647_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6435_ _6435_/A vssd1 vssd1 vccd1 vccd1 _6435_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6366_ _7527_/Q hold126/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6366_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5317_ hold232/X _5015_/X _5319_/S vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__mux2_1
X_6297_ _7109_/B _7108_/B _6238_/X vssd1 vssd1 vccd1 vccd1 _6297_/X sky130_fd_sc_hd__a21o_1
X_5248_ _5022_/X hold536/X _5248_/S vssd1 vssd1 vccd1 vccd1 _7411_/D sky130_fd_sc_hd__mux2_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ hold531/X _4864_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__mux2_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6207__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold500_A _7523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4885__A2 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4193__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4496__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4161__A _4751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4550_ _4601_/B vssd1 vssd1 vccd1 vccd1 _4553_/B sky130_fd_sc_hd__inv_2
Xhold517 _7399_/Q vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 _5245_/X vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ _6120_/A _4986_/S _4525_/B _4480_/Y vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold528 _5198_/X vssd1 vssd1 vccd1 vccd1 _7388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _7405_/Q vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _6417_/A _6220_/B _6220_/C _6220_/D vssd1 vssd1 vccd1 vccd1 _6220_/X sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7479_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4420__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6151_ _4698_/C _6153_/B _6160_/S vssd1 vssd1 vccd1 vccd1 _6152_/A sky130_fd_sc_hd__mux2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5704__B _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5102_ _5101_/X _4897_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _7346_/D sky130_fd_sc_hd__mux2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6082_ _6025_/Y _6079_/Y _6081_/X vssd1 vssd1 vccd1 vccd1 _6082_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4628__A2 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4184__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5033_ _5032_/C _5032_/B _4376_/Y vssd1 vssd1 vccd1 vccd1 _5033_/Y sky130_fd_sc_hd__a21boi_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7027__B1 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6984_ _4030_/B _6982_/X _6983_/X vssd1 vssd1 vccd1 vccd1 _6984_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout169_A _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5935_ _5970_/A _5457_/S _5952_/A vssd1 vssd1 vccd1 vccd1 _5935_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5866_ _5866_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__nor2_1
X_4817_ hold211/X _4580_/X _4823_/S vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7605_ _7621_/CLK _7605_/D vssd1 vssd1 vccd1 vccd1 _7605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5797_ _5797_/A _5797_/B _5797_/C vssd1 vssd1 vccd1 vccd1 _5798_/C sky130_fd_sc_hd__nand3_1
X_4748_ _4748_/A _4825_/B vssd1 vssd1 vccd1 vccd1 _5375_/C sky130_fd_sc_hd__nor2_4
X_7536_ _7536_/CLK _7536_/D vssd1 vssd1 vccd1 vccd1 _7536_/Q sky130_fd_sc_hd__dfxtp_1
X_7467_ _7481_/CLK _7467_/D vssd1 vssd1 vccd1 vccd1 _7467_/Q sky130_fd_sc_hd__dfxtp_1
X_4679_ _4529_/S _4663_/X _4678_/X _4640_/Y vssd1 vssd1 vccd1 vccd1 _4679_/X sky130_fd_sc_hd__a31o_4
XANTENNA__5513__B1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6418_ _6417_/B _3988_/A _4139_/B vssd1 vssd1 vccd1 vccd1 _7168_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7398_ _7400_/CLK _7398_/D vssd1 vssd1 vccd1 vccd1 _7398_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput48 _5660_/B vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
Xoutput59 _7543_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6349_ _6349_/A _6419_/A vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4175__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__A _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5029__C1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4680__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5805__A _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5807__A1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3913__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4469__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _6223_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _3988_/C sky130_fd_sc_hd__or2_1
XFILLER_0_85_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5720_ _5843_/A _5718_/X _5658_/X _5662_/A vssd1 vssd1 vccd1 vccd1 _5720_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5991__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5651_ _5651_/A _5651_/B vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__nor2_1
X_4602_ _4999_/B _4698_/B vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5582_ _6442_/A _6437_/A vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__or2_1
XANTENNA__4641__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7321_ _7451_/CLK _7321_/D vssd1 vssd1 vccd1 vccd1 _7321_/Q sky130_fd_sc_hd__dfxtp_1
X_4533_ _6139_/A _4533_/B vssd1 vssd1 vccd1 vccd1 _4534_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold303 _7435_/Q vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _7592_/CLK _7252_/D vssd1 vssd1 vccd1 vccd1 _7252_/Q sky130_fd_sc_hd__dfxtp_1
Xhold314 _4781_/X vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _7376_/Q vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _5219_/X vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _5256_/X vssd1 vssd1 vccd1 vccd1 _7414_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _5184_/X vssd1 vssd1 vccd1 vccd1 _7382_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _5154_/X vssd1 vssd1 vccd1 vccd1 _7369_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ input2/X _5031_/S _4462_/X _4463_/X vssd1 vssd1 vccd1 vccd1 _4464_/X sky130_fd_sc_hd__o22a_1
X_6203_ _5999_/A hold68/X _6207_/S vssd1 vssd1 vccd1 vccd1 _6203_/X sky130_fd_sc_hd__mux2_1
X_4395_ _7277_/Q _7592_/Q _7261_/Q _7485_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4395_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7183_ hold626/X _4529_/X _7191_/S vssd1 vssd1 vccd1 vccd1 _7183_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6134_ _6134_/A vssd1 vssd1 vccd1 vccd1 _6134_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4765__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6065_ _6328_/A _4219_/B _6064_/X _6375_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6065_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5016_ hold423/X _5015_/X _5039_/S vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3904__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6980__S _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_as1802_217 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_217/HI io_out[28] sky130_fd_sc_hd__conb_1
X_6967_ _6961_/X _6964_/Y _6966_/X _6220_/C vssd1 vssd1 vccd1 vccd1 _6967_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4785__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5918_ _5916_/Y _5941_/A _6516_/A _5918_/D vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__and4bb_1
XFILLER_0_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6898_ _4084_/A _6909_/B _6897_/S _5879_/A vssd1 vssd1 vccd1 vccd1 _6898_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_91_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5849_ _6808_/A _5811_/Y _5848_/X _5811_/A _5810_/X vssd1 vssd1 vccd1 vccd1 _5849_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4537__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7519_ _7534_/CLK _7519_/D vssd1 vssd1 vccd1 vccd1 _7519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4396__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4776__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7226__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4180_ _4271_/A vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6821_ _6841_/A _6817_/B _6817_/C _6838_/B _6819_/X vssd1 vssd1 vccd1 vccd1 _6821_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4216__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5413__C1 _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4767__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6752_ _6756_/A _6675_/X _6751_/B _6711_/Y _6673_/B vssd1 vssd1 vccd1 vccd1 _6752_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3964_ _4113_/B _6375_/C vssd1 vssd1 vccd1 vccd1 _6331_/A sky130_fd_sc_hd__or2_1
X_3895_ _7323_/Q _7339_/Q _7315_/Q _7451_/Q _7360_/Q _7361_/Q vssd1 vssd1 vccd1 vccd1
+ _3895_/X sky130_fd_sc_hd__mux4_1
X_6683_ _6683_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _6685_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5703_ _5705_/D vssd1 vssd1 vccd1 vccd1 _5703_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5634_ _5634_/A _5634_/B _5634_/C vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__or3_1
XANTENNA__4614__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7304_ _7487_/CLK _7304_/D vssd1 vssd1 vccd1 vccd1 _7304_/Q sky130_fd_sc_hd__dfxtp_1
Xhold100 _7246_/X vssd1 vssd1 vccd1 vccd1 _7568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ _6532_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _6431_/A sky130_fd_sc_hd__xnor2_2
X_4516_ _7279_/Q _7594_/Q _7263_/Q _7487_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4516_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout201_A _7341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 _4053_/X vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _5854_/C _5497_/A vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__or2_4
Xhold122 _7536_/Q vssd1 vssd1 vccd1 vccd1 _5999_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _6362_/X vssd1 vssd1 vccd1 vccd1 _6363_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold144 _7525_/Q vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4445_/X _4446_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4448_/B sky130_fd_sc_hd__mux2_1
Xhold177 _5075_/X vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _7213_/X vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _7534_/Q vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7235_ _6328_/A _7230_/C _6220_/C _5980_/B vssd1 vssd1 vccd1 vccd1 _7235_/X sky130_fd_sc_hd__a31o_1
X_7166_ hold201/X _4719_/Y _7166_/S vssd1 vssd1 vccd1 vccd1 _7166_/X sky130_fd_sc_hd__mux2_1
Xhold199 _5093_/X vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _7614_/Q vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _7602_/Q _6153_/A _6116_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6117_/X sky130_fd_sc_hd__a211o_1
X_4378_ _5011_/A _5012_/A _4376_/Y _4377_/X vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__o31ai_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _6235_/A _7025_/A _7551_/Q vssd1 vssd1 vccd1 vccd1 _7098_/B sky130_fd_sc_hd__mux2_1
X_6048_ _6048_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6048_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4508__B _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4302__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4758__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5183__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4247__A1_N _7455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4369__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6986__A2 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3992__B _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3680_ _3680_/A vssd1 vssd1 vccd1 vccd1 _7546_/D sky130_fd_sc_hd__inv_2
XANTENNA__5174__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5350_ _4538_/X _5349_/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7460_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4301_ _7440_/Q _7432_/Q _7416_/Q _7408_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4301_/X sky130_fd_sc_hd__mux4_1
X_5281_ hold446/X _5015_/X _5283_/S vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4232_ _4688_/S _4232_/B vssd1 vssd1 vccd1 vccd1 _4232_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7020_ _7020_/A _7020_/B _7020_/C vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__and3_1
XANTENNA__6808__B _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5204__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6096__A _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4163_ _4163_/A _4163_/B _4658_/A _4850_/B vssd1 vssd1 vccd1 vccd1 _7212_/B sky130_fd_sc_hd__or4b_4
X_4094_ _6198_/A _4440_/A _4846_/C vssd1 vssd1 vccd1 vccd1 _7211_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4996_ _3939_/X _4083_/X _5022_/A _4995_/X vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__a211o_4
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6804_ _6832_/A _6802_/Y _6801_/Y vssd1 vssd1 vccd1 vccd1 _6807_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6735_ _6869_/A _6735_/B vssd1 vssd1 vccd1 vccd1 _6786_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3947_ _4036_/A _3962_/B vssd1 vssd1 vccd1 vccd1 _7070_/A sky130_fd_sc_hd__or2_4
XFILLER_0_46_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3878_ _6057_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _4940_/B sky130_fd_sc_hd__and2_1
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6666_ _6666_/A _6666_/B vssd1 vssd1 vccd1 vccd1 _6666_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5165__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5617_ _5603_/X _5607_/B _5614_/B _5605_/X _5589_/X vssd1 vssd1 vccd1 vccd1 _5617_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6362__A0 _7570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6597_ _6597_/A _6597_/B vssd1 vssd1 vccd1 vccd1 _6643_/B sky130_fd_sc_hd__and2_1
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4912__A1 _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5548_ _5545_/X _5572_/B _5525_/Y _5529_/Y vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__a211o_4
XANTENNA__6114__A0 _4460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7218_ hold291/X _4443_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7618_/D sky130_fd_sc_hd__mux2_1
X_5479_ _6568_/A _5479_/B vssd1 vssd1 vccd1 vccd1 _5479_/Y sky130_fd_sc_hd__nand2_1
X_7149_ _6235_/A _6926_/Y _7147_/X _7148_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7590_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4979__A1 _6882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout83 _4685_/A vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7145__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout94 _3975_/X vssd1 vssd1 vccd1 vccd1 _6922_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6105__A0 _4407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6909__A _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6408__A1 _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output45_A _7540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4850_ _4850_/A _4850_/B vssd1 vssd1 vccd1 vccd1 _5322_/C sky130_fd_sc_hd__nand2_8
XANTENNA__5395__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3801_ _7273_/Q _7613_/Q _7605_/Q _7621_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3801_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4781_ hold313/X _4629_/X _4785_/S vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6520_ _6518_/A _6518_/B _6576_/A vssd1 vssd1 vccd1 vccd1 _6569_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3732_ _6383_/A _4122_/C _3988_/B vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__and3_1
XANTENNA__5147__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3663_ _3663_/A vssd1 vssd1 vccd1 vccd1 _3663_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6451_ _6451_/A _6451_/B vssd1 vssd1 vccd1 vccd1 _6451_/Y sky130_fd_sc_hd__xnor2_1
X_5402_ _4492_/X hold408/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7487_/D sky130_fd_sc_hd__mux2_1
X_6382_ hold136/X _6415_/A _6356_/B hold66/X vssd1 vssd1 vccd1 vccd1 _6382_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5333_ hold417/X _4990_/Y _5337_/S vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5264_ _5263_/X _4996_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _7418_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5195_ _5357_/A _5321_/B _7193_/C vssd1 vssd1 vccd1 vccd1 _5212_/S sky130_fd_sc_hd__or3b_4
X_4215_ _4213_/X _4214_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4215_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7003_ _6989_/A _5793_/X _7002_/Y split7/X _5970_/A vssd1 vssd1 vccd1 vccd1 _7003_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout199_A _7341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ _6329_/A _4279_/C _6162_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__and3_4
XANTENNA__4773__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4077_ _4076_/X hold558/X _7249_/S vssd1 vssd1 vccd1 vccd1 _4077_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6554__A _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6273__B _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5386__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4979_ _6882_/A _4905_/B _4978_/X vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6718_ _6718_/A _6718_/B vssd1 vssd1 vccd1 vccd1 _6766_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6649_ _6617_/A _6616_/X _6708_/A _6648_/A vssd1 vssd1 vccd1 vccd1 _6658_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6099__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__A _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5310__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6464__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5129__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6639__A _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5301__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4159__A _7527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ _3970_/B _3999_/X _3997_/X _7244_/A vssd1 vssd1 vccd1 vccd1 _4002_/C sky130_fd_sc_hd__a211o_1
XANTENNA__6374__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6093__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5951_ _5955_/A _5434_/S _5964_/B _5950_/Y vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4902_ _4902_/A _4902_/B vssd1 vssd1 vccd1 vccd1 _4902_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _6802_/A _5811_/Y _5810_/X vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__a21o_1
X_4833_ hold272/X _4483_/X _4843_/S vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__mux2_1
X_7621_ _7621_/CLK _7621_/D vssd1 vssd1 vccd1 vccd1 _7621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4764_ hold349/X _4589_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7273_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4622__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7552_ _7599_/CLK _7552_/D vssd1 vssd1 vccd1 vccd1 _7552_/Q sky130_fd_sc_hd__dfxtp_1
X_7483_ _7483_/CLK _7483_/D vssd1 vssd1 vccd1 vccd1 _7483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6503_ _6611_/A _6503_/B _6503_/C vssd1 vssd1 vccd1 vccd1 _6505_/D sky130_fd_sc_hd__and3_1
X_3715_ _4036_/A _6326_/B hold97/A vssd1 vssd1 vccd1 vccd1 _7020_/A sky130_fd_sc_hd__and3_4
XFILLER_0_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4695_ _4695_/A _4699_/A vssd1 vssd1 vccd1 vccd1 _4701_/C sky130_fd_sc_hd__xnor2_1
X_6434_ _6840_/A _6434_/B vssd1 vssd1 vccd1 vccd1 _6435_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout114_A _3665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _3646_/A vssd1 vssd1 vccd1 vccd1 _3646_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4768__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6365_ _6373_/A _6365_/B vssd1 vssd1 vccd1 vccd1 _7563_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5316_ _5315_/X _4973_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _5316_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6296_ _6240_/X _7051_/B _6242_/X vssd1 vssd1 vccd1 vccd1 _7108_/B sky130_fd_sc_hd__o21a_1
X_5247_ hold535/X _5038_/X _5247_/S vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__mux2_1
X_5178_ _5376_/A _7212_/A _5322_/C vssd1 vssd1 vccd1 vccd1 _5193_/S sky130_fd_sc_hd__and3_4
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7045__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
X_4129_ _5974_/C _4128_/X _4127_/X vssd1 vssd1 vccd1 vccd1 _4163_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3701__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5359__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4532__A _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4193__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6194__A _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7036__A1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7036__B2 _6338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5302__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6922__A _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6133__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__B _4827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold507 _5246_/X vssd1 vssd1 vccd1 vccd1 _7410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _7265_/Q vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4480_ _4479_/A _4479_/B _5034_/B vssd1 vssd1 vccd1 vccd1 _4480_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold529 _7440_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6150_ _6149_/X hold68/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__mux2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5101_ hold633/X _4912_/Y _5111_/S vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__mux2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6081_ _7350_/Q _6153_/A _6080_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4708__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4184__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5032_ _4376_/Y _5032_/B _5032_/C vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__and3b_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5212__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6983_ _6048_/A _5804_/C _4029_/Y _6120_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _6983_/X
+ sky130_fd_sc_hd__a221o_1
X_5934_ _5932_/X _5933_/Y _5955_/A vssd1 vssd1 vccd1 vccd1 _5934_/Y sky130_fd_sc_hd__o21ai_1
X_5865_ _5866_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__and2_1
X_4816_ hold183/X _4492_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7295_/D sky130_fd_sc_hd__mux2_1
X_7604_ _7608_/CLK _7604_/D vssd1 vssd1 vccd1 vccd1 _7604_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5210__A0 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5796_ _7069_/B _7069_/C _7069_/A vssd1 vssd1 vccd1 vccd1 _7073_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747_ _4747_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _7211_/C sky130_fd_sc_hd__nor2_2
X_7535_ _7538_/CLK _7535_/D vssd1 vssd1 vccd1 vccd1 _7535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7466_ _7592_/CLK _7466_/D vssd1 vssd1 vccd1 vccd1 _7466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4678_ _4986_/S _4676_/Y _4677_/Y _4144_/Y vssd1 vssd1 vccd1 vccd1 _4678_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7397_ _4004_/A _7397_/D vssd1 vssd1 vccd1 vccd1 _7397_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4498__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6417_ _6417_/A _6417_/B _4009_/A vssd1 vssd1 vccd1 vccd1 _6417_/X sky130_fd_sc_hd__or3b_1
Xoutput49 _5788_/D vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6348_ _6374_/A _5977_/B _6225_/A _5988_/A _4021_/A vssd1 vssd1 vccd1 vccd1 _6419_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6279_ _7035_/B _6279_/B vssd1 vssd1 vccd1 vccd1 _7009_/B sky130_fd_sc_hd__nor2_4
XANTENNA__4175__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7018__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__B _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5122__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6226__C1 _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6742__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold610_A _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5077__B _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4437__A _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3913__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4491__A1 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3980_ _3980_/A _6328_/B _3980_/C vssd1 vssd1 vccd1 vccd1 _3980_/X sky130_fd_sc_hd__and3_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5991__A1 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _6273_/A _5788_/D _5630_/X _5634_/A vssd1 vssd1 vccd1 vccd1 _5651_/B sky130_fd_sc_hd__a211oi_1
XFILLER_0_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4601_ _4601_/A _4601_/B _4601_/C vssd1 vssd1 vccd1 vccd1 _4698_/B sky130_fd_sc_hd__or3_2
XFILLER_0_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _6442_/A _6437_/A vssd1 vssd1 vccd1 vccd1 _5621_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_108_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7320_ _7424_/CLK _7320_/D vssd1 vssd1 vccd1 vccd1 _7320_/Q sky130_fd_sc_hd__dfxtp_1
X_4532_ _6139_/A _4533_/B vssd1 vssd1 vccd1 vccd1 _4632_/C sky130_fd_sc_hd__or2_1
XFILLER_0_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold304 _5301_/X vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ _7485_/CLK _7251_/D vssd1 vssd1 vccd1 vccd1 _7251_/Q sky130_fd_sc_hd__dfxtp_1
Xhold326 _7386_/Q vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _4118_/B _4455_/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4463_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold315 _6827_/A vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__5207__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold337 _7439_/Q vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 _7332_/Q vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _7273_/Q vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6218_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _7535_/D sky130_fd_sc_hd__nand2_1
X_7182_ _7181_/X _4443_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7602_/D sky130_fd_sc_hd__mux2_1
X_4394_ _5022_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__or2_4
XANTENNA__7248__A1 hold558/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6133_ _4601_/B _6135_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6827__A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6025_/Y _6061_/Y _6063_/X vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__o21a_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _4964_/S _5010_/X _5014_/X _4998_/Y vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__a31o_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3904__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4781__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6966_ _3716_/Y _6959_/Y _6965_/X _6913_/A vssd1 vssd1 vccd1 vccd1 _6966_/X sky130_fd_sc_hd__o22a_1
Xwrapped_as1802_218 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_218/HI io_out[29] sky130_fd_sc_hd__conb_1
XFILLER_0_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5917_ _6273_/A _6827_/A _6341_/A vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__and3_1
XANTENNA__4082__A _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6897_ _6311_/A _6909_/B _6897_/S vssd1 vssd1 vccd1 vccd1 _6897_/X sky130_fd_sc_hd__mux2_4
XANTENNA__5982__A1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _5879_/A _5579_/S _5877_/B _5847_/Y vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_51_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5779_ _5775_/A _5775_/B _5775_/C vssd1 vssd1 vccd1 vccd1 _5780_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7518_ _7537_/CLK hold89/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3745__B1 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3840__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7449_ _7449_/CLK _7449_/D vssd1 vssd1 vccd1 vccd1 _7449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5117__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4396__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_A _3975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4956__S _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7239__A1 hold60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6737__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold658_A _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5816__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3831__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5535__B _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6686__C1 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4866__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6647__A _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output75_A _7524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4464__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4216__A1 _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6820_ _6844_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6838_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5413__B1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6751_ _6751_/A _6751_/B vssd1 vssd1 vccd1 vccd1 _6751_/Y sky130_fd_sc_hd__xnor2_1
X_3963_ _6326_/C _4140_/B vssd1 vssd1 vccd1 vccd1 _6375_/C sky130_fd_sc_hd__and2_2
X_3894_ _7363_/Q _3894_/B vssd1 vssd1 vccd1 vccd1 _3894_/X sky130_fd_sc_hd__and2_1
XFILLER_0_73_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6682_ split18/X _6648_/X _6658_/X _6683_/A vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__a211o_1
X_5702_ _6802_/A _6771_/A _6773_/A _6808_/A vssd1 vssd1 vccd1 vccd1 _5705_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_5_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5633_ _6311_/A _6716_/A vssd1 vssd1 vccd1 vccd1 _5634_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _5556_/B _5563_/Y _5579_/S vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__mux2_2
XANTENNA__3822__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7303_ _7378_/CLK _7303_/D vssd1 vssd1 vccd1 vccd1 _7303_/Q sky130_fd_sc_hd__dfxtp_1
X_4515_ input3/X _4514_/Y _5031_/S vssd1 vssd1 vccd1 vccd1 _4515_/X sky130_fd_sc_hd__mux2_1
Xhold101 _7497_/Q vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold112 _7239_/X vssd1 vssd1 vccd1 vccd1 _7528_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ _5464_/B _5494_/Y _5495_/S vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__mux2_4
Xhold123 _6203_/X vssd1 vssd1 vccd1 vccd1 _6204_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 _7500_/Q vssd1 vssd1 vccd1 vccd1 _6216_/C sky130_fd_sc_hd__buf_2
X_4446_ _7478_/Q _7466_/Q _7458_/Q _7252_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4446_/X sky130_fd_sc_hd__mux4_1
Xhold156 _6199_/X vssd1 vssd1 vccd1 vccd1 _6200_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _6189_/X vssd1 vssd1 vccd1 vccd1 _7525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _7526_/Q vssd1 vssd1 vccd1 vccd1 _6191_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7234_ _7555_/Q _3698_/A _7230_/B vssd1 vssd1 vccd1 vccd1 _7234_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4776__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7165_ _7164_/X _4637_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7597_/D sky130_fd_sc_hd__mux2_1
Xhold189 _7469_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _7621_/Q vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _6071_/B _6062_/B _6080_/B _6089_/B _4320_/A vssd1 vssd1 vccd1 vccd1 _4377_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__7152__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6116_ _6153_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/A _7109_/B vssd1 vssd1 vccd1 vccd1 _7096_/Y sky130_fd_sc_hd__xnor2_1
X_6047_ _6328_/A _4902_/B _6046_/X _6375_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6047_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4455__B2 _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6991__S _7551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5404__A0 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5400__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4302__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6949_ _6949_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6949_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5636__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3813__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6380__A1 _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4369__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__B1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6467__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4906__C1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5546__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6141__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4382__B1 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5280_ _5279_/X _4973_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__mux2_1
X_4300_ _4474_/A _6071_/B vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__xnor2_1
X_4231_ _7402_/Q _7394_/Q _7370_/Q _7386_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4232_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5882__B1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _4846_/A _4162_/B _4964_/S vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__and3_2
X_4093_ _6198_/A _4440_/A _4846_/C vssd1 vssd1 vccd1 vccd1 _5393_/B sky130_fd_sc_hd__and3_2
XFILLER_0_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5220__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4344__B _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4296__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4995_ _4918_/Y _4993_/Y _4994_/X vssd1 vssd1 vccd1 vccd1 _4995_/X sky130_fd_sc_hd__o21a_1
X_6803_ _6803_/A1 _6774_/Y _6738_/A _6765_/X vssd1 vssd1 vccd1 vccd1 _6803_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout144_A _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6734_ _6734_/A _6734_/B vssd1 vssd1 vccd1 vccd1 _6781_/B sky130_fd_sc_hd__and2_1
XANTENNA__6840__A _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ _4037_/A _3962_/B vssd1 vssd1 vccd1 vccd1 _3946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6051__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3877_ _6048_/A _4862_/A _6039_/A vssd1 vssd1 vccd1 vccd1 _4915_/B sky130_fd_sc_hd__and3_1
X_6665_ _6670_/A _6670_/B _6640_/A vssd1 vssd1 vccd1 vccd1 _6666_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6898__C1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6596_ _6597_/B _6596_/B vssd1 vssd1 vccd1 vccd1 _6596_/X sky130_fd_sc_hd__and2_1
X_5616_ _5598_/B _5598_/C _6799_/A _5616_/C1 vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5547_ _5547_/A1 _5572_/B _5529_/Y vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5478_ _5454_/A _5454_/B _5452_/Y _5479_/B vssd1 vssd1 vccd1 vccd1 _5486_/C sky130_fd_sc_hd__a31o_1
X_7217_ hold290/X _4483_/X _7227_/S vssd1 vssd1 vccd1 vccd1 _7217_/X sky130_fd_sc_hd__mux2_1
X_4429_ _4428_/A _4428_/B _4986_/S vssd1 vssd1 vccd1 vccd1 _4429_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4220__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6287__A _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3704__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7148_ input38/X _4723_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _7148_/X sky130_fd_sc_hd__a21o_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ _7064_/X _7078_/X _7078_/A _6339_/A vssd1 vssd1 vccd1 vccd1 _7079_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5130__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6050__A0 _6049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout84 _4147_/X vssd1 vssd1 vccd1 vccd1 _4964_/S sky130_fd_sc_hd__buf_6
XFILLER_0_52_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout95 _3702_/Y vssd1 vssd1 vccd1 vccd1 _6328_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6353__A1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4903__A2 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4211__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5616__B1 _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5040__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4780_ _4779_/X _4538_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7280_/D sky130_fd_sc_hd__mux2_1
X_3800_ _7377_/Q _7305_/Q _7297_/Q _7289_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3800_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3731_ _7553_/Q _5988_/A _3960_/C vssd1 vssd1 vccd1 vccd1 _3988_/B sky130_fd_sc_hd__or3_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5667__A1_N _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7481_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4180__A _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6450_ _6568_/A _6471_/B vssd1 vssd1 vccd1 vccd1 _6485_/B sky130_fd_sc_hd__or2_1
X_3662_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__inv_2
X_5401_ hold407/X _4529_/X _5409_/S vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__mux2_1
X_6381_ _3989_/X _6378_/Y _6380_/X _6927_/A vssd1 vssd1 vccd1 vccd1 _6414_/S sky130_fd_sc_hd__a211o_4
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5332_ _4947_/X hold283/X _5338_/S vssd1 vssd1 vccd1 vccd1 _7448_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4450__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5215__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4202__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5263_ hold202/X _5015_/X _5265_/S vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__mux2_1
X_5194_ _5022_/X hold293/X _5194_/S vssd1 vssd1 vccd1 vccd1 _7387_/D sky130_fd_sc_hd__mux2_1
X_4214_ _7424_/Q _7356_/Q _7348_/Q _7328_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4214_/X sky130_fd_sc_hd__mux4_1
X_7002_ _7002_/A _7002_/B vssd1 vssd1 vccd1 vccd1 _7002_/Y sky130_fd_sc_hd__nand2_1
X_4145_ hold8/A input16/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4145_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5083__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4076_ _4039_/C _4057_/X _4075_/Y input15/X _7244_/A vssd1 vssd1 vccd1 vccd1 _4076_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4830__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _5002_/A _4957_/X _4977_/X _4953_/Y _4977_/B vssd1 vssd1 vccd1 vccd1 _4978_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3929_ _7379_/Q _7307_/Q _7299_/Q _7291_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3929_/X sky130_fd_sc_hd__mux4_1
X_6717_ _6718_/A _6718_/B vssd1 vssd1 vccd1 vccd1 _6717_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6648_ _6648_/A _6666_/A _6670_/B _6708_/A vssd1 vssd1 vccd1 vccd1 _6648_/X sky130_fd_sc_hd__and4_2
XFILLER_0_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5543__C1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6579_ _6742_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _6579_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5914__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5125__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4249__B _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4964__S _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5074__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4821__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4888__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5824__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4159__B _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5065__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _5931_/A _5932_/X _5948_/Y _5955_/A vssd1 vssd1 vccd1 vccd1 _5950_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__4812__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4901_ _4199_/B _4900_/Y _6096_/A vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7620_ _7620_/CLK _7620_/D vssd1 vssd1 vccd1 vccd1 _7620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5881_ _5952_/A _5881_/B vssd1 vssd1 vccd1 vccd1 _5881_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6014__B1 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4832_ _4831_/X _4394_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7301_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ hold348/X _4629_/X _4767_/S vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7551_ _7587_/CLK _7551_/D vssd1 vssd1 vccd1 vccd1 _7551_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7482_ _7596_/CLK _7482_/D vssd1 vssd1 vccd1 vccd1 _7482_/Q sky130_fd_sc_hd__dfxtp_1
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__inv_2
XFILLER_0_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6502_ _6503_/B _6503_/C _6611_/A vssd1 vssd1 vccd1 vccd1 _6505_/C sky130_fd_sc_hd__a21oi_2
X_3714_ _6326_/B hold97/X vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6433_ _5568_/B _6432_/S _6434_/B _6710_/A _6656_/A vssd1 vssd1 vccd1 vccd1 _6521_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4879__A1 _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3645_ hold88/X vssd1 vssd1 vccd1 vccd1 _3645_/Y sky130_fd_sc_hd__inv_2
X_6364_ hold92/X hold124/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6364_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout107_A _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5315_ hold419/X _4990_/Y _5319_/S vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__mux2_1
X_6295_ _6295_/A _7020_/B vssd1 vssd1 vccd1 vccd1 _7051_/B sky130_fd_sc_hd__nand2_1
X_5246_ _4996_/X hold506/X _5248_/S vssd1 vssd1 vccd1 vccd1 _5246_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4784__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7160__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5177_ _5357_/A _5393_/A _5321_/B vssd1 vssd1 vccd1 vccd1 _5194_/S sky130_fd_sc_hd__or3_4
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5056__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4128_ _4128_/A _4279_/C _4128_/C vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__and3_1
XANTENNA__7045__A2 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4059_ _4058_/X hold601/X _7241_/S vssd1 vssd1 vccd1 vccd1 _4059_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4803__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5295__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5047__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4723__A _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold508 _7494_/Q vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 _4741_/X vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6180__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5100_ hold619/X _4871_/Y _5112_/S vssd1 vssd1 vccd1 vccd1 _7345_/D sky130_fd_sc_hd__mux2_1
X_6080_ _6153_/A _6080_/B vssd1 vssd1 vccd1 vccd1 _6080_/Y sky130_fd_sc_hd__nor2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4708__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ input28/X _5030_/Y _5031_/S vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5038__A1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6982_ _6935_/A _6799_/A _4037_/X _6971_/X _6981_/X vssd1 vssd1 vccd1 vccd1 _6982_/X
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_50_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7538_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5933_ _5933_/A _5933_/B _5933_/C vssd1 vssd1 vccd1 vccd1 _5933_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4633__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5864_ _5864_/A _5864_/B vssd1 vssd1 vccd1 vccd1 _5866_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ hold182/X _4529_/X _4823_/S vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__mux2_1
X_7603_ _7623_/CLK _7603_/D vssd1 vssd1 vccd1 vccd1 _7603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7534_ _7534_/CLK _7534_/D vssd1 vssd1 vccd1 vccd1 _7534_/Q sky130_fd_sc_hd__dfxtp_1
X_5795_ _7033_/B _7033_/A vssd1 vssd1 vccd1 vccd1 _7069_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4746_ _4745_/X _4685_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7267_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7155__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4779__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7465_ _7485_/CLK _7465_/D vssd1 vssd1 vccd1 vccd1 _7465_/Q sky130_fd_sc_hd__dfxtp_1
X_4677_ _6157_/A _4986_/S vssd1 vssd1 vccd1 vccd1 _4677_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5464__A _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7396_ _7396_/CLK _7396_/D vssd1 vssd1 vccd1 vccd1 _7396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6416_ _6416_/A _6416_/B vssd1 vssd1 vccd1 vccd1 _6419_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6171__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4721__A0 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6347_ _6373_/A _6347_/B vssd1 vssd1 vccd1 vccd1 _7558_/D sky130_fd_sc_hd__and2_1
XANTENNA__5277__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6278_ _6311_/A _6808_/B vssd1 vssd1 vccd1 vccd1 _6949_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5403__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5229_ hold374/X _5038_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4808__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3712__A _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__C _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5029__A1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5358__B _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4960__A0 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6409__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6933__A _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6768__A1 _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4453__A _4460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4600_ _4601_/C vssd1 vssd1 vccd1 vccd1 _4600_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5580_ _6445_/A _5580_/B vssd1 vssd1 vccd1 vccd1 _6437_/A sky130_fd_sc_hd__xnor2_1
X_4531_ _4492_/X hold448/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7253_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7250_ _7485_/CLK _7250_/D vssd1 vssd1 vccd1 vccd1 _7250_/Q sky130_fd_sc_hd__dfxtp_1
Xhold305 _7470_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ _4116_/Y _4459_/X _4461_/X _4113_/Y vssd1 vssd1 vccd1 vccd1 _4462_/X sky130_fd_sc_hd__o211a_1
Xhold316 _4060_/X vssd1 vssd1 vccd1 vccd1 _4061_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold327 _5191_/X vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _7456_/Q vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _4763_/X vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4703__B1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6201_ _3646_/Y _3647_/Y _6207_/S vssd1 vssd1 vccd1 vccd1 _6201_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7181_ _4444_/A _4483_/X _7191_/S vssd1 vssd1 vccd1 vccd1 _7181_/X sky130_fd_sc_hd__mux2_1
X_4393_ _4107_/Y _4390_/X _4391_/Y _4392_/Y _3934_/A vssd1 vssd1 vccd1 vccd1 _4394_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5259__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6132_ hold64/X _6168_/S _6131_/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__a21bo_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _7348_/Q _6356_/B _6062_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6063_/X sky130_fd_sc_hd__a211o_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5223__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5014_ _4101_/A _5034_/B _5032_/B _5013_/Y _4162_/B vssd1 vssd1 vccd1 vccd1 _5014_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6843__A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5967__C1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6965_ _6978_/B _6318_/B _6319_/B _6253_/Y vssd1 vssd1 vccd1 vccd1 _6965_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5459__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _6273_/A _6827_/A _6341_/A vssd1 vssd1 vccd1 vccd1 _5916_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6896_ split4/A _6900_/A vssd1 vssd1 vccd1 vccd1 _6897_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4617__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7184__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5847_ _5723_/A _5802_/C _5845_/Y _5879_/A vssd1 vssd1 vccd1 vccd1 _5847_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_91_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5778_ _7069_/B _5778_/B vssd1 vssd1 vccd1 vccd1 _7033_/A sky130_fd_sc_hd__and2_1
X_4729_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _7176_/B sky130_fd_sc_hd__nor2_4
X_7517_ _7537_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7448_ _7448_/CLK _7448_/D vssd1 vssd1 vccd1 vccd1 _7448_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3840__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3707__A _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7379_ _7379_/CLK _7379_/D vssd1 vssd1 vccd1 vccd1 _7379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4538__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5422__A1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5186__A0 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5816__B _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3831__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A _7544_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4448__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4464__A2 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5661__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6750_ _6773_/A _6773_/B vssd1 vssd1 vccd1 vccd1 _6750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3962_ _6920_/A _3962_/B _3962_/C _3962_/D vssd1 vssd1 vccd1 vccd1 _4140_/B sky130_fd_sc_hd__and4_2
X_5701_ _5701_/A _5701_/B vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__or2_1
XANTENNA__7166__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3893_ _3891_/X _3892_/X _3915_/A vssd1 vssd1 vccd1 vccd1 _3894_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6681_ _6742_/A _6681_/B vssd1 vssd1 vccd1 vccd1 _6723_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5632_ _6691_/A _6871_/A _5629_/Y _5630_/X vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__o22a_1
X_5563_ _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5563_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5218__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3822__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7302_ _7618_/CLK _7302_/D vssd1 vssd1 vccd1 vccd1 _7302_/Q sky130_fd_sc_hd__dfxtp_1
X_4514_ _4930_/S _4513_/X _4512_/X vssd1 vssd1 vccd1 vccd1 _4514_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5494_ _5494_/A _5494_/B vssd1 vssd1 vccd1 vccd1 _5494_/Y sky130_fd_sc_hd__xnor2_1
Xhold102 _5954_/X vssd1 vssd1 vccd1 vccd1 _7497_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _7537_/Q vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _7563_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _6009_/Y vssd1 vssd1 vccd1 vccd1 _7501_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _7278_/Q _7593_/Q _7262_/Q _7486_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4445_/X sky130_fd_sc_hd__mux4_1
Xhold157 _7499_/Q vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _7522_/Q vssd1 vssd1 vccd1 vccd1 _6179_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7233_ _7233_/A _7233_/B _7232_/X vssd1 vssd1 vccd1 vccd1 _7237_/S sky130_fd_sc_hd__or3b_1
Xhold168 _6192_/X vssd1 vssd1 vccd1 vccd1 _7526_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7164_ hold242/X _4679_/X _7166_/S vssd1 vssd1 vccd1 vccd1 _7164_/X sky130_fd_sc_hd__mux2_1
Xhold179 _7223_/X vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
X_4376_ _4672_/B _6089_/B vssd1 vssd1 vccd1 vccd1 _4376_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6115_ _6115_/A vssd1 vssd1 vccd1 vccd1 _6115_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6429__B1 _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7095_/A _7095_/B _5798_/Y vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__or3b_1
X_6046_ _6025_/Y _6043_/Y _6045_/X vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__o21a_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4792__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6573__A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4093__A _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6948_ _6949_/A _6948_/B vssd1 vssd1 vccd1 vccd1 _6948_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__7157__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6879_ _6868_/Y _6870_/X _6880_/A vssd1 vssd1 vccd1 vccd1 _6879_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6904__A1 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5917__A _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5636__B _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3813__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5128__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6380__A2 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6117__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6132__A2 _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7093__B1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6483__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3900__A _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7148__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6108__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4230_ _7442_/Q _7434_/Q _7418_/Q _7410_/Q _7452_/Q _7453_/Q vssd1 vssd1 vccd1 vccd1
+ _4230_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5562__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4161_ _4751_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _7212_/A sky130_fd_sc_hd__and2_2
XANTENNA__5882__A1 _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4092_ _4748_/A _4825_/B vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5398__A0 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6802_ _6802_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6802_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _7123_/A _4945_/B _4942_/B _3939_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4994_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4296__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3945_ _3933_/Y _3935_/X _3944_/X _3788_/X vssd1 vssd1 vccd1 vccd1 _5974_/C sky130_fd_sc_hd__a31oi_4
XFILLER_0_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6733_ _6869_/A _6735_/B _6742_/B _6871_/A vssd1 vssd1 vccd1 vccd1 _6734_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7139__A1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6664_ _6773_/A _6710_/B vssd1 vssd1 vccd1 vccd1 _6756_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _4862_/A _6039_/A vssd1 vssd1 vccd1 vccd1 _4867_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout137_A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5615_ _5615_/A _5615_/B _6462_/B _6448_/A vssd1 vssd1 vccd1 vccd1 _5621_/D sky130_fd_sc_hd__nor4b_1
XANTENNA__4360__B _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6595_ _6603_/A _6603_/B _6596_/B vssd1 vssd1 vccd1 vccd1 _6643_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5546_ _5854_/C _5546_/B vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__nand2_1
X_5477_ _5483_/B _5482_/A _5476_/B _5458_/Y vssd1 vssd1 vccd1 vccd1 _5477_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6568__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7163__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7216_ _7215_/X _4394_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7617_/D sky130_fd_sc_hd__mux2_1
X_4428_ _4428_/A _4428_/B vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4220__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4359_ _4357_/X _4358_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__mux2_1
X_7147_ _7127_/X _7146_/Y _6413_/S vssd1 vssd1 vccd1 vccd1 _7147_/X sky130_fd_sc_hd__o21a_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _7078_/A _7078_/B _7078_/C _7078_/D vssd1 vssd1 vccd1 vccd1 _7078_/X sky130_fd_sc_hd__or4_1
XANTENNA__7075__B1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7424_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6029_ _6922_/C _6023_/X _6024_/X _6025_/Y _6028_/X vssd1 vssd1 vccd1 vccd1 _6029_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5625__B2 _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5625__A1 _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout85 _4147_/X vssd1 vssd1 vccd1 vccd1 _4529_/S sky130_fd_sc_hd__buf_4
XFILLER_0_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout96 _6022_/B vssd1 vssd1 vccd1 vccd1 _6375_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4270__B _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6353__A2 _5811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4364__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4211__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3630__A _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4164__C _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5919__A2 _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4052__A0 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _6223_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _4122_/C sky130_fd_sc_hd__or2_4
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3661_ _6920_/A vssd1 vssd1 vccd1 vccd1 _5132_/A sky130_fd_sc_hd__inv_2
X_5400_ _4443_/X hold440/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7486_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3789__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6380_ _7230_/A _5990_/A _6415_/B _6379_/X vssd1 vssd1 vccd1 vccd1 _6380_/X sky130_fd_sc_hd__a31o_1
X_5331_ hold282/X _4964_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4450__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5262_ _5261_/X _4973_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4202__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7001_ _6900_/A _6988_/A _6999_/Y _7000_/X _3949_/Y vssd1 vssd1 vccd1 vccd1 _7001_/X
+ sky130_fd_sc_hd__o221a_1
X_5193_ hold292/X _5038_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3866__B1 _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4213_ _7320_/Q _7336_/Q _7312_/Q _7448_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4213_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4144_ _4139_/Y _4142_/X _4846_/A vssd1 vssd1 vccd1 vccd1 _4144_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__7057__B1 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4075_ _6871_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _4075_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7012__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6851__A _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7158__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4977_ _4977_/A _4977_/B vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__and2_1
X_6716_ _6716_/A _6718_/B vssd1 vssd1 vccd1 vccd1 _6716_/Y sky130_fd_sc_hd__nor2_1
X_3928_ _7363_/Q _3928_/B vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__and2_1
XFILLER_0_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3859_ _3827_/S _3857_/X _3858_/X vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__a21oi_4
X_6647_ _6840_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6708_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578_ _6580_/B vssd1 vssd1 vccd1 vccd1 _6578_/Y sky130_fd_sc_hd__inv_2
X_5529_ _5854_/C _5546_/B vssd1 vssd1 vccd1 vccd1 _5529_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5914__B _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5406__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7048__B1 _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5824__B _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output50_A _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5051__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _4902_/B _4900_/B vssd1 vssd1 vccd1 vccd1 _4900_/Y sky130_fd_sc_hd__xnor2_1
X_5880_ _5879_/A split1/X _5877_/X _5879_/X vssd1 vssd1 vccd1 vccd1 _5881_/B sky130_fd_sc_hd__o2bb2a_1
X_4831_ hold221/X _4434_/Y _4843_/S vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4762_ _4761_/X _4538_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7272_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6970__C1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7550_ _7599_/CLK _7550_/D vssd1 vssd1 vccd1 vccd1 _7550_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5773__B1 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7481_ _7481_/CLK _7481_/D vssd1 vssd1 vccd1 vccd1 _7481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4693_ _3668_/Y _4692_/X _4689_/X vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__a21oi_2
X_6501_ _6503_/B _6503_/C vssd1 vssd1 vccd1 vccd1 _6501_/X sky130_fd_sc_hd__and2_1
X_3713_ _6326_/B hold97/A vssd1 vssd1 vccd1 vccd1 _3716_/B sky130_fd_sc_hd__and2_2
XFILLER_0_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3644_ _3644_/A vssd1 vssd1 vccd1 vccd1 _3644_/Y sky130_fd_sc_hd__inv_2
X_6432_ _5565_/B _6431_/X _6432_/S vssd1 vssd1 vccd1 vccd1 _6434_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5226__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6363_ _6373_/A _6363_/B vssd1 vssd1 vccd1 vccd1 _7562_/D sky130_fd_sc_hd__and2_1
XFILLER_0_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5314_ hold530/X _4947_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _7440_/D sky130_fd_sc_hd__mux2_1
X_6294_ _7019_/A _7019_/B vssd1 vssd1 vccd1 vccd1 _7020_/B sky130_fd_sc_hd__or2_1
X_5245_ hold505/X _5015_/X _5247_/S vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5750__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5176_ _5175_/X _4685_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7379_/D sky130_fd_sc_hd__mux2_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4366__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4127_ _4267_/C _4267_/D _4127_/C vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__and3_1
X_4058_ _4039_/C _4056_/X _4057_/X input10/X _7244_/A vssd1 vssd1 vccd1 vccd1 _4058_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6581__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4319__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5819__B2 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5660__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3925__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6922__C _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4215__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold509 _5883_/X vssd1 vssd1 vccd1 vccd1 _7494_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5046__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7172__A1_N _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _4930_/S _5024_/X _5029_/X vssd1 vssd1 vccd1 vccd1 _5030_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3916__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ _7078_/A _6981_/B _6981_/C _6975_/X vssd1 vssd1 vccd1 vccd1 _6981_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4341__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4797__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5932_ _5933_/A _5933_/B _5933_/C vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863_ _5864_/A _5864_/B vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4549__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4814_ hold281/X _4443_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7294_/D sky130_fd_sc_hd__mux2_1
X_7602_ _7608_/CLK _7602_/D vssd1 vssd1 vccd1 vccd1 _7602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5794_ _5792_/A _5792_/B _5793_/X vssd1 vssd1 vccd1 vccd1 _7033_/B sky130_fd_sc_hd__a21boi_1
X_4745_ hold215/X _4719_/Y _4745_/S vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7533_ _7534_/CLK _7533_/D vssd1 vssd1 vccd1 vccd1 _7533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7464_ _7592_/CLK _7464_/D vssd1 vssd1 vccd1 vccd1 _7464_/Q sky130_fd_sc_hd__dfxtp_1
X_4676_ _4676_/A _4713_/S vssd1 vssd1 vccd1 vccd1 _4676_/Y sky130_fd_sc_hd__xnor2_1
X_7395_ _7403_/CLK _7395_/D vssd1 vssd1 vccd1 vccd1 _7395_/Q sky130_fd_sc_hd__dfxtp_1
X_6415_ _6415_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6416_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6346_ _6413_/S _6415_/A _6415_/B _6220_/B _4084_/A vssd1 vssd1 vccd1 vccd1 _6347_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4795__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5480__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6277_ _7109_/B vssd1 vssd1 vccd1 vccd1 _7110_/A sky130_fd_sc_hd__inv_2
XANTENNA__4485__A0 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5228_ hold384/X _4996_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _7402_/D sky130_fd_sc_hd__mux2_1
X_5159_ _7211_/B _5375_/C _5159_/C vssd1 vssd1 vccd1 vccd1 _5176_/S sky130_fd_sc_hd__and3_4
XANTENNA__4096__A _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__D _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6226__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4332__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3874__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4399__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4712__A1 _7343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3903__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6465__A1 _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4476__B1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6217__A1 _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4323__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4779__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5268__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5565__A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ hold447/X _4529_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4530_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6160__S _6160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold306 _7615_/Q vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _5024_/S _4455_/X _4460_/Y _4930_/S vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__a211o_1
Xhold317 _4064_/X vssd1 vssd1 vccd1 vccd1 _7343_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold339 _5341_/X vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _7285_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
X_7180_ _7179_/X _4394_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7601_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6200_ _6218_/A _6200_/B vssd1 vssd1 vccd1 vccd1 _7534_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4392_ _6111_/A _3901_/B _4107_/Y vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__o21ai_1
X_6131_ _6374_/A _6129_/X _6130_/X _6168_/S _6123_/X vssd1 vssd1 vccd1 vccd1 _6131_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6356_/B _6062_/B vssd1 vssd1 vccd1 vccd1 _6062_/Y sky130_fd_sc_hd__nor2_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5013_ _5012_/A _5012_/B _5034_/B vssd1 vssd1 vccd1 vccd1 _5013_/Y sky130_fd_sc_hd__a21oi_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4644__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6964_ _7123_/A _6922_/B _6981_/C vssd1 vssd1 vccd1 vccd1 _6964_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__7020__A _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout167_A _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6895_ _7129_/A _7085_/A _7085_/B _6893_/Y _6894_/Y vssd1 vssd1 vccd1 vccd1 split4/A
+ sky130_fd_sc_hd__o311a_4
X_5915_ _7123_/A _6844_/A vssd1 vssd1 vccd1 vccd1 _5958_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5178__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5846_ _5723_/A _5802_/C _5845_/Y vssd1 vssd1 vccd1 vccd1 _5877_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4617__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7166__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5777_ _5777_/A _5777_/B _5777_/C vssd1 vssd1 vccd1 vccd1 _5778_/B sky130_fd_sc_hd__or3_1
X_4728_ _4964_/S _4728_/B _4750_/B vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__and3_2
X_7516_ _7537_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7447_ _4004_/A _7447_/D vssd1 vssd1 vccd1 vccd1 _7447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4659_ _6844_/A _4658_/A _4658_/Y _4116_/Y vssd1 vssd1 vccd1 vccd1 _4659_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3707__B _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _7378_/CLK _7378_/D vssd1 vssd1 vccd1 vccd1 _7378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _6329_/A _6329_/B vssd1 vssd1 vccd1 vccd1 _6331_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4305__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5816__C _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5324__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3633__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5110__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5661__A2 _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7476_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5413__A2 _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3961_ _4036_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _3962_/D sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5700_ _5700_/A _5700_/B vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__nor2_1
X_3892_ _7403_/Q _7395_/Q _7371_/Q _7387_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3892_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6680_ _6742_/A _6681_/B vssd1 vssd1 vccd1 vccd1 _6680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5631_ _5630_/X _6742_/A _6690_/A _5631_/D vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__and4b_1
XFILLER_0_79_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5562_ _6710_/A _5591_/B vssd1 vssd1 vccd1 vccd1 _5579_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7301_ _7476_/CLK _7301_/D vssd1 vssd1 vccd1 vccd1 _7301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4513_ _6123_/B _4507_/X _6096_/A vssd1 vssd1 vccd1 vccd1 _4513_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5493_ _5493_/A _5493_/B vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__nand2_1
Xhold114 _6205_/X vssd1 vssd1 vccd1 vccd1 _6206_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold125 _6364_/X vssd1 vssd1 vccd1 vccd1 _6365_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _7580_/Q vssd1 vssd1 vccd1 vccd1 _6420_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ _7232_/A _7232_/B _7232_/C vssd1 vssd1 vccd1 vccd1 _7232_/X sky130_fd_sc_hd__and3_1
X_4444_ _4444_/A _4493_/C vssd1 vssd1 vccd1 vccd1 _4444_/Y sky130_fd_sc_hd__xnor2_1
Xhold158 _5973_/X vssd1 vssd1 vccd1 vccd1 _7499_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _6180_/X vssd1 vssd1 vccd1 vccd1 _7522_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold136 _7560_/Q vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5234__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7163_ hold467/X _4589_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7596_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_95_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4375_ _4667_/B _4370_/X _4374_/X vssd1 vssd1 vccd1 vccd1 _6089_/B sky130_fd_sc_hd__a21oi_4
Xhold169 _7312_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_6114_ _4460_/B _6116_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6115_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6429__A1 _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _5798_/A _5798_/C _7073_/A vssd1 vssd1 vccd1 vccd1 _7095_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5101__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6045_ _7346_/Q _6356_/B _6044_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__a211o_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4860__B1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4093__B _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6947_ _7020_/A _6974_/C _6945_/Y _6946_/Y vssd1 vssd1 vccd1 vccd1 _6952_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6878_ _6939_/A _6877_/B _6875_/X vssd1 vssd1 vccd1 vccd1 _6968_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5168__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6904__A2 _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5829_ _5829_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5831_/B sky130_fd_sc_hd__xor2_1
XANTENNA__5917__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5409__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3718__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5144__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold663_A _7587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7148__A2 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5331__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5054__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4160_ _4963_/S _4158_/X _4159_/X _4964_/S vssd1 vssd1 vccd1 vccd1 _4827_/B sky130_fd_sc_hd__o211a_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7084__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4517__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4091_ hold97/A input8/X _5022_/A vssd1 vssd1 vccd1 vccd1 _4825_/B sky130_fd_sc_hd__mux2_4
X_6801_ _6801_/A1 _6774_/Y _6802_/A _6765_/X vssd1 vssd1 vccd1 vccd1 _6801_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _6084_/A _4993_/B vssd1 vssd1 vccd1 vccd1 _4993_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3944_ _3937_/Y _3939_/X _3944_/C _3944_/D vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4070__A1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6732_ _6742_/A _6732_/B vssd1 vssd1 vccd1 vccd1 _6732_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3875_ _3827_/S _3874_/X _3871_/X vssd1 vssd1 vccd1 vccd1 _6039_/A sky130_fd_sc_hd__a21oi_4
X_6663_ _6773_/A _6710_/B vssd1 vssd1 vccd1 vccd1 _6663_/X sky130_fd_sc_hd__and2_4
XANTENNA__5229__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5614_ _5620_/B _5614_/B vssd1 vssd1 vccd1 vccd1 _6448_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6898__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6594_ _6593_/B _6574_/Y _6613_/B _6592_/Y _6567_/A vssd1 vssd1 vccd1 vccd1 _6603_/B
+ sky130_fd_sc_hd__o311ai_4
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5545_ _5583_/B _5585_/A _5533_/Y vssd1 vssd1 vccd1 vccd1 _5545_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5476_ _5482_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5489_/A sky130_fd_sc_hd__and2_1
XFILLER_0_41_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7215_ hold380/X _4434_/Y _7227_/S vssd1 vssd1 vccd1 vccd1 _7215_/X sky130_fd_sc_hd__mux2_1
X_4427_ _6098_/B _4320_/A _4383_/Y vssd1 vssd1 vccd1 vccd1 _4428_/B sky130_fd_sc_hd__o21a_1
X_7146_ _4031_/B _7144_/X _7145_/X vssd1 vssd1 vccd1 vccd1 _7146_/Y sky130_fd_sc_hd__a21oi_1
X_4358_ _7402_/Q _7394_/Q _7370_/Q _7386_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4358_/X sky130_fd_sc_hd__mux4_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _6911_/B _4290_/B _6220_/C _4290_/D vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__or4_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _7020_/A _7071_/X _7072_/Y _7076_/X _7068_/X vssd1 vssd1 vccd1 vccd1 _7078_/D
+ sky130_fd_sc_hd__a311o_1
X_6028_ _6328_/A _4999_/B _6166_/B _4122_/C vssd1 vssd1 vccd1 vccd1 _6028_/X sky130_fd_sc_hd__o211a_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4551__B _4879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout86 _6166_/B vssd1 vssd1 vccd1 vccd1 _6157_/B sky130_fd_sc_hd__buf_4
Xfanout97 _3711_/X vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5313__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4279__A _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5849__C1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3875__A1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5049__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3660_ hold76/A vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__inv_2
XANTENNA__3789__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4888__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5330_ _4921_/X _5329_/X _5338_/S vssd1 vssd1 vccd1 vccd1 _7447_/D sky130_fd_sc_hd__mux2_1
X_5261_ hold390/X _4990_/Y _5265_/S vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4212_ _4688_/S _4212_/B vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4189__A _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7000_ _6869_/B split4/X _7043_/S vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__a21o_1
X_5192_ _4996_/X hold327/X _5194_/S vssd1 vssd1 vccd1 vccd1 _7386_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3866__A1 _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7378_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4512__C1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4143_ _4139_/Y _4142_/X _4846_/A vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__o21a_1
XANTENNA__7057__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _4073_/X hold524/X _7249_/S vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5240__A0 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4579__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4976_ _5008_/A _4976_/B _5001_/A _4980_/B vssd1 vssd1 vccd1 vccd1 _4976_/X sky130_fd_sc_hd__or4_1
X_6715_ _6701_/Y _6714_/Y split7/A vssd1 vssd1 vccd1 vccd1 _6718_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3927_ _3925_/X _3926_/X _7362_/Q vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3858_ _3915_/A _3852_/X _3854_/X _7363_/Q vssd1 vssd1 vccd1 vccd1 _3858_/X sky130_fd_sc_hd__o211a_1
X_6646_ _6773_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3789_ _7282_/Q _7597_/Q _7266_/Q _7490_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3789_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4798__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6577_ _6518_/B _6576_/X _7090_/B vssd1 vssd1 vccd1 vccd1 _6580_/B sky130_fd_sc_hd__mux2_1
XANTENNA__6579__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5528_ _5503_/B _5527_/Y _5528_/S vssd1 vssd1 vccd1 vccd1 _5546_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6099__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3715__B _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6298__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5459_ _5854_/C _5459_/B vssd1 vssd1 vccd1 vccd1 _5483_/B sky130_fd_sc_hd__nand2_1
Xfanout210 _4846_/A vssd1 vssd1 vccd1 vccd1 _6345_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7129_ _7129_/A _7129_/B vssd1 vssd1 vccd1 vccd1 _7130_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4806__A0 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7220__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5658__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5096__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5332__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3641__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5470__B1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6952__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4830_ hold579/X _4111_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7300_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5568__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4761_ hold445/X _4580_/X _4767_/S vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5773__B2 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5773__A1 _6874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7480_ _7483_/CLK _7480_/D vssd1 vssd1 vccd1 vccd1 _7480_/Q sky130_fd_sc_hd__dfxtp_1
X_4692_ _4690_/X _4691_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4692_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4981__C1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6500_ _6521_/A _6521_/D _6498_/Y vssd1 vssd1 vccd1 vccd1 _6503_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3712_ _4037_/A _3712_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3643_ _3643_/A vssd1 vssd1 vccd1 vccd1 _3643_/Y sky130_fd_sc_hd__inv_2
X_6431_ _6431_/A _6431_/B vssd1 vssd1 vccd1 vccd1 _6431_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6362_ _7570_/Q hold132/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6362_/X sky130_fd_sc_hd__mux2_1
X_5313_ hold529/X _4964_/X _5319_/S vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6293_ _6249_/A _6988_/B _6279_/B vssd1 vssd1 vccd1 vccd1 _7019_/B sky130_fd_sc_hd__a21o_1
X_5244_ _4973_/X _5243_/X _5248_/S vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__mux2_1
X_5175_ hold322/X _4719_/Y _5175_/S vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5242__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A _7342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4126_ _6920_/A _4846_/A _4128_/A vssd1 vssd1 vccd1 vccd1 _4127_/C sky130_fd_sc_hd__and3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__or2_1
XANTENNA__6581__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7202__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4016__A1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _5008_/A _4956_/X _4958_/X _4952_/X vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6629_ _6629_/A _6629_/B _6629_/C vssd1 vssd1 vccd1 vccd1 _6629_/X sky130_fd_sc_hd__and3_1
XFILLER_0_15_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5660__B _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3925__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5152__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4557__A _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4991__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A0 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_7__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5327__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5062__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3916__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__A1 _7454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6980_ _6973_/X _6979_/X _7043_/S vssd1 vssd1 vccd1 vccd1 _6981_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5931_ _5931_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5933_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4341__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5862_ _7109_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5864_/B sky130_fd_sc_hd__xnor2_1
X_4813_ hold280/X _4483_/X _4823_/S vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__mux2_1
X_7601_ _7617_/CLK _7601_/D vssd1 vssd1 vccd1 vccd1 _7601_/Q sky130_fd_sc_hd__dfxtp_2
X_5793_ _7002_/A _7002_/B vssd1 vssd1 vccd1 vccd1 _5793_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _4743_/X _4637_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7266_/D sky130_fd_sc_hd__mux2_1
X_7532_ _7534_/CLK _7532_/D vssd1 vssd1 vccd1 vccd1 _7532_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3852__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7463_ _7596_/CLK _7463_/D vssd1 vssd1 vccd1 vccd1 _7463_/Q sky130_fd_sc_hd__dfxtp_1
X_4675_ _4625_/B _4625_/C _4624_/B _4625_/A vssd1 vssd1 vccd1 vccd1 _4713_/S sky130_fd_sc_hd__a211o_1
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7394_ _7485_/CLK _7394_/D vssd1 vssd1 vccd1 vccd1 _7394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6414_ _6413_/X hold315/X _6414_/S vssd1 vssd1 vccd1 vccd1 _7579_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6857__A _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6345_ _6345_/A _6345_/B vssd1 vssd1 vccd1 vccd1 _7557_/D sky130_fd_sc_hd__and2_1
X_6276_ _6238_/X _6276_/B vssd1 vssd1 vccd1 vccd1 _7109_/B sky130_fd_sc_hd__and2b_2
X_5227_ hold383/X _5015_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6068__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5158_ _5022_/X hold548/X _5158_/S vssd1 vssd1 vccd1 vccd1 _7371_/D sky130_fd_sc_hd__mux2_1
X_5089_ hold163/X _4990_/Y _5093_/S vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__mux2_1
X_4109_ _4103_/A _3937_/A _4106_/X vssd1 vssd1 vccd1 vccd1 _4109_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4332__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5147__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4399__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4986__S _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4712__A2 _4707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5425__B1 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4323__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5057__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold307 _7270_/Q vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
X_4460_ _5024_/S _4460_/B vssd1 vssd1 vccd1 vccd1 _4460_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6689__C1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold318 _7416_/Q vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _7309_/Q vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_4391_ _6874_/A _4440_/A vssd1 vssd1 vccd1 vccd1 _4391_/Y sky130_fd_sc_hd__nor2_1
X_6130_ _6130_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6130_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6061_/A vssd1 vssd1 vccd1 vccd1 _6061_/Y sky130_fd_sc_hd__inv_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5012_ _5012_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__or2_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5416__B1 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5967__B2 _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5967__A1 _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6963_ _6872_/A _6911_/A _7098_/A _6962_/X vssd1 vssd1 vccd1 vccd1 _6981_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6894_ _6840_/A _6840_/B _6845_/A vssd1 vssd1 vccd1 vccd1 _6894_/Y sky130_fd_sc_hd__o21ai_1
X_5914_ _7123_/A _6844_/A vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__and2_1
X_5845_ _5877_/A _5845_/B vssd1 vssd1 vccd1 vccd1 _5845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6916__B1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3825__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6392__A1 _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5776_ _5777_/B _5777_/C _5777_/A vssd1 vssd1 vccd1 vccd1 _7069_/B sky130_fd_sc_hd__o21ai_1
X_4727_ _7211_/B _7150_/B _7175_/B vssd1 vssd1 vccd1 vccd1 _4746_/S sky130_fd_sc_hd__and3_4
X_7515_ _7538_/CLK hold81/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
X_7446_ _7446_/CLK _7446_/D vssd1 vssd1 vccd1 vccd1 _7446_/Q sky130_fd_sc_hd__dfxtp_1
X_4658_ _4658_/A _4658_/B vssd1 vssd1 vccd1 vccd1 _4658_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4155__B1 _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7377_ _7620_/CLK _7377_/D vssd1 vssd1 vccd1 vccd1 _7377_/Q sky130_fd_sc_hd__dfxtp_1
X_4589_ _4685_/A _4589_/B vssd1 vssd1 vccd1 vccd1 _4589_/X sky130_fd_sc_hd__or2_4
XANTENNA__5491__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6328_ _6328_/A _6328_/B vssd1 vssd1 vccd1 vccd1 _6919_/B sky130_fd_sc_hd__nand2_1
X_6259_ _6974_/B _6259_/B vssd1 vssd1 vccd1 vccd1 _6949_/A sky130_fd_sc_hd__nand2_2
XANTENNA__4305__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4554__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4630__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3816__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4570__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5816__D _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4697__A1 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4729__B _4827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3960_ _6225_/A _6223_/A _3960_/C vssd1 vssd1 vccd1 vccd1 _6220_/C sky130_fd_sc_hd__or3_4
XANTENNA__6960__A _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4621__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3891_ _7443_/Q _7435_/Q _7419_/Q _7411_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3891_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5576__A _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5630_ _6802_/A _6808_/A _6637_/A _6702_/A vssd1 vssd1 vccd1 vccd1 _5630_/X sky130_fd_sc_hd__and4_1
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5561_ _5577_/A _5561_/A2 _5561_/A3 _5559_/Y vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7300_ _7476_/CLK _7300_/D vssd1 vssd1 vccd1 vccd1 _7300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5492_ _6568_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5493_/B sky130_fd_sc_hd__nand2_1
X_4512_ _6869_/A _4658_/A _4511_/X _5008_/A vssd1 vssd1 vccd1 vccd1 _4512_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold126 _7564_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _6420_/Y vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
X_7231_ _7231_/A _7231_/B _7231_/C _7231_/D vssd1 vssd1 vccd1 vccd1 _7232_/C sky130_fd_sc_hd__and4_1
Xhold115 _7531_/Q vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4443_ _5022_/A _4443_/B vssd1 vssd1 vccd1 vccd1 _4443_/X sky130_fd_sc_hd__or2_4
Xhold159 _7538_/Q vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 _6358_/X vssd1 vssd1 vccd1 vccd1 _6359_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5885__B1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 _7599_/Q vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__clkbuf_4
X_7162_ hold466/X _4629_/X _7166_/S vssd1 vssd1 vccd1 vccd1 _7162_/X sky130_fd_sc_hd__mux2_1
X_4374_ _4667_/B _4374_/B vssd1 vssd1 vccd1 vccd1 _4374_/X sky130_fd_sc_hd__and2b_1
XANTENNA__6200__A _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6113_ _6112_/X hold72/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__mux2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6429__A2 _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7091_/X _7092_/X _6900_/A vssd1 vssd1 vccd1 vccd1 _7093_/X sky130_fd_sc_hd__a21o_1
X_6044_ _6356_/B _6044_/B vssd1 vssd1 vccd1 vccd1 _6044_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5637__B1 _7040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4860__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6946_ _7070_/A _6978_/A vssd1 vssd1 vccd1 vccd1 _6946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4093__C _4846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5486__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6877_ _6875_/X _6877_/B vssd1 vssd1 vccd1 vccd1 _6939_/B sky130_fd_sc_hd__and2b_1
XANTENNA__3966__A3 _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4390__A _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5828_ _5829_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5759_ _5769_/A _5760_/B vssd1 vssd1 vccd1 vccd1 _5797_/A sky130_fd_sc_hd__or2_1
XANTENNA__3718__B _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4223__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7429_ _7449_/CLK _7429_/D vssd1 vssd1 vccd1 vccd1 _7429_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4679__A1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout92_A _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 _6799_/A vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5628__B1 _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6780__A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5335__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4214__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output73_A _7522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4517__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4090_ _5805_/A input9/X _5022_/A vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4842__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5070__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6690__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6800_ _6790_/S _6796_/Y _6797_/Y _6799_/A vssd1 vssd1 vccd1 vccd1 _6859_/B sky130_fd_sc_hd__a211o_1
X_4992_ _4991_/X _4973_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _4992_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3943_ _6148_/A _6139_/A _6130_/A _3943_/D vssd1 vssd1 vccd1 vccd1 _3944_/D sky130_fd_sc_hd__and4_1
XFILLER_0_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6731_ _6742_/B vssd1 vssd1 vccd1 vccd1 _6732_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3874_ _3872_/X _3873_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__mux2_1
X_6662_ _6606_/B _6659_/Y _6661_/X _6642_/Y vssd1 vssd1 vccd1 vccd1 _6710_/B sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5613_ _5615_/B _6451_/B _5612_/X _5597_/X vssd1 vssd1 vccd1 vccd1 _5620_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6593_ _6593_/A _6593_/B vssd1 vssd1 vccd1 vccd1 _6608_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5544_ _5542_/Y _5543_/X _5541_/Y vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5475_ _5504_/A _5465_/B _5472_/B _5499_/B _5470_/Y vssd1 vssd1 vccd1 vccd1 _5476_/B
+ sky130_fd_sc_hd__a221o_1
X_7214_ hold166/X _4111_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7616_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4426_ _4477_/B _4477_/C vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__nor2_1
X_7145_ _6093_/A _5804_/C _4029_/Y _6166_/A _6326_/C vssd1 vssd1 vccd1 vccd1 _7145_/X
+ sky130_fd_sc_hd__a221o_1
X_4357_ _7442_/Q _7434_/Q _7418_/Q _7410_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4357_/X sky130_fd_sc_hd__mux4_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4288_ _4667_/B _4283_/X _4287_/X vssd1 vssd1 vccd1 vccd1 _6098_/B sky130_fd_sc_hd__a21oi_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7043_/S _7073_/Y _7074_/X _7075_/Y _3705_/X vssd1 vssd1 vccd1 vccd1 _7076_/X
+ sky130_fd_sc_hd__o221a_1
X_6027_ _6166_/B vssd1 vssd1 vccd1 vccd1 _6027_/Y sky130_fd_sc_hd__inv_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4833__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6311_/A _6926_/Y _6928_/X _6917_/Y _6373_/A vssd1 vssd1 vccd1 vccd1 _7583_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3729__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout87 _6026_/X vssd1 vssd1 vccd1 vccd1 _6166_/B sky130_fd_sc_hd__buf_4
Xfanout98 _3711_/X vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__buf_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5010__A1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5155__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold490 _5165_/X vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4824__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6015__A _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5854__A _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5065__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5260_ hold319/X _4947_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _7416_/D sky130_fd_sc_hd__mux2_1
X_4211_ _7400_/Q _7392_/Q _7368_/Q _7384_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4212_/B sky130_fd_sc_hd__mux4_1
X_5191_ hold326/X _5015_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5068__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4142_ _4267_/D _4142_/B vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__and2_1
XANTENNA__7057__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4073_ _7244_/A input14/X _4039_/C _4072_/X vssd1 vssd1 vccd1 vccd1 _4073_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4815__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7396_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ _5002_/A _4974_/B _4949_/X _4977_/B vssd1 vssd1 vccd1 vccd1 _4980_/B sky130_fd_sc_hd__a22o_1
X_3926_ _7483_/Q _7471_/Q _7463_/Q _7257_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3926_/X sky130_fd_sc_hd__mux4_1
X_6714_ _6714_/A _6714_/B vssd1 vssd1 vccd1 vccd1 _6714_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3857_ _3855_/X _3856_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6645_ _6773_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6576_ _6576_/A _6576_/B vssd1 vssd1 vccd1 vccd1 _6576_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ _3962_/B _3771_/Y _3772_/X _3777_/X _3787_/X vssd1 vssd1 vccd1 vccd1 _3788_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5527_ _5527_/A _5527_/B vssd1 vssd1 vccd1 vccd1 _5527_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3715__C hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5458_ _5854_/C _5459_/B vssd1 vssd1 vccd1 vccd1 _5458_/Y sky130_fd_sc_hd__nor2_1
X_5389_ hold396/X _4679_/X _5391_/S vssd1 vssd1 vccd1 vccd1 _5389_/X sky130_fd_sc_hd__mux2_1
Xfanout200 _4709_/S1 vssd1 vssd1 vccd1 vccd1 _4706_/S1 sky130_fd_sc_hd__buf_6
X_4409_ _4269_/A _4403_/Y _4408_/X _4658_/A vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout211 input44/X vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__buf_6
XANTENNA__4827__B _4827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7128_ _6887_/A _6887_/B _6845_/A vssd1 vssd1 vccd1 vccd1 _7129_/B sky130_fd_sc_hd__a21oi_1
X_7059_ _7054_/X _7055_/X _7058_/Y _6220_/C vssd1 vssd1 vccd1 vccd1 _7059_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3731__B _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5939__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5658__B _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4665__S0 _7340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3867__A1_N _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3893__S _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4417__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6192__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5298__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6495__B1 _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3922__A _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5222__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ hold470/X _4492_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7271_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4430__C1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5773__A2 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4691_ _7275_/Q _7615_/Q _7607_/Q _7623_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4691_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3711_ _4037_/A _3712_/B vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__and2_1
XFILLER_0_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3642_ hold97/X vssd1 vssd1 vccd1 vccd1 _6421_/B sky130_fd_sc_hd__inv_2
X_6430_ _6430_/A _6430_/B vssd1 vssd1 vccd1 vccd1 _6431_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6183__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6361_ _6373_/A _6361_/B vssd1 vssd1 vccd1 vccd1 _7561_/D sky130_fd_sc_hd__and2_1
X_5312_ _5311_/X _4921_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _7439_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5289__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6292_ _6319_/A _6959_/B _6264_/A vssd1 vssd1 vccd1 vccd1 _6988_/B sky130_fd_sc_hd__o21ba_1
X_5243_ hold498/X _4990_/Y _5247_/S vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5174_ _5173_/X _4637_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7378_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5750__C _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4125_ _6328_/A _5985_/B _4124_/B vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__or3b_1
X_4056_ _6220_/C _4056_/B vssd1 vssd1 vccd1 vccd1 _4056_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4016__A2 _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4958_ _5001_/A _4951_/Y _4955_/Y _4957_/X _4954_/X vssd1 vssd1 vccd1 vccd1 _4958_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3909_ _3827_/S _3907_/X _3908_/Y _3903_/Y vssd1 vssd1 vccd1 vccd1 _6120_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4889_ hold330/X _4871_/Y _5040_/S vssd1 vssd1 vccd1 vccd1 _7309_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6628_ _6628_/A split9/X vssd1 vssd1 vccd1 vccd1 _6629_/C sky130_fd_sc_hd__or2_1
XANTENNA__6174__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3726__B _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6559_ _6494_/Y _6558_/Y _7090_/B vssd1 vssd1 vccd1 vccd1 _6561_/B sky130_fd_sc_hd__mux2_2
XANTENNA__3742__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4660__C1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6401__A0 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6165__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6704__A1 _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4715__A0 _6166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5912__C1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5343__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5930_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5931_/B sky130_fd_sc_hd__and2_1
XANTENNA__7196__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7600_ _7617_/CLK _7600_/D vssd1 vssd1 vccd1 vccd1 _7600_/Q sky130_fd_sc_hd__dfxtp_2
X_5861_ _5861_/A _5861_/B vssd1 vssd1 vccd1 vccd1 _5862_/B sky130_fd_sc_hd__nor2_1
X_4812_ _4811_/X _4394_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7293_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6943__A1 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5792_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _7002_/B sky130_fd_sc_hd__xnor2_1
X_4743_ hold203/X _4679_/X _4745_/S vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7531_ _7582_/CLK _7531_/D vssd1 vssd1 vccd1 vccd1 _7531_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3852__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7462_ _7596_/CLK _7462_/D vssd1 vssd1 vccd1 vccd1 _7462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6156__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4674_ _4674_/A _4674_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__and2_1
X_6413_ input38/X _6412_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6413_/X sky130_fd_sc_hd__mux2_1
X_7393_ _7441_/CLK _7393_/D vssd1 vssd1 vccd1 vccd1 _7393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6344_ _6343_/X _6301_/A _6344_/S vssd1 vssd1 vccd1 vccd1 _6345_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5880__A1_N _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6275_ _7109_/A _6275_/B vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__nand2_2
X_5226_ _5225_/X _4973_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5157_ hold547/X _5038_/X _5157_/S vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__mux2_1
X_5088_ hold333/X _4947_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _7336_/D sky130_fd_sc_hd__mux2_1
X_4108_ _6261_/A _4440_/A _4389_/B _4104_/X vssd1 vssd1 vccd1 vccd1 _4108_/X sky130_fd_sc_hd__a2bb2o_1
X_4039_ _4039_/A _5980_/B _4039_/C _4039_/D vssd1 vssd1 vccd1 vccd1 _4067_/C sky130_fd_sc_hd__and4_1
XANTENNA__6631__B1 _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7187__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5198__A0 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6147__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5952__A _5952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5370__A0 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__B _6718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5163__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7111__B2 _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6870__B1 _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5425__A1 _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7178__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4936__B1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5338__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6138__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold308 _4757_/X vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 _5259_/X vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_4390_ _4440_/A _4438_/B _4390_/C vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__and3_1
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5073__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _4955_/B _6062_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6061_/A sky130_fd_sc_hd__mux2_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5011_ _5011_/A _5011_/B vssd1 vssd1 vccd1 vccd1 _5012_/B sky130_fd_sc_hd__and2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6962_ _6962_/A _7230_/A vssd1 vssd1 vccd1 vccd1 _6962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6893_ _6893_/A _6893_/B vssd1 vssd1 vccd1 vccd1 _6893_/Y sky130_fd_sc_hd__nor2_1
X_5913_ _5913_/A _5913_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_76_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5844_ _5844_/A vssd1 vssd1 vccd1 vccd1 _5845_/B sky130_fd_sc_hd__inv_2
XANTENNA__5248__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3825__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7514_ _7582_/CLK hold65/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
X_5775_ _5775_/A _5775_/B _5775_/C vssd1 vssd1 vccd1 vccd1 _5777_/C sky130_fd_sc_hd__and3_1
X_4726_ _4825_/B _4748_/A vssd1 vssd1 vccd1 vccd1 _7175_/B sky130_fd_sc_hd__and2b_2
X_7445_ _7446_/CLK _7445_/D vssd1 vssd1 vccd1 vccd1 _7445_/Q sky130_fd_sc_hd__dfxtp_1
X_4657_ _4266_/Y _4652_/Y _4656_/X vssd1 vssd1 vccd1 vccd1 _4658_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5352__A0 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7376_ _7378_/CLK _7376_/D vssd1 vssd1 vccd1 vccd1 _7376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4588_ _3924_/B _4106_/X _4587_/Y _4586_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _4589_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6327_ _4037_/A _6326_/X _3980_/A vssd1 vssd1 vccd1 vccd1 _6332_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4388__A _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6258_ _6258_/A vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__inv_2
X_5209_ hold588/X _5015_/X _5211_/S vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__mux2_1
X_6189_ _3751_/Y _6187_/X _6188_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6189_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5407__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4091__A0 hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold601_A _7529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6907__B2 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5666__B _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5158__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5857__A _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3890_ _6075_/A _4971_/B _6084_/A vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__and3_1
XANTENNA__4909__B1 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5068__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4385__A1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5560_ _5577_/A _5549_/B _5557_/Y _5559_/Y vssd1 vssd1 vccd1 vccd1 _5591_/B sky130_fd_sc_hd__a31oi_4
XFILLER_0_110_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7598_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5491_ _6568_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__or2_4
X_4511_ _4701_/B _4507_/X _4510_/X vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5334__A0 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4442_ _3935_/X _4107_/Y _4441_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _4443_/B sky130_fd_sc_hd__o2bb2a_1
Xhold116 _6193_/X vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 _6422_/Y vssd1 vssd1 vccd1 vccd1 _7580_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7230_ _7230_/A _7230_/B _7230_/C _7230_/D vssd1 vssd1 vccd1 vccd1 _7231_/D sky130_fd_sc_hd__or4_1
Xhold127 _6366_/X vssd1 vssd1 vccd1 vccd1 _6367_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _6006_/X vssd1 vssd1 vccd1 vccd1 _6007_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _7502_/Q vssd1 vssd1 vccd1 vccd1 _6216_/A sky130_fd_sc_hd__buf_2
X_7161_ _7160_/X _4538_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7595_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4373_ _4372_/X _4371_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4374_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5885__B2 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6112_ _6427_/B _6110_/X _6111_/Y _4403_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6112_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7092_/A _7109_/B _7065_/X vssd1 vssd1 vccd1 vccd1 _7092_/X sky130_fd_sc_hd__or3b_1
X_6043_ _6043_/A vssd1 vssd1 vccd1 vccd1 _6043_/Y sky130_fd_sc_hd__inv_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A1 _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4655__B _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4860__A2 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout172_A _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6945_ _6949_/A _6945_/B vssd1 vssd1 vccd1 vccd1 _6945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6876_ _6875_/B _6875_/C _6875_/A vssd1 vssd1 vccd1 vccd1 _6877_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5827_ _5856_/B _5827_/B vssd1 vssd1 vccd1 vccd1 _5829_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5758_ _5758_/A _5758_/B vssd1 vssd1 vccd1 vccd1 _5760_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6117__A2 _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4709_ _7275_/Q _7615_/Q _7607_/Q _7623_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4709_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7428_ _7449_/CLK _7428_/D vssd1 vssd1 vccd1 vccd1 _7428_/Q sky130_fd_sc_hd__dfxtp_1
X_5689_ _5745_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5689_/X sky130_fd_sc_hd__and2_1
XFILLER_0_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4223__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3887__B1 _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7359_ _7427_/CLK _7359_/D vssd1 vssd1 vccd1 vccd1 _7359_/Q sky130_fd_sc_hd__dfxtp_1
Xhold650 _7604_/Q vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _6851_/A vssd1 vssd1 vccd1 vccd1 split20/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4846__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A _4147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5628__B2 _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5628__A1 _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4603__A2 _4601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3811__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6108__A2 _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4214__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output66_A hold94/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5351__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4055__A0 hold558/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4991_ hold553/X _4990_/Y _5039_/S vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5587__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6690__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6730_ _6687_/X _6729_/Y split7/A vssd1 vssd1 vccd1 vccd1 _6742_/B sky130_fd_sc_hd__mux2_4
X_3942_ _4103_/A _6157_/A _6111_/A _6075_/A vssd1 vssd1 vccd1 vccd1 _3943_/D sky130_fd_sc_hd__and4b_1
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3873_ _7421_/Q _7353_/Q _7345_/Q _7325_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3873_/X sky130_fd_sc_hd__mux4_1
X_6661_ _6648_/A _6642_/B _6659_/Y vssd1 vssd1 vccd1 vccd1 _6661_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6592_ _6593_/B _6592_/B vssd1 vssd1 vccd1 vccd1 _6592_/Y sky130_fd_sc_hd__nand2b_1
X_5612_ _6637_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5612_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5543_ _5535_/A split1/X _5539_/X _6518_/A vssd1 vssd1 vccd1 vccd1 _5543_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5474_ _5472_/B _5499_/B _5470_/Y vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__5858__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5753__C _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6211__A _7540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7213_ hold165/X _4385_/X _7227_/S vssd1 vssd1 vccd1 vccd1 _7213_/X sky130_fd_sc_hd__mux2_1
X_4425_ _4672_/B _6107_/B vssd1 vssd1 vccd1 vccd1 _4477_/C sky130_fd_sc_hd__nor2_1
XANTENNA__5858__B2 _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4530__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ _4985_/A _4984_/B vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__or2_1
X_7144_ _7132_/X _7143_/X _7078_/A _6234_/Y vssd1 vssd1 vccd1 vccd1 _7144_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4667_/B _4287_/B vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__and2b_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7074_/A _7074_/B _7043_/S vssd1 vssd1 vccd1 vccd1 _7075_/Y sky130_fd_sc_hd__o21ai_1
X_6026_ _7555_/Q _3698_/A _3728_/A vssd1 vssd1 vccd1 vccd1 _6026_/X sky130_fd_sc_hd__o21a_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6928_ input31/X _4723_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _6928_/X sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_A _7544_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6859_ _6813_/B _6859_/B vssd1 vssd1 vccd1 vccd1 _6860_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout88 _6022_/Y vssd1 vssd1 vccd1 vccd1 _7236_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout77 _6086_/S vssd1 vssd1 vccd1 vccd1 _6168_/S sky130_fd_sc_hd__clkbuf_8
Xfanout99 _6326_/C vssd1 vssd1 vccd1 vccd1 _6329_/A sky130_fd_sc_hd__buf_4
XFILLER_0_107_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold599_A _7259_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5849__A1 _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5849__B2 _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold480 _7364_/Q vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 _7427_/Q vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5171__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4588__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4515__S _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5854__B _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5346__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4760__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _7440_/Q _7432_/Q _7416_/Q _7408_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4210_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4512__A1 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _4973_/X _5189_/X _5194_/S vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5081__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4141_ _3780_/B _6329_/A _4140_/Y _5804_/B _6900_/A vssd1 vssd1 vccd1 vccd1 _4142_/B
+ sky130_fd_sc_hd__a32o_1
X_4072_ _5805_/A hold610/X _6329_/A vssd1 vssd1 vccd1 vccd1 _4072_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4371__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6017__A1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4028__B1 _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4579__A1 _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ _5002_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4974_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6206__A _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3925_ _7283_/Q _7598_/Q _7267_/Q _7491_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3925_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6713_ _6719_/A _6719_/B _6698_/A vssd1 vssd1 vccd1 vccd1 _6714_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6644_ _6553_/Y _6643_/Y split9/A vssd1 vssd1 vccd1 vccd1 _6647_/B sky130_fd_sc_hd__mux2_2
X_3856_ _7422_/Q _7354_/Q _7346_/Q _7326_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3856_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6575_ _6575_/A _6575_/B vssd1 vssd1 vccd1 vccd1 _6576_/B sky130_fd_sc_hd__and2_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3787_ _3779_/X _7230_/C _3787_/C _3787_/D vssd1 vssd1 vccd1 vccd1 _3787_/X sky130_fd_sc_hd__and4bb_1
X_5526_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5527_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5457_ _5456_/Y _5455_/B _5457_/S vssd1 vssd1 vccd1 vccd1 _5459_/B sky130_fd_sc_hd__mux2_2
XANTENNA__4503__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4408_ _4876_/B _4454_/A _4408_/C vssd1 vssd1 vccd1 vccd1 _4408_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5388_ hold460/X _4589_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7481_/D sky130_fd_sc_hd__mux2_1
Xfanout201 _7341_/Q vssd1 vssd1 vccd1 vccd1 _4709_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout212 input44/X vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__clkbuf_8
X_4339_ _4360_/B _4338_/X _4335_/Y vssd1 vssd1 vccd1 vccd1 _6035_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__6087__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7127_ _7118_/X _7120_/X _7126_/X _6326_/C vssd1 vssd1 vccd1 vccd1 _7127_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4197__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7058_ _6872_/A _6922_/B _7051_/Y _7052_/X _7078_/B vssd1 vssd1 vccd1 vccd1 _7058_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__4362__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6009_ _6216_/B _3751_/Y _6190_/S _6216_/C _6007_/A vssd1 vssd1 vccd1 vccd1 _6009_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5939__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6116__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4665__S1 _7341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5955__A _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4417__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4990__A1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5166__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4742__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4245__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3710_ _6326_/B _6421_/B vssd1 vssd1 vccd1 vccd1 _3712_/B sky130_fd_sc_hd__nor2_2
X_4690_ _7379_/Q _7307_/Q _7299_/Q _7291_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4690_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5076__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3641_ _7230_/A vssd1 vssd1 vccd1 vccd1 _6160_/S sky130_fd_sc_hd__inv_2
XANTENNA__4733__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6360_ _7569_/Q hold128/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__mux2_1
X_5311_ hold337/X _4937_/Y _5319_/S vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6696__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6291_ _6872_/A _6290_/C _6290_/B vssd1 vssd1 vccd1 vccd1 _6959_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _4947_/X hold513/X _5248_/S vssd1 vssd1 vccd1 vccd1 _7408_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4592__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5173_ hold229/X _4679_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5750__D _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4124_ _3724_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _4128_/C sky130_fd_sc_hd__and2b_1
Xinput1 custom_settings[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
X_4055_ hold558/X _6844_/A _6023_/S vssd1 vssd1 vccd1 vccd1 _4056_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4957_ _4263_/B _4953_/B _4698_/A vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__o21a_1
X_3908_ _3931_/S _3904_/X _7363_/Q vssd1 vssd1 vccd1 vccd1 _3908_/Y sky130_fd_sc_hd__o21ai_1
X_4888_ hold329/X _4887_/X _5039_/S vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3839_ _7320_/Q _7336_/Q _7312_/Q _7448_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3839_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6627_ _6622_/A split9/X _6627_/C vssd1 vssd1 vccd1 vccd1 _6629_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6558_ _6558_/A _6558_/B vssd1 vssd1 vccd1 vccd1 _6558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5509_ _6518_/A _5509_/B vssd1 vssd1 vccd1 vccd1 _5530_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6489_ _6532_/B vssd1 vssd1 vccd1 vccd1 _6489_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6229__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7230__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold631_A _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4412__A0 _4407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5140__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5860_ _6244_/A _6690_/A _6771_/A _6773_/A vssd1 vssd1 vccd1 vccd1 _5861_/B sky130_fd_sc_hd__and4_1
X_4811_ hold224/X _4434_/Y _4823_/S vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6943__A2 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5791_ _6972_/A _6972_/B vssd1 vssd1 vccd1 vccd1 _7002_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4742_ hold519/X _4589_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7265_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4954__A1 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7530_ _7569_/CLK _7530_/D vssd1 vssd1 vccd1 vccd1 _7530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7461_ _7476_/CLK _7461_/D vssd1 vssd1 vccd1 vccd1 _7461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4673_ _4672_/B _6153_/B vssd1 vssd1 vccd1 vccd1 _4674_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6412_ _6235_/A _6383_/Y _6411_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6412_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7392_ _7396_/CLK _7392_/D vssd1 vssd1 vccd1 vccd1 _7392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3851__A1_N _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6343_ _6220_/C _6333_/X _6342_/Y _6325_/X vssd1 vssd1 vccd1 vccd1 _6343_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6274_ _7109_/A _6275_/B vssd1 vssd1 vccd1 vccd1 _7074_/A sky130_fd_sc_hd__and2_2
X_5225_ hold381/X _4990_/Y _5229_/S vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4565__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ _4996_/X hold586/X _5158_/S vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ hold332/X _4964_/X _5093_/S vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__mux2_1
X_4107_ _4946_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4107_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__6092__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4038_ _6911_/A _7078_/A vssd1 vssd1 vccd1 vccd1 _4039_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7196__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6395__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5989_ _6374_/A _5988_/X _6357_/A _3741_/B _4021_/A vssd1 vssd1 vccd1 vccd1 _5994_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3804__A1_N _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4849__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__C _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5122__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4881__B1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4584__A _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5425__A2 _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5189__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3928__A _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5361__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5354__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 _7320_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5649__C1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4547__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5010_ _5031_/S _5006_/X _5008_/Y _5009_/X vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__a31o_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6074__C1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6961_ _6978_/A _6978_/B _6933_/B _6960_/Y vssd1 vssd1 vccd1 vccd1 _6961_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5912_ hold86/X wire79/X _5911_/X _6218_/A vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__o211a_1
X_6892_ _6840_/A _6840_/B _6890_/Y _6891_/Y _6835_/X vssd1 vssd1 vccd1 vccd1 _6893_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5843_ _5843_/A _5843_/B _5843_/C vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__and3_1
XANTENNA__3838__A _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6214__A _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7513_ _7537_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5774_ _5774_/A _5774_/B vssd1 vssd1 vccd1 vccd1 _5775_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_29_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4725_ _4787_/B _4747_/A vssd1 vssd1 vccd1 vccd1 _7150_/B sky130_fd_sc_hd__and2b_2
XANTENNA__6129__B1 _6128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7444_ _7448_/CLK _7444_/D vssd1 vssd1 vccd1 vccd1 _7444_/Q sky130_fd_sc_hd__dfxtp_1
X_4656_ _4876_/B _4651_/B _4655_/Y _4654_/Y _4953_/A vssd1 vssd1 vccd1 vccd1 _4656_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7375_ _7379_/CLK _7375_/D vssd1 vssd1 vccd1 vccd1 _7375_/Q sky130_fd_sc_hd__dfxtp_1
X_4587_ _6139_/A _4536_/B _6148_/A vssd1 vssd1 vccd1 vccd1 _4587_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4155__A2 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6326_ _7043_/S _6326_/B _6326_/C _6326_/D vssd1 vssd1 vccd1 vccd1 _6326_/X sky130_fd_sc_hd__or4_1
XANTENNA__5104__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ _6872_/A _6875_/A vssd1 vssd1 vccd1 vccd1 _6258_/A sky130_fd_sc_hd__nor2_1
X_5208_ _4973_/X _5207_/X _5212_/S vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__mux2_1
X_6188_ _6188_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6188_/X sky130_fd_sc_hd__or2_1
XANTENNA__4863__B1 _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6095__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5139_ _6911_/A _6225_/B vssd1 vssd1 vccd1 vccd1 _5139_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6065__C1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5812__C1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6368__A0 hold60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4343__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5666__C _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5343__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5174__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4518__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4854__B1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6056__C1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5857__B _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5349__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5031__A0 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5490_ _5459_/B _5489_/Y _5495_/S vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4510_ _5024_/S _4263_/B _6123_/B _4509_/Y _4700_/B vssd1 vssd1 vccd1 vccd1 _4510_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4441_ _6935_/A _4440_/A _4439_/Y _4440_/Y vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__o22a_1
Xhold106 _7581_/Q vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _7524_/Q vssd1 vssd1 vccd1 vccd1 _6185_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ hold245/X _4580_/X _7166_/S vssd1 vssd1 vccd1 vccd1 _7160_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5084__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold128 _7561_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _6212_/X vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4372_ _7427_/Q _7359_/Q _7351_/Q _7331_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4372_/X sky130_fd_sc_hd__mux4_1
X_6111_ _6111_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6111_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _6242_/X _7065_/X _7110_/A vssd1 vssd1 vccd1 vccd1 _7091_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4001__B _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6042_ _4199_/B _6044_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__mux2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A2 _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6047__C1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4073__A1 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout165_A _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6944_ _6989_/A _5789_/Y _6943_/Y _6891_/B _5879_/A vssd1 vssd1 vccd1 vccd1 _6944_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _6875_/A _6875_/B _6875_/C vssd1 vssd1 vccd1 vccd1 _6875_/X sky130_fd_sc_hd__and3_1
X_5826_ _6630_/A _6673_/A _5823_/Y _5856_/A vssd1 vssd1 vccd1 vccd1 _5827_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_106_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5757_ _5757_/A _5757_/B vssd1 vssd1 vccd1 vccd1 _5758_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4708_ _7379_/Q _7307_/Q _7299_/Q _7291_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4708_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5325__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7427_ _7427_/CLK _7427_/D vssd1 vssd1 vccd1 vccd1 _7427_/Q sky130_fd_sc_hd__dfxtp_1
X_5688_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__nor2_1
X_4639_ hold668/X _4638_/C _7606_/Q vssd1 vssd1 vccd1 vccd1 _4639_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3887__A1 _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7358_ _7427_/CLK _7358_/D vssd1 vssd1 vccd1 vccd1 _7358_/Q sky130_fd_sc_hd__dfxtp_1
Xhold651 _7606_/Q vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold640 _7584_/Q vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _7583_/Q vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
X_7289_ _7481_/CLK _7289_/D vssd1 vssd1 vccd1 vccd1 _7289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6309_ _6341_/A _6309_/B vssd1 vssd1 vccd1 vccd1 _6309_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5628__A2 _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4338__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6038__C1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4862__A _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3811__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5169__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5013__B1 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4801__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5316__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4102__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3941__A _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output59_A _7543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4055__A1 _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4990_ _4964_/S _4987_/X _4989_/X vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5079__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3941_ _4084_/A _6057_/A _3941_/C vssd1 vssd1 vccd1 vccd1 _3944_/C sky130_fd_sc_hd__and3_1
X_3872_ _7317_/Q _7333_/Q _7309_/Q _7445_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3872_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6660_ _6670_/A _6648_/X _6658_/X vssd1 vssd1 vccd1 vccd1 _6709_/S sky130_fd_sc_hd__a21o_4
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5611_ _5589_/B _5611_/A2 _5854_/C vssd1 vssd1 vccd1 vccd1 _5614_/B sky130_fd_sc_hd__a21oi_1
X_6591_ _6574_/Y _6613_/B _6592_/B vssd1 vssd1 vccd1 vccd1 _6608_/A sky130_fd_sc_hd__o21ba_1
X_5542_ hold82/A _6808_/B vssd1 vssd1 vccd1 vccd1 _5542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5307__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5473_ hold86/A _6683_/B vssd1 vssd1 vccd1 vccd1 _5499_/B sky130_fd_sc_hd__or2_2
XFILLER_0_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5753__D _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7212_ _7212_/A _7212_/B _7212_/C vssd1 vssd1 vccd1 vccd1 _7227_/S sky130_fd_sc_hd__and3_4
X_4424_ _4672_/B _6107_/B vssd1 vssd1 vccd1 vccd1 _4477_/B sky130_fd_sc_hd__and2_1
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4355_ _4355_/A _4355_/B vssd1 vssd1 vccd1 vccd1 _4984_/B sky130_fd_sc_hd__or2_1
X_7143_ _6989_/A _7140_/Y _7142_/X _7135_/X _7139_/X vssd1 vssd1 vccd1 vccd1 _7143_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ _7074_/A _7074_/B vssd1 vssd1 vccd1 vccd1 _7074_/X sky130_fd_sc_hd__and2_1
X_4286_ _4285_/X _4284_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4287_/B sky130_fd_sc_hd__mux2_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4158__S _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6025_ _6328_/A _6220_/C _6375_/C vssd1 vssd1 vccd1 vccd1 _6025_/Y sky130_fd_sc_hd__a21oi_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4682__A _6166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5497__B _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6991__A0 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6927_ _6927_/A _6927_/B _6925_/X vssd1 vssd1 vccd1 vccd1 _6927_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6858_ _6858_/A vssd1 vssd1 vccd1 vccd1 _7030_/A sky130_fd_sc_hd__inv_2
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 _4290_/X vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__buf_4
Xfanout78 _4612_/B vssd1 vssd1 vccd1 vccd1 _5031_/S sky130_fd_sc_hd__clkbuf_8
X_5809_ _5810_/A _5810_/B _5810_/C _5810_/D vssd1 vssd1 vccd1 vccd1 wire79/A sky130_fd_sc_hd__nor4_1
XFILLER_0_91_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6789_ _6789_/A _6789_/B vssd1 vssd1 vccd1 vccd1 _6789_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5018__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 _5143_/X vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold470 _4759_/X vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold492 _5283_/X vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold661_A _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3761__A _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7223__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5234__A0 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3891__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4531__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5854__C _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5362__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _6326_/B _4140_/B vssd1 vssd1 vccd1 vccd1 _4140_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__3671__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ hold99/A hold66/X _7249_/S vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__mux2_1
XANTENNA__4371__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7214__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5598__A _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6193__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4028__A1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4973_ _4083_/X _4972_/X _4970_/X _5022_/A vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__a211o_4
XANTENNA__4579__A2 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3924_ _6157_/A _3924_/B vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__nand2_1
X_6712_ _6756_/A _6675_/X _6751_/B _6711_/Y vssd1 vssd1 vccd1 vccd1 split7/A sky130_fd_sc_hd__a31o_4
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6643_ _6643_/A _6643_/B vssd1 vssd1 vccd1 vccd1 _6643_/Y sky130_fd_sc_hd__xnor2_1
X_3855_ _7318_/Q _7334_/Q _7310_/Q _7446_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3855_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6574_ _6613_/A vssd1 vssd1 vccd1 vccd1 _6574_/Y sky130_fd_sc_hd__inv_2
X_3786_ _3780_/B _7123_/C _3785_/X vssd1 vssd1 vccd1 vccd1 _3787_/C sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout128_A _7587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7434_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5525_ _5525_/A vssd1 vssd1 vccd1 vccd1 _5525_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5456_ _5456_/A _5456_/B vssd1 vssd1 vccd1 vccd1 _5456_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4407_ _4407_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4408_/C sky130_fd_sc_hd__nand2_1
X_5387_ hold459/X _4629_/X _5391_/S vssd1 vssd1 vccd1 vccd1 _5387_/X sky130_fd_sc_hd__mux2_1
Xfanout202 _4369_/S0 vssd1 vssd1 vccd1 vccd1 _4371_/S0 sky130_fd_sc_hd__buf_8
XANTENNA__5272__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4677__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 input44/X vssd1 vssd1 vccd1 vccd1 _6218_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4337_/X _4336_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4338_/X sky130_fd_sc_hd__mux2_1
X_7126_ _7023_/A _7122_/X _7125_/X vssd1 vssd1 vccd1 vccd1 _7126_/X sky130_fd_sc_hd__a21o_1
X_4269_ _4269_/A _4879_/S vssd1 vssd1 vccd1 vccd1 _4701_/B sky130_fd_sc_hd__or2_2
X_7057_ _6244_/A _6911_/A _7098_/A _7056_/X vssd1 vssd1 vccd1 vccd1 _7078_/B sky130_fd_sc_hd__o211a_1
X_6008_ _6216_/B _6008_/B vssd1 vssd1 vccd1 vccd1 _6190_/S sky130_fd_sc_hd__nand2_4
XANTENNA__7199__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4362__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7205__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4616__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3873__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3756__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7141__B1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5182__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3864__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4430__A1 _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4718__C1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3640_ _5988_/A vssd1 vssd1 vccd1 vccd1 _6223_/A sky130_fd_sc_hd__inv_6
X_5310_ hold239/X _4897_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5881__A _5952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6290_ _6872_/A _6290_/B _6290_/C vssd1 vssd1 vccd1 vccd1 _6290_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ hold512/X _4964_/X _5247_/S vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5092__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4592__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5172_ hold477/X _4589_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7377_/D sky130_fd_sc_hd__mux2_1
X_4123_ _4123_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4905_/B sky130_fd_sc_hd__nand2_2
X_4054_ _4053_/X hold60/X _7241_/S vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
Xinput2 custom_settings[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4436__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3855__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ _4955_/B _4951_/A _6096_/A vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3907_ _3905_/X _3906_/X _3931_/S vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__mux2_1
X_4887_ _4872_/Y _4886_/X _4964_/S vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__mux2_8
X_3838_ _3886_/S _3838_/B vssd1 vssd1 vccd1 vccd1 _3838_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6626_ _6628_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _6627_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6557_ _6557_/A _6557_/B _6557_/C vssd1 vssd1 vccd1 vccd1 _6558_/B sky130_fd_sc_hd__nor3_1
X_5508_ _5507_/A _5507_/B _6518_/A vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__a21o_1
X_3769_ _6235_/A _7123_/A _7025_/A _6244_/A vssd1 vssd1 vccd1 vccd1 _3770_/B sky130_fd_sc_hd__or4_1
XFILLER_0_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6488_ _6481_/S _6486_/X _6487_/X vssd1 vssd1 vccd1 vccd1 _6532_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5439_ _5438_/A _5438_/B _5438_/C _7497_/Q vssd1 vssd1 vccd1 vccd1 _5444_/C sky130_fd_sc_hd__o31ai_2
XFILLER_0_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7109_ _7109_/A _7109_/B _7109_/C vssd1 vssd1 vccd1 vccd1 _7109_/X sky130_fd_sc_hd__and3_1
XFILLER_0_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3846__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6165__A1 _3702_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6165__B2 _6022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7114__B1 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3933__B _6166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4256__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ hold217/X _4111_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7292_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3837__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5790_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _6972_/B sky130_fd_sc_hd__xnor2_1
X_4741_ hold518/X _4629_/X _4745_/S vssd1 vssd1 vccd1 vccd1 _4741_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5087__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7460_ _7596_/CLK _7460_/D vssd1 vssd1 vccd1 vccd1 _7460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4672_ _6153_/B _4672_/B vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__6156__A1 _3702_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6156__B2 _6022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6411_ hold130/X _6415_/A _6356_/B hold254/X vssd1 vssd1 vccd1 vccd1 _6411_/X sky130_fd_sc_hd__a22o_1
X_7391_ _7400_/CLK _7391_/D vssd1 vssd1 vccd1 vccd1 _7391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6342_ _6234_/Y _6341_/Y _6333_/A _6236_/A vssd1 vssd1 vccd1 vccd1 _6342_/Y sky130_fd_sc_hd__o211ai_1
X_6273_ _6273_/A _6851_/A vssd1 vssd1 vccd1 vccd1 _6275_/B sky130_fd_sc_hd__or2_1
X_5224_ hold483/X _4947_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _7400_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4020__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5155_ hold585/X _5015_/X _5157_/S vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4890__A1 _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _7343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6616__C1 _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5086_ _5085_/X _4921_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _7335_/D sky130_fd_sc_hd__mux2_1
X_4106_ _4946_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__and2_2
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4037_ _4037_/A _5805_/A vssd1 vssd1 vccd1 vccd1 _4037_/X sky130_fd_sc_hd__or2_4
XFILLER_0_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3828__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6395__B2 hold92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5988_ _5988_/A _5988_/B _5811_/B vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__or3b_1
X_4939_ _4938_/X _4921_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _7311_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6147__A1 _3702_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6147__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6609_ _6565_/Y _6608_/Y split9/A vssd1 vssd1 vccd1 vccd1 _6612_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7589_ _7590_/CLK _7589_/D vssd1 vssd1 vccd1 vccd1 _7589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4881__A1 _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5696__A _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4804__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6138__A1 _3702_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6138__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4244__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5649__B1 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4547__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5370__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7151__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6960_ _6989_/A _6960_/B vssd1 vssd1 vccd1 vccd1 _6960_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5911_ _6962_/A _5811_/Y _5910_/X _5811_/A _5810_/X vssd1 vssd1 vccd1 vccd1 _5911_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ _6891_/A _6891_/B vssd1 vssd1 vccd1 vccd1 _6891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ _5843_/A _5843_/B _5843_/C vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4927__A2 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5773_ _6874_/A _6871_/A _6869_/A _6261_/A vssd1 vssd1 vccd1 vccd1 _5774_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7512_ _7582_/CLK hold73/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
X_4724_ _4723_/Y hold599/X _4724_/S vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6129__B2 _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7443_ _7443_/CLK _7443_/D vssd1 vssd1 vccd1 vccd1 _7443_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3854__A _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4655_ _4698_/B _4698_/C vssd1 vssd1 vccd1 vccd1 _4655_/Y sky130_fd_sc_hd__nand2_1
X_7374_ _7618_/CLK _7374_/D vssd1 vssd1 vccd1 vccd1 _7374_/Q sky130_fd_sc_hd__dfxtp_1
X_4586_ _6628_/A _4440_/A _4440_/Y _4585_/Y vssd1 vssd1 vccd1 vccd1 _4586_/X sky130_fd_sc_hd__o22a_1
XANTENNA_fanout110_A _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6230__A _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4560__B1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6325_ _6233_/Y _6313_/X _7122_/A _6315_/X _6326_/C vssd1 vssd1 vccd1 vccd1 _6325_/X
+ sky130_fd_sc_hd__o311a_1
X_6256_ _6872_/A _6875_/A vssd1 vssd1 vccd1 vccd1 _6974_/B sky130_fd_sc_hd__nand2_2
X_5207_ hold415/X _4990_/Y _5211_/S vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5280__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4685__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4863__A1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6187_ hold62/X hold40/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6187_/X sky130_fd_sc_hd__mux2_1
X_5138_ _7244_/A _7244_/B vssd1 vssd1 vccd1 vccd1 _7362_/D sky130_fd_sc_hd__or2_1
XFILLER_0_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5069_ hold252/X _4964_/X _5075_/S vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7014__C1 _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__B1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5040__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4000__C1 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5190__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4595__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4465__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5365__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _4440_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4440_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 _6423_/Y vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3674__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 _6360_/X vssd1 vssd1 vccd1 vccd1 _6361_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _6185_/X vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4371_ _7323_/Q _7339_/Q _7315_/Q _7451_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4371_/X sky130_fd_sc_hd__mux4_1
X_6110_ _6328_/A _4403_/Y _6109_/X _6375_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6110_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6819__C1 _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5098__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7090_/A _7090_/B vssd1 vssd1 vccd1 vccd1 _7090_/X sky130_fd_sc_hd__or2_1
XANTENNA__4001__C _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6041_ _6040_/X hold50/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__mux2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7621_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__B _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5270__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6943_ _6261_/A _6875_/A _5787_/Y vssd1 vssd1 vccd1 vccd1 _6943_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6874_ _6874_/A _6888_/A _6874_/C vssd1 vssd1 vccd1 vccd1 _6875_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5558__C1 _5556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5825_ _5856_/A _5918_/D _6683_/A _5825_/D vssd1 vssd1 vccd1 vccd1 _5856_/B sky130_fd_sc_hd__and4b_1
XANTENNA__4455__A2_N _4460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5756_ _5768_/A _5768_/B vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__nand2_1
X_4707_ _4705_/X _4706_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5275__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5783__B _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5687_ _5683_/X _5684_/Y _5654_/A _5740_/A vssd1 vssd1 vccd1 vccd1 _5688_/B sky130_fd_sc_hd__o211a_1
X_7426_ _7427_/CLK _7426_/D vssd1 vssd1 vccd1 vccd1 _7426_/Q sky130_fd_sc_hd__dfxtp_1
X_4638_ _7605_/Q _7606_/Q _4638_/C vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__or3_1
XANTENNA__7056__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold630 _5108_/X vssd1 vssd1 vccd1 vccd1 _7349_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4569_ _4667_/B _4564_/X _4568_/X vssd1 vssd1 vccd1 vccd1 _6135_/B sky130_fd_sc_hd__a21oi_2
X_7357_ _7424_/CLK _7357_/D vssd1 vssd1 vccd1 vccd1 _7357_/Q sky130_fd_sc_hd__dfxtp_1
Xhold652 _7190_/X vssd1 vssd1 vccd1 vccd1 _7606_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold641 _6844_/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold663 _7587_/Q vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5089__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7288_ _7487_/CLK _7288_/D vssd1 vssd1 vccd1 vccd1 _7288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6308_ _7109_/A _7109_/C _7109_/B vssd1 vssd1 vccd1 vccd1 _6309_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4619__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6239_ _7123_/A _6754_/A vssd1 vssd1 vccd1 vccd1 _6276_/B sky130_fd_sc_hd__or2_2
XANTENNA__5304__A _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4846__C _4846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4862__B _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5261__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6135__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5974__A _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5185__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4529__S _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3941__B _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4686__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5252__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ _4862_/A _6039_/A _6066_/A _6048_/A vssd1 vssd1 vccd1 vccd1 _3941_/C sky130_fd_sc_hd__and4b_1
XANTENNA__4264__S _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3669__A _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3871_ _7363_/Q _3871_/B vssd1 vssd1 vccd1 vccd1 _3871_/X sky130_fd_sc_hd__and2_1
XANTENNA__5004__A1 _4238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5610_ _5604_/A _5660_/B _5603_/X _5609_/B vssd1 vssd1 vccd1 vccd1 _6451_/B sky130_fd_sc_hd__a31o_1
X_6590_ _6618_/B _6619_/A _6579_/Y vssd1 vssd1 vccd1 vccd1 _6613_/B sky130_fd_sc_hd__a21oi_4
X_5541_ _7494_/Q _5541_/A2 _5538_/X _6875_/A vssd1 vssd1 vccd1 vccd1 _5541_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_14_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7211_ _5393_/A _7211_/B _7211_/C vssd1 vssd1 vccd1 vccd1 _7228_/S sky130_fd_sc_hd__and3b_4
X_5472_ _5470_/Y _5472_/B vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4515__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4423_ _4667_/B _4418_/X _4422_/X vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4354_ _4321_/X _4933_/A _4353_/A vssd1 vssd1 vccd1 vccd1 _4355_/B sky130_fd_sc_hd__o21a_1
X_7142_ _6282_/A _6341_/Y _7141_/Y vssd1 vssd1 vccd1 vccd1 _7142_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7073_ _7073_/A _7073_/B vssd1 vssd1 vccd1 vccd1 _7073_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4818__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4285_ _7268_/Q _7608_/Q _7600_/Q _7616_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4285_/X sky130_fd_sc_hd__mux4_1
X_6024_ _6096_/A _4861_/B _4953_/B vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__o21a_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5243__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6926_ _6927_/A _6927_/B _6925_/X vssd1 vssd1 vccd1 vccd1 _6926_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6991__A1 _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6857_ _6857_/A _7029_/A vssd1 vssd1 vccd1 vccd1 _6858_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5808_ _5808_/A _6329_/B vssd1 vssd1 vccd1 vccd1 _5810_/D sky130_fd_sc_hd__nor2_1
X_6788_ _6793_/A _6793_/B vssd1 vssd1 vccd1 vccd1 _6817_/B sky130_fd_sc_hd__and2_1
XFILLER_0_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5739_ _5739_/A _5739_/B vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7409_ _7441_/CLK _7409_/D vssd1 vssd1 vccd1 vccd1 _7409_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4506__B1 _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold471 _7256_/Q vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 _5387_/X vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A _4290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 _7400_/Q vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _7305_/Q vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4962__A2_N _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4809__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5034__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4873__A _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4668__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6982__A1 _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3891__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4812__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3936__B _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5854__D _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4113__A _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output71_A _7520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3720__A1 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4846_/A input13/X _4021_/B hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__o22a_1
XFILLER_0_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5879__A _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6422__B1 _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _4972_/A _4972_/B vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__or2_1
XANTENNA__6973__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6973__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3923_ _6148_/A _6139_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _3924_/B sky130_fd_sc_hd__and3_1
XFILLER_0_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6711_ _6663_/X _6668_/X _6706_/X _6709_/X _6756_/B vssd1 vssd1 vccd1 vccd1 _6711_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_0_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3854_ _3886_/S _3854_/B vssd1 vssd1 vccd1 vccd1 _3854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6642_ _6648_/A _6642_/B vssd1 vssd1 vccd1 vccd1 _6642_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6503__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6186__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6573_ _6637_/A _6573_/B vssd1 vssd1 vccd1 vccd1 _6613_/A sky130_fd_sc_hd__xnor2_1
X_3785_ _7543_/Q _3712_/B _3716_/B _7557_/Q vssd1 vssd1 vccd1 vccd1 _3785_/X sky130_fd_sc_hd__a22o_1
X_5524_ _6568_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5525_/A sky130_fd_sc_hd__or2_4
XFILLER_0_41_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4023__A _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5455_ _6871_/A _5455_/B vssd1 vssd1 vccd1 vccd1 _5456_/B sky130_fd_sc_hd__xnor2_1
X_4406_ _4260_/X _4407_/B _4405_/X vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7579_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5386_ _5385_/X _4538_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7480_/D sky130_fd_sc_hd__mux2_1
Xfanout203 _7340_/Q vssd1 vssd1 vccd1 vccd1 _4369_/S0 sky130_fd_sc_hd__buf_8
XANTENNA__4677__B _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7125_ _6301_/A _6911_/A _7098_/A _7124_/X vssd1 vssd1 vccd1 vccd1 _7125_/X sky130_fd_sc_hd__a31o_1
X_4337_ _7421_/Q _7353_/Q _7345_/Q _7325_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4337_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6110__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4268_ _5974_/C _3989_/X _4131_/X _4267_/X vssd1 vssd1 vccd1 vccd1 _4879_/S sky130_fd_sc_hd__a31o_2
X_7056_ _7123_/A _7230_/A vssd1 vssd1 vccd1 vccd1 _7056_/X sky130_fd_sc_hd__or2_1
X_6007_ _6007_/A _6007_/B vssd1 vssd1 vccd1 vccd1 _6007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4199_ _4873_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4209_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5216__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6413__A0 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6964__A1 _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _7557_/Q _6909_/B vssd1 vssd1 vccd1 vccd1 _6910_/C sky130_fd_sc_hd__or2_1
XANTENNA__3873__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6177__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3756__B _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3950__B2 _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5152__A0 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7244__A _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3702__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 _7618_/Q vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4663__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6955__A1 _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3864__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4430__A2 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7132__A1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5240_ _4921_/X _5239_/X _5248_/S vssd1 vssd1 vccd1 vccd1 _7407_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5373__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ hold476/X _4629_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__mux2_1
X_4122_ _6922_/A _6920_/A _4122_/C _4122_/D vssd1 vssd1 vccd1 vccd1 _4123_/B sky130_fd_sc_hd__or4_4
X_4053_ _4846_/A input9/X _4021_/B hold110/X vssd1 vssd1 vccd1 vccd1 _4053_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 custom_settings[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7199__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4955_ _4955_/A _4955_/B vssd1 vssd1 vccd1 vccd1 _4955_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4957__B1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3855__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3906_ _7270_/Q _7610_/Q _7602_/Q _7618_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3906_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4886_ _4963_/S _4883_/X _4885_/X vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout140_A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3837_ _7400_/Q _7392_/Q _7368_/Q _7384_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3838_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6625_ _6742_/A _6625_/B vssd1 vssd1 vccd1 vccd1 _6694_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6556_ _6754_/A _6556_/B vssd1 vssd1 vccd1 vccd1 _6597_/B sky130_fd_sc_hd__or2_1
X_3768_ _6962_/A _6935_/A _6872_/A _6311_/A vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__or4_1
XANTENNA__3932__A1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5507_ _5507_/A _5507_/B vssd1 vssd1 vccd1 vccd1 _5509_/B sky130_fd_sc_hd__and2_1
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5283__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6487_ _6521_/A _6487_/B _6509_/B vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__and3_1
X_3699_ _7555_/Q _7554_/Q _6225_/A vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__or3_4
X_5438_ _5438_/A _5438_/B _5438_/C _5437_/Y vssd1 vssd1 vccd1 vccd1 _5444_/B sky130_fd_sc_hd__or4b_1
X_5369_ hold189/X _4629_/X _5373_/S vssd1 vssd1 vccd1 vccd1 _5369_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7108_ _7109_/B _7108_/B vssd1 vssd1 vccd1 vccd1 _7108_/Y sky130_fd_sc_hd__xnor2_1
X_7039_ _7040_/B _7039_/B vssd1 vssd1 vccd1 vccd1 _7039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6937__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3846__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3767__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5193__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6928__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5368__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3837__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5600__A1 _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ _4739_/X _4538_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7264_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6053__A _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4671_ _4667_/B _4670_/X _4667_/Y vssd1 vssd1 vccd1 vccd1 _6153_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5364__A0 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7390_ _7400_/CLK _7390_/D vssd1 vssd1 vccd1 vccd1 _7390_/Q sky130_fd_sc_hd__dfxtp_1
X_6410_ _6409_/X hold641/X _6414_/S vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6341_ _6341_/A _7101_/B vssd1 vssd1 vccd1 vccd1 _6341_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6199__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6272_ _7025_/A _6882_/A vssd1 vssd1 vccd1 vccd1 _6339_/A sky130_fd_sc_hd__nor2_1
X_5223_ hold482/X _4964_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4020__B _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5154_ _4973_/X _5153_/X _5158_/S vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4105_ _4119_/A _4279_/C vssd1 vssd1 vccd1 vccd1 _4942_/B sky130_fd_sc_hd__nand2_4
XANTENNA__4955__B _4955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5085_ hold298/X _4937_/Y _5093_/S vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6092__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6228__A _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6092__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4036_ _4036_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_79_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4971__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3850__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3828__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5278__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _6417_/B _3988_/C _4139_/B vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__o21a_1
X_4938_ hold576/X _4937_/Y _5039_/S vssd1 vssd1 vccd1 vccd1 _4938_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4869_ _6874_/A _4868_/Y _4945_/B vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6608_ _6608_/A _6608_/B vssd1 vssd1 vccd1 vccd1 _6608_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7588_ _7590_/CLK _7588_/D vssd1 vssd1 vccd1 vccd1 _7588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6539_ _6538_/Y _6509_/B _6434_/B _6481_/S vssd1 vssd1 vccd1 vccd1 _6540_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5026__B _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4330__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5977__A _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5696__B _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5188__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5346__A0 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4820__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4244__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7151__B _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6074__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6074__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4085__B1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5910_ _5933_/B _5909_/Y _5970_/A _5495_/S vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6890_ _6780_/X _6821_/X _6828_/Y _6888_/Y vssd1 vssd1 vccd1 vccd1 _6890_/Y sky130_fd_sc_hd__a31oi_1
X_5841_ _5841_/A _5841_/B vssd1 vssd1 vccd1 vccd1 _5843_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5772_ _6690_/A _6802_/B _5788_/D _6802_/A vssd1 vssd1 vccd1 vccd1 _5775_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7511_ _7581_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4723_ _4723_/A _6015_/C vssd1 vssd1 vccd1 vccd1 _4723_/Y sky130_fd_sc_hd__nor2_1
X_7442_ _7443_/CLK _7442_/D vssd1 vssd1 vccd1 vccd1 _7442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6129__A2 _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ _4654_/A vssd1 vssd1 vccd1 vccd1 _4654_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7373_ _7476_/CLK _7373_/D vssd1 vssd1 vccd1 vccd1 _7373_/Q sky130_fd_sc_hd__dfxtp_1
X_4585_ _4633_/B _4585_/B vssd1 vssd1 vccd1 vccd1 _4585_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4560__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6324_ _7137_/A _7121_/B vssd1 vssd1 vccd1 vccd1 _7122_/A sky130_fd_sc_hd__and2_1
XANTENNA__4031__A _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6255_ _6264_/A _6319_/A vssd1 vssd1 vccd1 vccd1 _6974_/A sky130_fd_sc_hd__or2_2
XFILLER_0_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5206_ _4947_/X hold362/X _5212_/S vssd1 vssd1 vccd1 vccd1 _7392_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6186_ _3751_/Y _6184_/X hold118/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6186_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4177__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5137_ _4036_/A input33/X _6229_/S vssd1 vssd1 vccd1 vccd1 _7244_/B sky130_fd_sc_hd__mux2_1
X_5068_ _5067_/X _4921_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _7327_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6065__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6065__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4076__B1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4019_ _6417_/B _7244_/A vssd1 vssd1 vccd1 vccd1 _4039_/C sky130_fd_sc_hd__nor2_4
XANTENNA__5812__B2 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5812__A1 _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7014__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold315_A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5328__A0 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6421__A _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4876__A _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4087__S _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6056__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6056__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5803__A1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4815__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4465__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3955__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold108 _6425_/Y vssd1 vssd1 vccd1 vccd1 _7581_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _4368_/X _4369_/X _7342_/Q vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold119 _6186_/X vssd1 vssd1 vccd1 vccd1 _7524_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5381__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3690__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6922_/A _6038_/X _6039_/Y _4902_/A _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6040_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6047__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6047__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4058__B1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ _4084_/A _6949_/A _6940_/Y _6941_/X _3949_/Y vssd1 vssd1 vccd1 vccd1 _6942_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6873_ _6888_/A _6874_/C _6872_/X _5787_/Y vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__a22o_1
X_5824_ _6690_/A _6802_/A _6771_/A _6773_/A vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__and4_1
XANTENNA__4026__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _5766_/B _5755_/B vssd1 vssd1 vccd1 vccd1 _5768_/B sky130_fd_sc_hd__nor2_1
X_4706_ _7483_/Q _7471_/Q _7463_/Q _7257_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4706_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4781__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6241__A _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5686_ _6581_/A _6802_/B _5652_/B _5651_/A vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__a31o_1
X_7425_ _7450_/CLK _7425_/D vssd1 vssd1 vccd1 vccd1 _7425_/Q sky130_fd_sc_hd__dfxtp_1
X_4637_ _4685_/A _4637_/B vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__or2_4
XANTENNA__7056__B _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 _7605_/Q vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4568_ _4667_/B _4568_/B vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__and2b_1
X_7356_ _7423_/CLK _7356_/D vssd1 vssd1 vccd1 vccd1 _7356_/Q sky130_fd_sc_hd__dfxtp_1
Xhold631 _6864_/A vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 _6410_/X vssd1 vssd1 vccd1 vccd1 _7578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _7557_/Q vssd1 vssd1 vccd1 vccd1 _6301_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4499_ _4689_/A _4499_/B vssd1 vssd1 vccd1 vccd1 _4499_/X sky130_fd_sc_hd__and2_1
X_7287_ _7379_/CLK _7287_/D vssd1 vssd1 vccd1 vccd1 _7287_/Q sky130_fd_sc_hd__dfxtp_1
X_6307_ _6339_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _7109_/C sky130_fd_sc_hd__or2_1
Xhold664 _7552_/Q vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
X_6238_ _7123_/A _6754_/A vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__and2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ hold74/X hold54/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6169_/X sky130_fd_sc_hd__mux2_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6038__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6038__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7011__S _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4772__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4370__S _7342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5990__A _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6029__B2 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6029__A1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6326__A _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4686__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _3868_/X _3869_/X _3915_/A vssd1 vssd1 vccd1 vccd1 _3871_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4763__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5540_ _7494_/Q split1/X _5538_/X vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5471_ _6518_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5472_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4422_ _4667_/B _4422_/B vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__and2b_1
X_7210_ _7209_/X _4685_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7615_/D sky130_fd_sc_hd__mux2_1
X_4353_ _4353_/A _4353_/B vssd1 vssd1 vccd1 vccd1 _4933_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7141_ _6282_/A _6341_/Y _7043_/S vssd1 vssd1 vccd1 vccd1 _7141_/Y sky130_fd_sc_hd__o21ai_1
X_4284_ _7372_/Q _7300_/Q _7292_/Q _7284_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4284_/X sky130_fd_sc_hd__mux4_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7072_ _7072_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7072_/Y sky130_fd_sc_hd__nand2_1
X_6023_ _3663_/Y _4861_/B _6023_/S vssd1 vssd1 vccd1 vccd1 _6023_/X sky130_fd_sc_hd__mux2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6925_ _6925_/A _6925_/B _6925_/C _6925_/D vssd1 vssd1 vccd1 vccd1 _6925_/X sky130_fd_sc_hd__and4_1
XFILLER_0_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6856_ _6857_/A _7029_/A vssd1 vssd1 vccd1 vccd1 _6856_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5807_ _6900_/A _4119_/A _4128_/A vssd1 vssd1 vccd1 vccd1 _6329_/B sky130_fd_sc_hd__a21o_1
X_3999_ _4001_/D _7473_/Q _5985_/B _4124_/B _5810_/A vssd1 vssd1 vccd1 vccd1 _3999_/X
+ sky130_fd_sc_hd__o221a_1
X_6787_ _6726_/Y _6786_/Y _6790_/S vssd1 vssd1 vccd1 vccd1 _6793_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4754__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5738_ _5757_/A _5757_/B vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4506__A1 _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5669_ _5671_/D vssd1 vssd1 vccd1 vccd1 _5669_/Y sky130_fd_sc_hd__inv_2
X_7408_ _7439_/CLK _7408_/D vssd1 vssd1 vccd1 vccd1 _7408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold450 _5381_/X vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _7463_/Q vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
X_7339_ _7434_/CLK _7339_/D vssd1 vssd1 vccd1 vccd1 _7339_/Q sky130_fd_sc_hd__dfxtp_1
Xhold472 _7286_/Q vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _5223_/X vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _4839_/X vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5034__B _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4873__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold647_A _7556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4668__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6982__A2 _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4745__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3953__C1 _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5170__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output64_A _7580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__A0 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4971_ _6075_/A _4971_/B vssd1 vssd1 vccd1 vccd1 _4972_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3922_ _6139_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6710_ _6710_/A _6710_/B vssd1 vssd1 vccd1 vccd1 _6756_/B sky130_fd_sc_hd__or2_4
X_3853_ _7398_/Q _7390_/Q _7366_/Q _7382_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3854_/B sky130_fd_sc_hd__mux4_1
X_6641_ _6666_/A _6670_/A _6670_/B _6616_/X _6617_/A vssd1 vssd1 vccd1 vccd1 _6642_/B
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4736__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6572_ _6869_/A _6573_/B vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__and2_1
X_3784_ _5811_/B _6415_/A vssd1 vssd1 vccd1 vccd1 _7230_/C sky130_fd_sc_hd__or2_2
XFILLER_0_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5523_ _6568_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7135__C1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5454_ _5454_/A _5454_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _5457_/S sky130_fd_sc_hd__nand3_4
X_5385_ hold427/X _4580_/X _5391_/S vssd1 vssd1 vccd1 vccd1 _5385_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5161__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4405_ _4999_/B _4454_/A vssd1 vssd1 vccd1 vccd1 _4405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout204 _4709_/S0 vssd1 vssd1 vccd1 vccd1 _4706_/S0 sky130_fd_sc_hd__buf_8
X_4336_ _7317_/Q _7333_/Q _7309_/Q _7445_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4336_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5135__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7124_ _6962_/A _6922_/B _7123_/X vssd1 vssd1 vccd1 vccd1 _7124_/X sky130_fd_sc_hd__a21o_1
X_4267_ _5974_/C _4267_/B _4267_/C _4267_/D vssd1 vssd1 vccd1 vccd1 _4267_/X sky130_fd_sc_hd__and4b_1
X_7055_ _6247_/B _7074_/A _7023_/C _6913_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _7055_/X
+ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4198_ _4199_/B vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__inv_2
X_6006_ _5132_/B _6005_/X _6216_/C vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4913__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4975__B2 _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6908_ _6872_/A _6911_/A _7098_/A _6907_/X vssd1 vssd1 vccd1 vccd1 _6908_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6839_ _6779_/Y _6838_/Y _6891_/B vssd1 vssd1 vccd1 vccd1 _6840_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3950__A2 _3705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold280 _7294_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _7217_/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6404__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4966__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4823__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4718__A1 _4144_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5391__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3963__A _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5143__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ _5169_/X _4538_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7376_/D sky130_fd_sc_hd__mux2_1
X_4121_ _4267_/C _4121_/B _4134_/D vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__nand3_2
X_4052_ _5805_/A _4051_/X _6329_/A vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__mux2_1
Xinput4 custom_settings[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
XANTENNA__4733__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4501__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4954_ _6793_/A _4123_/B _4219_/B _4953_/Y _4123_/A vssd1 vssd1 vccd1 vccd1 _4954_/X
+ sky130_fd_sc_hd__o221a_1
X_3905_ _7374_/Q _7302_/Q _7294_/Q _7286_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3905_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4885_ _6039_/A _4986_/S _4349_/Y _4884_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4885_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6233__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3836_ _7440_/Q _7432_/Q _7416_/Q _7408_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3836_/X sky130_fd_sc_hd__mux4_1
X_6624_ _6871_/A _6625_/B vssd1 vssd1 vccd1 vccd1 _6624_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4034__A _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5382__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6555_ _6597_/A vssd1 vssd1 vccd1 vccd1 _6555_/Y sky130_fd_sc_hd__inv_2
X_3767_ _7230_/A _4036_/A vssd1 vssd1 vccd1 vccd1 _7123_/C sky130_fd_sc_hd__and2_2
X_5506_ _5499_/B _5481_/Y _5500_/B split8/X vssd1 vssd1 vccd1 vccd1 _5507_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3698_ _3698_/A _3992_/C vssd1 vssd1 vccd1 vccd1 _5985_/A sky130_fd_sc_hd__nor2_4
XANTENNA__5134__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6486_ _6486_/A _6486_/B vssd1 vssd1 vccd1 vccd1 _6486_/X sky130_fd_sc_hd__or2_1
X_5437_ _5437_/A _5437_/B vssd1 vssd1 vccd1 vccd1 _5437_/Y sky130_fd_sc_hd__nand2_1
X_5368_ _4538_/X _5367_/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7468_/D sky130_fd_sc_hd__mux2_1
X_5299_ hold196/X _5015_/X _5301_/S vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__mux2_1
X_4319_ _4360_/B _4314_/X _4318_/X vssd1 vssd1 vccd1 vccd1 _6053_/B sky130_fd_sc_hd__a21oi_2
X_7107_ _6084_/A _5804_/C _7105_/Y _7106_/X _6326_/C vssd1 vssd1 vccd1 vccd1 _7107_/X
+ sky130_fd_sc_hd__a221o_1
X_7038_ _7040_/B _7039_/B vssd1 vssd1 vccd1 vccd1 _7038_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4643__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__A _6427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5373__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3783__A hold97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5125__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4818__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4884__B1 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__A _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6389__A0 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4939__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7050__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6928__A2 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5600__A2 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4670_ _4669_/X _4668_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4670_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4789__A _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5384__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3693__A _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6340_ _7109_/A _7100_/C _7109_/B vssd1 vssd1 vccd1 vccd1 _7101_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5116__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6271_ _7137_/A _7137_/B _6233_/Y vssd1 vssd1 vccd1 vccd1 _6271_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6313__B1 _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5222_ _5221_/X _4921_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _7399_/D sky130_fd_sc_hd__mux2_1
X_5153_ hold346/X _4990_/Y _5157_/S vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__mux2_1
X_4104_ _4103_/A _5019_/A _4440_/A vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6616__A1 _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5084_ _5083_/X _4897_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _7334_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4627__B1 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4035_ _4035_/A _6383_/B vssd1 vssd1 vccd1 vccd1 _6023_/S sky130_fd_sc_hd__nand2_4
XANTENNA__4029__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3850__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6244__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _3980_/A _4125_/X _5985_/Y _4011_/X vssd1 vssd1 vccd1 vccd1 _5994_/C sky130_fd_sc_hd__a31o_1
X_4937_ _4948_/B _4936_/Y _4935_/X vssd1 vssd1 vccd1 vccd1 _4937_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_47_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4868_ _4942_/B _4868_/B vssd1 vssd1 vccd1 vccd1 _4868_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5355__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ _3915_/A _3815_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _3819_/Y sky130_fd_sc_hd__a21oi_1
X_6607_ _6608_/A _6608_/B vssd1 vssd1 vccd1 vccd1 _6607_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5294__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4799_ hold414/X _4580_/X _4805_/S vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7587_ _7587_/CLK _7587_/D vssd1 vssd1 vccd1 vccd1 _7587_/Q sky130_fd_sc_hd__dfxtp_1
X_6538_ _6435_/Y _6441_/Y _6475_/X _6477_/X _6521_/A vssd1 vssd1 vccd1 vccd1 _6538_/Y
+ sky130_fd_sc_hd__a41oi_1
XANTENNA__5107__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6469_ _6468_/A _6468_/B _6506_/B _6453_/X vssd1 vssd1 vccd1 vccd1 _6498_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4373__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7032__A1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3778__A _7543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5696__C _6338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7099__A1 _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7099__B2 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5988__C_N _5811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4548__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__B _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6329__A _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6048__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4283__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5379__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5840_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5841_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5771_ _6691_/A _6738_/A _6683_/B _6629_/A vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__or4_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7510_ _7537_/CLK hold43/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4722_ _3682_/Y _4724_/S _3763_/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__a21boi_1
X_7441_ _7441_/CLK _7441_/D vssd1 vssd1 vccd1 vccd1 _7441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5337__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4653_ _5024_/S _4698_/C vssd1 vssd1 vccd1 vccd1 _4654_/A sky130_fd_sc_hd__or2_1
XFILLER_0_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput40 io_in[26] vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__clkbuf_1
X_7372_ _7372_/CLK _7372_/D vssd1 vssd1 vccd1 vccd1 _7372_/Q sky130_fd_sc_hd__dfxtp_1
X_4584_ _6148_/A _4632_/C vssd1 vssd1 vccd1 vccd1 _4585_/B sky130_fd_sc_hd__and2_1
XFILLER_0_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6323_ _6238_/X _7110_/B _6276_/B vssd1 vssd1 vccd1 vccd1 _7121_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6254_ _6264_/A _6319_/A vssd1 vssd1 vccd1 vccd1 _6978_/B sky130_fd_sc_hd__nor2_2
X_5205_ hold361/X _4964_/X _5211_/S vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4848__A0 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6239__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6185_ _6185_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6185_/X sky130_fd_sc_hd__or2_1
X_5136_ input32/X _6225_/B _5135_/X _6373_/A vssd1 vssd1 vccd1 vccd1 _7361_/D sky130_fd_sc_hd__o211a_1
X_5067_ hold611/X _4937_/Y _5075_/S vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4982__A _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4076__B2 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4018_ _4021_/A _3741_/B _6357_/A _4017_/X _6015_/A vssd1 vssd1 vccd1 vccd1 _4067_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7014__B2 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7014__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5025__B1 _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5969_ _5960_/A _5958_/Y _6236_/A vssd1 vssd1 vccd1 vccd1 _5970_/D sky130_fd_sc_hd__o21ba_1
XANTENNA__6702__A _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5981__D1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6421__B _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5988__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5199__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4831__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6612__A _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5319__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold109 _7549_/Q vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6819__A1 _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7229__D1 _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4058__B2 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6941_ _6875_/B _6875_/C split4/A _7043_/S vssd1 vssd1 vccd1 vccd1 _6941_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5007__A0 _4238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6872_ _6872_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _6872_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5558__A1 _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5823_ _5825_/D vssd1 vssd1 vccd1 vccd1 _5823_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4026__B _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4741__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_wb_clk_i _7544_/CLK vssd1 vssd1 vccd1 vccd1 _7536_/CLK sky130_fd_sc_hd__clkbuf_16
X_5754_ _6630_/A _6808_/B _5751_/Y _5766_/A vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__o22a_1
X_4705_ _7283_/Q _7598_/Q _7267_/Q _7491_/Q _7340_/Q _7341_/Q vssd1 vssd1 vccd1 vccd1
+ _4705_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6241__B _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5685_ _5654_/A _5740_/A _5683_/X _5684_/Y vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__a211oi_2
X_7424_ _7424_/CLK _7424_/D vssd1 vssd1 vccd1 vccd1 _7424_/Q sky130_fd_sc_hd__dfxtp_1
X_4636_ _3933_/A _4635_/X _4634_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _4637_/B sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout213_A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5138__A _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7355_ _7423_/CLK _7355_/D vssd1 vssd1 vccd1 vccd1 _7355_/Q sky130_fd_sc_hd__dfxtp_1
Xhold621 _7344_/Q vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5730__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold610 _6807_/A vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__clkbuf_2
X_4567_ _4566_/X _4565_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4568_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold654 _7586_/Q vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 _6398_/X vssd1 vssd1 vccd1 vccd1 _7575_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _6338_/A _6306_/B vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__nor2_1
Xhold643 _7589_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _4496_/X _4497_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__mux2_1
X_7286_ _7618_/CLK _7286_/D vssd1 vssd1 vccd1 vccd1 _7286_/Q sky130_fd_sc_hd__dfxtp_1
Xhold665 _7472_/Q vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6237_ _7137_/A vssd1 vssd1 vccd1 vccd1 _6282_/A sky130_fd_sc_hd__inv_2
XANTENNA__5304__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6167_/X hold88/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
X_5119_ hold373/X _4912_/Y _5129_/S vssd1 vssd1 vccd1 vccd1 _5119_/X sky130_fd_sc_hd__mux2_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7235__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5246__A0 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6099_ _7600_/Q _6153_/A _6098_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6100_/B sky130_fd_sc_hd__a211o_1
XANTENNA__4049__A1 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6994__B1 _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5974__C _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3791__A _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4288__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5214__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6682__C1 _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7226__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7202__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6985__B1 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6326__B _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5470_ _5471_/B _5471_/C _6518_/A vssd1 vssd1 vccd1 vccd1 _5470_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4421_ _4420_/X _4419_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5392__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4352_ _4474_/A _6044_/B _4351_/X vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7140_ _5800_/C _7136_/X _7558_/Q vssd1 vssd1 vccd1 vccd1 _7140_/Y sky130_fd_sc_hd__o21ai_1
X_4283_ _4281_/X _4282_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__mux2_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7071_ _7072_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7071_/X sky130_fd_sc_hd__or2_1
X_6022_ _6427_/B _6022_/B vssd1 vssd1 vccd1 vccd1 _6022_/Y sky130_fd_sc_hd__nor2_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7217__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4736__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6517__A _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6951__S _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4037__A _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6924_ _6220_/B _6919_/Y _6920_/X _3761_/B _4013_/Y vssd1 vssd1 vccd1 vccd1 _6925_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3885__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4471__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3876__A _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6855_ _6791_/Y _6854_/Y _6891_/B vssd1 vssd1 vccd1 vccd1 _7029_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5400__A0 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3998_ _6920_/A _7473_/Q vssd1 vssd1 vccd1 vccd1 _4121_/B sky130_fd_sc_hd__nor2_2
X_5806_ _3973_/B _4081_/A _5805_/X _7043_/S vssd1 vssd1 vccd1 vccd1 _5810_/C sky130_fd_sc_hd__o22a_1
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6786_ _6786_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6786_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__6252__A _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5951__A1 _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5737_ _5737_/A vssd1 vssd1 vccd1 vccd1 _5757_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7407_ _7439_/CLK _7407_/D vssd1 vssd1 vccd1 vccd1 _7407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _6808_/A _6771_/A _6773_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _5671_/D sky130_fd_sc_hd__a22o_1
X_4619_ _4618_/X _4617_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4620_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5599_ _5615_/A _5615_/B vssd1 vssd1 vccd1 vccd1 _6451_/A sky130_fd_sc_hd__or2_1
Xhold440 _5399_/X vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7338_ _7450_/CLK _7338_/D vssd1 vssd1 vccd1 vccd1 _7338_/Q sky130_fd_sc_hd__dfxtp_1
Xhold462 _7423_/Q vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _7446_/Q vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold484 _7432_/Q vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _4795_/X vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
X_7269_ _7372_/CLK _7269_/D vssd1 vssd1 vccd1 vccd1 _7269_/Q sky130_fd_sc_hd__dfxtp_1
Xhold495 _7275_/Q vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7208__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6427__A _6427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6967__B1 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4442__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6162__A _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7144__B1 _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7624_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3800__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output57_A _7558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7080__C1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _7025_/A _4945_/B _4968_/X _4969_/Y _4946_/A vssd1 vssd1 vccd1 vccd1 _4970_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5387__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3921_ _3935_/A _4487_/A vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__nor2_1
X_3852_ _7438_/Q _7430_/Q _7414_/Q _7406_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3852_/X sky130_fd_sc_hd__mux4_1
X_6640_ _6640_/A _6640_/B vssd1 vssd1 vccd1 vccd1 _6670_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6571_ _6524_/B _6570_/X _7090_/B vssd1 vssd1 vccd1 vccd1 _6573_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4292__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4304__B _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5522_ _5497_/A _5521_/X _5528_/S vssd1 vssd1 vccd1 vccd1 _5524_/B sky130_fd_sc_hd__mux2_4
X_3783_ hold97/X _4034_/B vssd1 vssd1 vccd1 vccd1 _6415_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5453_ _5452_/A _5452_/B _5452_/C _5451_/Y vssd1 vssd1 vccd1 vccd1 _5454_/C sky130_fd_sc_hd__a31o_4
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5384_ hold297/X _4492_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7479_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4320__A _4320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4404_ _4407_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__or2_1
Xfanout205 _7340_/Q vssd1 vssd1 vccd1 vccd1 _4709_/S0 sky130_fd_sc_hd__buf_8
X_4335_ _4334_/X _4360_/B vssd1 vssd1 vccd1 vccd1 _4335_/Y sky130_fd_sc_hd__nand2b_1
X_7123_ _7123_/A _7123_/B _7123_/C vssd1 vssd1 vccd1 vccd1 _7123_/X sky130_fd_sc_hd__and3_1
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7631__A _7631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6110__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6110__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4266_ _4269_/A _4876_/B vssd1 vssd1 vccd1 vccd1 _4266_/Y sky130_fd_sc_hd__nor2_1
X_7054_ _7072_/B _6307_/B _7053_/Y vssd1 vssd1 vccd1 vccd1 _7054_/X sky130_fd_sc_hd__a21o_1
X_4197_ _4689_/A _4195_/X _4196_/Y _4192_/Y vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6005_ _3754_/X _6008_/B _3749_/Y vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__o21ba_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6907_ _6301_/A _7123_/B _7123_/C _6922_/B _6244_/A vssd1 vssd1 vccd1 vccd1 _6907_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6838_ _6838_/A _6838_/B vssd1 vssd1 vccd1 vccd1 _6838_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__7078__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6769_ _6789_/A _6766_/Y _6767_/Y _6768_/X vssd1 vssd1 vccd1 vccd1 _6823_/A sky130_fd_sc_hd__a211oi_1
XFILLER_0_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6710__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold270 _5292_/X vssd1 vssd1 vccd1 vccd1 _7430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _7387_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _4813_/X vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6101__B2 _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6157__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4663__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4415__A1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4405__A _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7117__B1 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ _4267_/C _4121_/B _4134_/D vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__and3_2
XANTENNA__4286__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4051_ _7569_/Q _6882_/A _6023_/S vssd1 vssd1 vccd1 vccd1 _4051_/X sky130_fd_sc_hd__mux2_1
Xinput5 custom_settings[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
XFILLER_0_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5603__B1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4501__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4953_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6800__C1 _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3904_ _7478_/Q _7466_/Q _7458_/Q _7252_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3904_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4884_ _4349_/A _4861_/B _5034_/B vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6623_ _6585_/Y _6622_/Y split9/A vssd1 vssd1 vccd1 vccd1 _6625_/B sky130_fd_sc_hd__mux2_2
X_3835_ _7363_/Q _3833_/X _3834_/Y _3829_/Y vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3766_ _6096_/A _7550_/Q vssd1 vssd1 vccd1 vccd1 _4290_/B sky130_fd_sc_hd__or2_1
X_6554_ _6754_/A _6556_/B vssd1 vssd1 vccd1 vccd1 _6597_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4590__B1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5505_ split8/X _5500_/B hold86/A vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6485_ _6485_/A _6485_/B _6485_/C _6485_/D vssd1 vssd1 vccd1 vccd1 _6486_/B sky130_fd_sc_hd__and4_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5436_ _7497_/Q _6683_/B vssd1 vssd1 vccd1 vccd1 _5437_/B sky130_fd_sc_hd__nand2_1
X_3697_ _7555_/Q _7554_/Q vssd1 vssd1 vccd1 vccd1 _3992_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5367_ hold474/X _4580_/X _5373_/S vssd1 vssd1 vccd1 vccd1 _5367_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5298_ _5297_/X _4973_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__mux2_1
X_4318_ _4360_/B _4318_/B vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__and2b_1
X_7106_ _5988_/A _6157_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _7106_/X sky130_fd_sc_hd__a21o_1
X_4249_ _5026_/A _5026_/B vssd1 vssd1 vccd1 vccd1 _5027_/A sky130_fd_sc_hd__or2_1
X_7037_ _6249_/A _7008_/B _6279_/B vssd1 vssd1 vccd1 vccd1 _7039_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__B _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5070__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3908__B1 _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6440__A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4636__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4834__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7210__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6615__A _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5061__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3974__A _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6270_ _7137_/A _7137_/B vssd1 vssd1 vccd1 vccd1 _6270_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6313__A1 _7551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5221_ hold517/X _4937_/Y _5229_/S vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5152_ _4947_/X hold561/X _5158_/S vssd1 vssd1 vccd1 vccd1 _7368_/D sky130_fd_sc_hd__mux2_1
X_4103_ _4103_/A _5019_/A vssd1 vssd1 vccd1 vccd1 _4389_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ hold557/X _4912_/Y _5093_/S vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__mux2_1
X_4034_ _6421_/B _4034_/B vssd1 vssd1 vccd1 vccd1 _4034_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4744__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5052__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6244__B _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5985_ _5985_/A _5985_/B vssd1 vssd1 vccd1 vccd1 _5985_/Y sky130_fd_sc_hd__nand2_1
X_4936_ _7347_/Q _4166_/B _4964_/S vssd1 vssd1 vccd1 vccd1 _4936_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4867_ _4867_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4868_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3818_ _3816_/X _3817_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3818_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7586_ _7587_/CLK _7586_/D vssd1 vssd1 vccd1 vccd1 _7586_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6260__A _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6606_ _6771_/A _6606_/B vssd1 vssd1 vccd1 vccd1 _6648_/A sky130_fd_sc_hd__xnor2_2
X_4798_ _4492_/X hold343/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7287_/D sky130_fd_sc_hd__mux2_1
X_6537_ _6483_/Y _6490_/X _6482_/Y vssd1 vssd1 vccd1 vccd1 _6540_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3749_ _6216_/A _6216_/B vssd1 vssd1 vccd1 vccd1 _3749_/Y sky130_fd_sc_hd__nor2_1
X_6468_ _6468_/A _6468_/B _6506_/B vssd1 vssd1 vccd1 vccd1 _6468_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3823__S _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5419_ _5818_/B _5854_/C _6702_/A split8/A vssd1 vssd1 vccd1 vccd1 _5955_/D sky130_fd_sc_hd__or4_4
X_6399_ hold126/X _6415_/A _6356_/B hold213/X vssd1 vssd1 vccd1 vccd1 _6399_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4866__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6068__A0 _6067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5815__B1 _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5042__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5043__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4829__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7205__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__A0 _6058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4564__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6345__A _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _6690_/A _6802_/A _6802_/B _5788_/D vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__and4_1
X_4721_ _4685_/X _4720_/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7257_/D sky130_fd_sc_hd__mux2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5395__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7440_ _7449_/CLK _7440_/D vssd1 vssd1 vccd1 vccd1 _7440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7176__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6080__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4652_ _4602_/X _4698_/C _4695_/A vssd1 vssd1 vccd1 vccd1 _4652_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 custom_settings[9] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
X_7371_ _7443_/CLK _7371_/D vssd1 vssd1 vccd1 vccd1 _7371_/Q sky130_fd_sc_hd__dfxtp_1
X_4583_ _6148_/A _4632_/C vssd1 vssd1 vccd1 vccd1 _4633_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput41 io_in[27] vssd1 vssd1 vccd1 vccd1 _3679_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6322_ _7092_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _7110_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4739__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6253_ _6738_/A _6799_/A vssd1 vssd1 vccd1 vccd1 _6253_/Y sky130_fd_sc_hd__nand2_1
X_5204_ _4921_/X _5203_/X _5212_/S vssd1 vssd1 vccd1 vccd1 _7391_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4848__A1 _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5424__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6184_ hold68/X hold38/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6239__B _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_A _7360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5135_ _6326_/B _6229_/S vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _5065_/X _4897_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5273__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4017_ _4267_/D _4015_/Y _4016_/Y _6374_/A vssd1 vssd1 vccd1 vccd1 _4017_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7014__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5025__A1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ hold78/X wire79/X _5967_/X _6218_/A vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__o211a_1
XFILLER_0_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4919_ _6962_/A _4945_/B _4917_/X _4918_/Y vssd1 vssd1 vccd1 vccd1 _4919_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3818__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5899_ _5927_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5901_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6421__C _6427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7569_ _7569_/CLK _7569_/D vssd1 vssd1 vccd1 vccd1 _7569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4839__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5264__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5805__C_N _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5509__A _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5972__C1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6104__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4413__A _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5255__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4294__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6940_ split4/X _6940_/B vssd1 vssd1 vccd1 vccd1 _6940_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6075__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6871_ _6871_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6968_/A sky130_fd_sc_hd__xnor2_2
X_5822_ _6690_/A _6771_/A _6773_/A _6802_/A vssd1 vssd1 vccd1 vccd1 _5825_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5753_ _5751_/Y _5766_/A _6683_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _5766_/B sky130_fd_sc_hd__and4bb_1
XANTENNA__4026__C _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4704_ _3677_/Y _4982_/A _4701_/X _4703_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4704_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5419__A _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5684_ _5684_/A _5684_/B vssd1 vssd1 vccd1 vccd1 _5684_/Y sky130_fd_sc_hd__nor2_1
X_7423_ _7423_/CLK _7423_/D vssd1 vssd1 vccd1 vccd1 _7423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7180__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4635_ _6157_/A _3924_/B _4107_/Y vssd1 vssd1 vccd1 vccd1 _4635_/X sky130_fd_sc_hd__o21a_1
Xhold611 _7327_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _7272_/Q _7612_/Q _7604_/Q _7620_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4566_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7354_ _7453_/CLK _7354_/D vssd1 vssd1 vccd1 vccd1 _7354_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout206_A _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold600 _4724_/X vssd1 vssd1 vccd1 vccd1 _7259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 _7600_/Q vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold633 _7346_/Q vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4977__B _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6305_ _7040_/A _6989_/B _7040_/B vssd1 vssd1 vccd1 vccd1 _6306_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5730__A2 _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold644 _7590_/Q vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _7479_/Q _7467_/Q _7459_/Q _7253_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4497_/X sky130_fd_sc_hd__mux4_1
X_7285_ _7477_/CLK _7285_/D vssd1 vssd1 vccd1 vccd1 _7285_/Q sky130_fd_sc_hd__dfxtp_1
Xhold655 _7348_/Q vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _7345_/Q vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ _6236_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _7137_/A sky130_fd_sc_hd__nand2_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4993__A _6084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6167_ _6427_/B _6165_/X _6166_/Y _4699_/A _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6167_/X
+ sky130_fd_sc_hd__o32a_1
X_5118_ hold278/X _4871_/Y _5130_/S vssd1 vssd1 vccd1 vccd1 _7353_/D sky130_fd_sc_hd__mux2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6098_ _6153_/A _6098_/B vssd1 vssd1 vccd1 vccd1 _6098_/Y sky130_fd_sc_hd__nor2_1
X_5049_ hold256/X _4937_/Y _5057_/S vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5954__C1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5182__A0 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5237__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6326__C _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4996__B1 _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4842__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7162__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _7269_/Q _7609_/Q _7601_/Q _7617_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4420_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4351_ _4351_/A _4351_/B vssd1 vssd1 vccd1 vccd1 _4351_/X sky130_fd_sc_hd__and2_1
X_4282_ _7476_/Q _7464_/Q _7456_/Q _7250_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4282_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7070_ _7070_/A _7109_/A vssd1 vssd1 vccd1 vccd1 _7078_/C sky130_fd_sc_hd__nor2_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _7169_/A _7171_/A _6021_/C vssd1 vssd1 vccd1 vccd1 _6086_/S sky130_fd_sc_hd__or3_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5228__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6425__B1 _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4037__B _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6923_ _4021_/A _5979_/A _5979_/B _6922_/X _4036_/A vssd1 vssd1 vccd1 vccd1 _6925_/C
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3885__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6189__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout156_A _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6854_ _6854_/A _6854_/B vssd1 vssd1 vccd1 vccd1 _6854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5805_ _5805_/A _6920_/A _4037_/A vssd1 vssd1 vccd1 vccd1 _5805_/X sky130_fd_sc_hd__or3b_1
XANTENNA__5936__C1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3997_ hold56/X _5990_/A _5985_/A _3996_/X _6922_/A vssd1 vssd1 vccd1 vccd1 _3997_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6252__B _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6785_ _6789_/A _6789_/B _6732_/Y vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5736_ _5736_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _5737_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7153__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667_ _6273_/A _5818_/B _5664_/Y _5665_/X vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__o2bb2a_1
X_7406_ _7430_/CLK _7406_/D vssd1 vssd1 vccd1 vccd1 _7406_/Q sky130_fd_sc_hd__dfxtp_1
X_4618_ _7273_/Q _7613_/Q _7605_/Q _7621_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4618_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5598_ _6799_/A _5598_/B _5598_/C vssd1 vssd1 vccd1 vccd1 _5615_/B sky130_fd_sc_hd__and3_1
Xhold441 _7485_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _7457_/Q vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
X_7337_ _7451_/CLK _7337_/D vssd1 vssd1 vccd1 vccd1 _7337_/Q sky130_fd_sc_hd__dfxtp_1
X_4549_ _3668_/Y _4548_/X _4545_/X vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__a21oi_4
Xhold452 _5328_/X vssd1 vssd1 vccd1 vccd1 _7446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _7450_/Q vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _7468_/Q vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _7252_/Q vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _5295_/X vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
X_7268_ _7621_/CLK _7268_/D vssd1 vssd1 vccd1 vccd1 _7268_/Q sky130_fd_sc_hd__dfxtp_1
X_6219_ _4084_/A hold97/X _3962_/D _6911_/A vssd1 vssd1 vccd1 vccd1 _6220_/D sky130_fd_sc_hd__a211o_1
X_7199_ hold219/X _4483_/X _7209_/S vssd1 vssd1 vccd1 vccd1 _7199_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5612__A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5219__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6427__B _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4228__A _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3953__A1 hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3800__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4837__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7213__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6407__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6958__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4138__A _5811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7080__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _3665_/Y _3917_/Y _3918_/X _3912_/X vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3851_ _7363_/Q _3849_/X _3850_/Y _3845_/Y vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__a2bb2o_2
XANTENNA__3696__B _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6570_ _6570_/A _6570_/B vssd1 vssd1 vccd1 vccd1 _6570_/X sky130_fd_sc_hd__and2_1
X_3782_ _6326_/B _3962_/C vssd1 vssd1 vccd1 vccd1 _4034_/B sky130_fd_sc_hd__or2_2
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4292__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5521_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5146__A0 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7135__A1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _5452_/A _5452_/B _5452_/C vssd1 vssd1 vccd1 vccd1 _5452_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5383_ hold296/X _4529_/X _5391_/S vssd1 vssd1 vccd1 vccd1 _5383_/X sky130_fd_sc_hd__mux2_1
X_4403_ _4407_/B vssd1 vssd1 vccd1 vccd1 _4403_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4334_ _4332_/X _4333_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4334_/X sky130_fd_sc_hd__mux2_1
X_7122_ _7122_/A _7122_/B vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__or2_1
Xfanout206 _6204_/A vssd1 vssd1 vccd1 vccd1 _7244_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7053_ _7072_/B _6307_/B _6989_/A vssd1 vssd1 vccd1 vccd1 _7053_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4207__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4265_ _4876_/B vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__inv_2
X_6004_ _6004_/A _6004_/B _6004_/C _6004_/D vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__or4_4
X_4196_ _4401_/S _4190_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4196_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4482__S _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6906_ _4862_/A _5804_/C _6429_/Y _6905_/Y _6326_/C vssd1 vssd1 vccd1 vccd1 _6906_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6837_ _6862_/B _6874_/C vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7487_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6768_ _6857_/A _6717_/Y _6722_/B _6716_/Y vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3826__S _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6699_ _6699_/A _6699_/B vssd1 vssd1 vccd1 vccd1 _6699_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5719_ _5658_/X _5662_/A _5843_/A _5718_/X vssd1 vssd1 vccd1 vccd1 _5843_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold271 _7373_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _7322_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold293 _5193_/X vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _7448_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6101__A2 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6157__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4663__A2 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7208__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6325__C1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6876__B1 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4567__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ _4049_/X hold213/X _7241_/S vssd1 vssd1 vccd1 vccd1 _4050_/X sky130_fd_sc_hd__mux2_1
Xinput6 custom_settings[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_1
XFILLER_0_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7053__B1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5398__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4406__A2 _4407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4952_ _6793_/A _4976_/B _5008_/A vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__a21o_1
X_3903_ _3915_/A _3903_/B vssd1 vssd1 vccd1 vccd1 _3903_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4883_ input12/X _4882_/X _5031_/S vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold94_A hold94/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3834_ _3915_/A _3830_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _3834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6622_ _6622_/A _6622_/B vssd1 vssd1 vccd1 vccd1 _6622_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3917__A1 _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6553_ _6556_/B vssd1 vssd1 vccd1 vccd1 _6553_/Y sky130_fd_sc_hd__inv_2
X_3765_ _7230_/A _4036_/A vssd1 vssd1 vccd1 vccd1 _3780_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4331__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5504_ _5504_/A _5504_/B vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__nor2_1
X_3696_ _7555_/Q _7554_/Q vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__and2_1
X_6484_ _6840_/A _6484_/B vssd1 vssd1 vccd1 vccd1 _6535_/A sky130_fd_sc_hd__xnor2_1
X_5435_ _5818_/B _5455_/B vssd1 vssd1 vccd1 vccd1 _5452_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout119_A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5366_ _4492_/X hold207/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7467_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5297_ hold284/X _4990_/Y _5301_/S vssd1 vssd1 vccd1 vccd1 _5297_/X sky130_fd_sc_hd__mux2_1
X_4317_ _4316_/X _4315_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__mux2_1
X_7105_ _7089_/X _7103_/X _7104_/X vssd1 vssd1 vccd1 vccd1 _7105_/Y sky130_fd_sc_hd__o21ai_1
X_4248_ _5026_/B vssd1 vssd1 vccd1 vccd1 _4248_/Y sky130_fd_sc_hd__inv_2
X_7036_ _7020_/A _6267_/B _7035_/X _3946_/Y _6338_/A vssd1 vssd1 vccd1 vccd1 _7044_/C
+ sky130_fd_sc_hd__a32o_1
X_4179_ _4689_/A _4177_/X _4178_/Y _4173_/Y vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__a2bb2o_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6721__A _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3908__A1 _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4581__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4241__A _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4387__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5597__B1 _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4789__C _4789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5220_ hold369/X _4897_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3990__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6313__A2 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4297__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5151_ hold560/X _4964_/X _5157_/S vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__mux2_1
X_5082_ hold581/X _4871_/Y _5094_/S vssd1 vssd1 vccd1 vccd1 _7333_/D sky130_fd_sc_hd__mux2_1
X_4102_ _6093_/A _5018_/B vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__nor2_1
X_4033_ _4065_/C _4033_/B vssd1 vssd1 vccd1 vccd1 _4033_/X sky130_fd_sc_hd__or2_1
XANTENNA__4183__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7026__B1 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3930__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5984_ _5977_/B _6220_/B _4280_/B _4065_/C _4011_/X vssd1 vssd1 vccd1 vccd1 _6925_/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4760__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4935_ _4162_/B _4934_/X _4932_/X _4964_/S vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4866_ hold172/X _4849_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _7308_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3817_ _7269_/Q _7609_/Q _7601_/Q _7617_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3817_/X sky130_fd_sc_hd__mux4_1
X_4797_ hold342/X _4529_/X _4805_/S vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7585_ _7587_/CLK _7585_/D vssd1 vssd1 vccd1 vccd1 _7585_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6260__B _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6605_ _6754_/A _6606_/B vssd1 vssd1 vccd1 vccd1 _6605_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4061__A _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6536_ _6531_/A _6531_/B _6535_/Y vssd1 vssd1 vccd1 vccd1 _6583_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3748_ _6920_/A _5132_/B _6920_/D vssd1 vssd1 vccd1 vccd1 _3762_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3679_ _3679_/A vssd1 vssd1 vccd1 vccd1 _7545_/D sky130_fd_sc_hd__inv_2
X_6467_ _6742_/A _6467_/B vssd1 vssd1 vccd1 vccd1 _6506_/B sky130_fd_sc_hd__and2_1
X_5418_ _5818_/B _5438_/A vssd1 vssd1 vccd1 vccd1 _5418_/Y sky130_fd_sc_hd__nor2_1
X_6398_ _6397_/X hold631/X _6414_/S vssd1 vssd1 vccd1 vccd1 _6398_/X sky130_fd_sc_hd__mux2_1
X_5349_ hold523/X _4580_/X _5355_/S vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5604__B _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5815__A1 _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5815__B2 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4079__B1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4174__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7019_ _7019_/A _7019_/B vssd1 vssd1 vccd1 vccd1 _7020_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold615_A _7559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4670__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5806__B2 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7221__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6626__A _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4146__A _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4720_ hold582/X _4719_/Y _4720_/S vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__mux2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4651_ _4999_/B _4651_/B vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__nor2_1
Xinput20 custom_settings[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput31 io_in[11] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
X_4582_ _4538_/X _4581_/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7254_/D sky130_fd_sc_hd__mux2_1
X_7370_ _7443_/CLK _7370_/D vssd1 vssd1 vccd1 vccd1 _7370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 io_in[28] vssd1 vssd1 vccd1 vccd1 _3680_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6321_ _7066_/A _7022_/B _7072_/B _6295_/A vssd1 vssd1 vccd1 vccd1 _6322_/B sky130_fd_sc_hd__o211a_1
X_6252_ _6935_/A _6871_/A vssd1 vssd1 vccd1 vccd1 _6319_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5203_ hold402/X _4937_/Y _5211_/S vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6183_ _3751_/Y _6181_/X _6182_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6183_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5134_ input31/X _6225_/B _5133_/Y _6373_/A vssd1 vssd1 vccd1 vccd1 _7360_/D sky130_fd_sc_hd__o211a_1
XANTENNA_fanout186_A _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4755__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5065_ hold412/X _4912_/Y _5075_/S vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3879__B _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6470__A1 _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4016_ _4021_/A _4122_/C _6374_/B vssd1 vssd1 vccd1 vccd1 _4016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4056__A _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5967_ _6581_/A _5811_/Y _5966_/Y _5811_/A _5810_/X vssd1 vssd1 vccd1 vccd1 _5967_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4784__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4918_ _4945_/B _4942_/B vssd1 vssd1 vccd1 vccd1 _4918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _5898_/A _5898_/B _5898_/C vssd1 vssd1 vccd1 vccd1 _5899_/B sky130_fd_sc_hd__nor3_1
X_4849_ _5022_/A _4849_/B vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__or2_4
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_7568_ _7569_/CLK _7568_/D vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7499_ _7538_/CLK _7499_/D vssd1 vssd1 vccd1 vccd1 _7499_/Q sky130_fd_sc_hd__dfxtp_1
X_6519_ _6581_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _6576_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4395__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout99_A _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4298__A_N _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4775__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7216__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__C1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6356__A _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3699__B _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6075__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4463__B1 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6870_ _6864_/B _6864_/C _6864_/A vssd1 vssd1 vccd1 vccd1 _6870_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5821_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5829_/A sky130_fd_sc_hd__or2_1
XANTENNA__4766__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5752_ _6690_/A _6807_/A _5774_/A vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__and3_1
X_4703_ _4701_/D _4702_/Y _5031_/S _4697_/X vssd1 vssd1 vccd1 vccd1 _4703_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5419__B _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5683_ _5684_/A _5684_/B vssd1 vssd1 vccd1 vccd1 _5683_/X sky130_fd_sc_hd__and2_2
X_7422_ _7454_/CLK _7422_/D vssd1 vssd1 vccd1 vccd1 _7422_/Q sky130_fd_sc_hd__dfxtp_1
X_4634_ _6581_/A _4440_/A _4440_/Y _4633_/Y vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5191__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4565_ _7376_/Q _7304_/Q _7296_/Q _7288_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4565_/X sky130_fd_sc_hd__mux4_1
X_7353_ _7453_/CLK _7353_/D vssd1 vssd1 vccd1 vccd1 _7353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold601 _7529_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold612 _7539_/Q vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold623 _7350_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold645 _7607_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5435__A _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6304_ _7009_/A _6960_/B _7009_/B vssd1 vssd1 vccd1 vccd1 _6989_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout101_A _3705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 _7553_/Q vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__clkbuf_2
X_4496_ _7279_/Q _7594_/Q _7263_/Q _7487_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4496_/X sky130_fd_sc_hd__mux4_1
X_7284_ _7476_/CLK _7284_/D vssd1 vssd1 vccd1 vccd1 _7284_/Q sky130_fd_sc_hd__dfxtp_1
Xhold656 _7602_/Q vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 _4898_/Y vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6235_ _6235_/A _6827_/A vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__or2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6166_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4485__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5117_ hold277/X _4887_/X _5129_/S vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__mux2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6096_/A _4180_/Y _6025_/Y _6096_/Y vssd1 vssd1 vccd1 vccd1 _6100_/A sky130_fd_sc_hd__a211o_1
XANTENNA__7235__A3 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5048_ _5047_/X _4897_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _7318_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4206__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold146_A _7522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4301__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4757__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6205__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6999_ split4/X _6999_/B vssd1 vssd1 vccd1 vccd1 _6999_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4368__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6131__B1 _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4424__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3971__A2 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5173__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3982__B _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6370__A0 _7529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4350_ _4474_/A _6035_/B _4349_/Y vssd1 vssd1 vccd1 vccd1 _4351_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__4920__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4281_ _7276_/Q _7591_/Q _7260_/Q _7484_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4281_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _7169_/B _6020_/B _6020_/C _7170_/B vssd1 vssd1 vccd1 vccd1 _6021_/C sky130_fd_sc_hd__or4b_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4436__A0 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4987__B2 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6922_ _6922_/A _6922_/B _6922_/C _6922_/D vssd1 vssd1 vccd1 vccd1 _6922_/X sky130_fd_sc_hd__or4_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6853_ _6813_/B _6813_/C _6813_/A vssd1 vssd1 vccd1 vccd1 _6854_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4739__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5804_ _6220_/B _5804_/B _5804_/C _5804_/D vssd1 vssd1 vccd1 vccd1 _5810_/B sky130_fd_sc_hd__or4_1
XFILLER_0_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6784_ _6851_/A _6784_/B vssd1 vssd1 vccd1 vccd1 _6841_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout149_A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3996_ _7539_/Q _4723_/A _3742_/C vssd1 vssd1 vccd1 vccd1 _3996_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _5634_/A _5634_/B _5634_/C vssd1 vssd1 vccd1 vccd1 _5736_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5666_ _5665_/X _5818_/B _6628_/A _5666_/D vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__and4b_1
X_7405_ _7449_/CLK _7405_/D vssd1 vssd1 vccd1 vccd1 _7405_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5164__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4617_ _7377_/Q _7305_/Q _7297_/Q _7289_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4617_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold420 _5316_/X vssd1 vssd1 vccd1 vccd1 _7441_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5597_ _5598_/B _5598_/C _5818_/B vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__a21o_1
Xhold442 _7431_/Q vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _7477_/Q vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
X_7336_ _7451_/CLK _7336_/D vssd1 vssd1 vccd1 vccd1 _7336_/Q sky130_fd_sc_hd__dfxtp_1
X_4548_ _4546_/X _4547_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4548_/X sky130_fd_sc_hd__mux2_1
Xhold431 _5335_/X vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4911__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7267_ _7598_/CLK _7267_/D vssd1 vssd1 vccd1 vccd1 _7267_/Q sky130_fd_sc_hd__dfxtp_1
Xhold475 _7282_/Q vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _7365_/Q vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _7299_/Q vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _4479_/A _4479_/B vssd1 vssd1 vccd1 vccd1 _4525_/B sky130_fd_sc_hd__or2_1
Xhold497 _4484_/X vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6218_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _7542_/D sky130_fd_sc_hd__and2_1
X_7198_ _7197_/X _4394_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7609_/D sky130_fd_sc_hd__mux2_1
X_6149_ _6427_/B _6147_/X _6148_/Y _4600_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6149_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4978__B2 _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5155__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6352__B1 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6407__B2 hold601/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__A1 _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7080__A1 _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7080__B2 _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _3915_/A _3846_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _3850_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ _6326_/B _3962_/C vssd1 vssd1 vccd1 vccd1 _6383_/B sky130_fd_sc_hd__nor2_2
X_5520_ _5553_/B _5520_/B _5520_/C vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__and3_1
XFILLER_0_42_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7135__A2 _6481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4601__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5451_ _5479_/B vssd1 vssd1 vccd1 vccd1 _5451_/Y sky130_fd_sc_hd__inv_2
X_5382_ hold450/X _4443_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7478_/D sky130_fd_sc_hd__mux2_1
X_4402_ _3668_/Y _4401_/X _4398_/X vssd1 vssd1 vccd1 vccd1 _4407_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__6894__A1 _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4333_ _7397_/Q _7389_/Q _7365_/Q _7381_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4333_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7121_ _7137_/A _7121_/B vssd1 vssd1 vccd1 vccd1 _7122_/B sky130_fd_sc_hd__nor2_1
X_4264_ _4127_/X _4128_/X _5974_/C vssd1 vssd1 vccd1 vccd1 _4876_/B sky130_fd_sc_hd__mux2_2
Xfanout207 _6015_/A vssd1 vssd1 vccd1 vccd1 _6373_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7052_ _7072_/B _7051_/B _7020_/A vssd1 vssd1 vccd1 vccd1 _7052_/X sky130_fd_sc_hd__o21a_1
X_6003_ _3650_/Y hold84/X _3652_/Y hold72/X _5999_/X vssd1 vssd1 vccd1 vccd1 _6004_/D
+ sky130_fd_sc_hd__a221o_1
X_4195_ _4193_/X _4194_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4763__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6905_ _6905_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6905_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6836_ _6835_/X _6836_/B _6836_/C vssd1 vssd1 vccd1 vccd1 _6874_/C sky130_fd_sc_hd__and3b_2
XANTENNA__5909__B1 _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5385__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6767_ _6734_/A _6734_/B _6766_/A _6781_/A vssd1 vssd1 vccd1 vccd1 _6767_/Y sky130_fd_sc_hd__a211oi_1
X_3979_ _4128_/A _3978_/Y _7553_/Q vssd1 vssd1 vccd1 vccd1 _3980_/C sky130_fd_sc_hd__mux2_1
X_5718_ _5814_/B _5716_/Y _5682_/A _5683_/X vssd1 vssd1 vccd1 vccd1 _5718_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6698_ _6698_/A _6698_/B vssd1 vssd1 vccd1 vccd1 _6719_/B sky130_fd_sc_hd__nor2_2
XANTENNA__5137__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5649_ _5630_/X _5634_/A _6273_/A _5788_/D vssd1 vssd1 vccd1 vccd1 _5651_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4938__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 _7321_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
X_7319_ _7446_/CLK _7319_/D vssd1 vssd1 vccd1 vccd1 _7319_/Q sky130_fd_sc_hd__dfxtp_1
Xhold261 _5055_/X vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold294 _7429_/Q vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _7302_/Q vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _5331_/X vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_3_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A _4143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4959__A1_N _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6454__A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5128__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7224__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5533__A _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6629__A _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output62_A _7259_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5300__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4149__A _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 custom_settings[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4951_ _4951_/A vssd1 vssd1 vccd1 vccd1 _4951_/Y sky130_fd_sc_hd__inv_2
X_3902_ _7278_/Q _7593_/Q _7262_/Q _7486_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3903_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _4930_/S _4877_/Y _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5367__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3833_ _3831_/X _3832_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3833_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6621_ _6621_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _6622_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3927__S _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4612__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6552_ _6501_/X _7090_/B _6550_/Y _6551_/X vssd1 vssd1 vccd1 vccd1 _6556_/B sky130_fd_sc_hd__a2bb2o_1
X_3764_ _6920_/A _3693_/Y _3763_/X vssd1 vssd1 vccd1 vccd1 _7474_/D sky130_fd_sc_hd__a21bo_1
XANTENNA__5119__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5503_ _5818_/B _5503_/B vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__nor2_1
X_3695_ _7553_/Q _5988_/A vssd1 vssd1 vccd1 vccd1 _3698_/A sky130_fd_sc_hd__or2_2
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6483_ _6710_/A _6484_/B vssd1 vssd1 vccd1 vccd1 _6483_/Y sky130_fd_sc_hd__nand2_1
X_5434_ _5433_/Y _5421_/Y _5434_/S vssd1 vssd1 vccd1 vccd1 _5455_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4758__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5365_ hold206/X _4529_/X _5373_/S vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7104_ _7123_/A _6844_/A _4037_/X _4030_/Y vssd1 vssd1 vccd1 vccd1 _7104_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5296_ hold485/X _4947_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _7432_/D sky130_fd_sc_hd__mux2_1
X_4316_ _7423_/Q _7355_/Q _7347_/Q _7327_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4316_/X sky130_fd_sc_hd__mux4_1
X_4247_ _7455_/Q _4245_/X _4246_/Y _4241_/Y vssd1 vssd1 vccd1 vccd1 _5026_/B sky130_fd_sc_hd__a2bb2o_2
X_7035_ _7040_/B _7035_/B _6265_/Y vssd1 vssd1 vccd1 vccd1 _7035_/X sky130_fd_sc_hd__or3b_1
X_4178_ _4688_/S _4174_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4178_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4802__A0 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6819_ _6844_/A _6820_/B _6784_/B _5918_/D vssd1 vssd1 vccd1 vccd1 _6819_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4869__A0 _6874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7219__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6313__A3 _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5150_ _4921_/X _5149_/X _5158_/S vssd1 vssd1 vccd1 vccd1 _7367_/D sky130_fd_sc_hd__mux2_1
X_5081_ hold580/X _4887_/X _5093_/S vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4088__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4101_ _4101_/A _4993_/B vssd1 vssd1 vccd1 vccd1 _5018_/B sky130_fd_sc_hd__nand2_1
X_4032_ _6922_/A _6326_/D vssd1 vssd1 vccd1 vccd1 _5979_/B sky130_fd_sc_hd__or2_1
XANTENNA__4183__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7026__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5202__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3930__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4607__A _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4326__B _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5983_ _5974_/X _5976_/A _5982_/Y _4021_/A vssd1 vssd1 vccd1 vccd1 _5995_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4934_ _6057_/A _4933_/Y _4986_/S vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7441_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4865_ hold171/X _4864_/X _5039_/S vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__mux2_1
X_3816_ _7373_/Q _7301_/Q _7293_/Q _7285_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3816_/X sky130_fd_sc_hd__mux4_1
X_4796_ _4443_/X hold473/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7286_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6033__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7584_ _7587_/CLK _7584_/D vssd1 vssd1 vccd1 vccd1 _7584_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout131_A _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6604_ _6561_/B _6603_/X split9/A vssd1 vssd1 vccd1 vccd1 _6606_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6535_ _6535_/A _6545_/B vssd1 vssd1 vccd1 vccd1 _6535_/Y sky130_fd_sc_hd__nand2_1
X_3747_ _3759_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _6920_/D sky130_fd_sc_hd__or2_2
XFILLER_0_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3678_ _3678_/A vssd1 vssd1 vccd1 vccd1 _7544_/D sky130_fd_sc_hd__inv_2
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6466_ _6507_/B _6466_/B vssd1 vssd1 vccd1 vccd1 _6468_/B sky130_fd_sc_hd__and2_1
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5417_ _5415_/Y _5417_/B vssd1 vssd1 vccd1 vccd1 _5955_/C sky130_fd_sc_hd__and2b_1
X_6397_ input34/X _6396_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6397_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5348_ _4492_/X hold511/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7459_/D sky130_fd_sc_hd__mux2_1
X_5279_ hold404/X _4990_/Y _5283_/S vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4079__B2 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7018_ _6962_/A _6926_/Y _7016_/Y _7017_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7586_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5815__A2 _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4174__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7017__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A _7544_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6732__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5200__A0 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4003__A1 _7542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5751__A1 _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5811__A _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6626__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4162__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4650_ _4698_/B _4698_/C vssd1 vssd1 vccd1 vccd1 _4651_/B sky130_fd_sc_hd__or2_1
XFILLER_0_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 custom_settings[28] vssd1 vssd1 vccd1 vccd1 _7630_/A sky130_fd_sc_hd__buf_2
Xinput10 custom_settings[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
X_4581_ hold434/X _4580_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__mux2_1
Xinput32 io_in[12] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 io_in[29] vssd1 vssd1 vccd1 vccd1 _3681_/A sky130_fd_sc_hd__clkbuf_1
X_6320_ _6249_/A _6993_/B _6279_/B vssd1 vssd1 vccd1 vccd1 _7022_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6089__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6251_ _6738_/A _6799_/A vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__nor2_2
X_5202_ _4897_/X hold258/X _5212_/S vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6182_ _6182_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__or2_1
XANTENNA__7247__A1 hold524/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5133_ _6421_/B _6225_/B vssd1 vssd1 vccd1 vccd1 _5133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5064_ hold378/X _4871_/Y _5076_/S vssd1 vssd1 vccd1 vccd1 _7325_/D sky130_fd_sc_hd__mux2_1
X_4015_ _6383_/A _4015_/B vssd1 vssd1 vccd1 vccd1 _4015_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout179_A _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4771__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5430__B1 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5966_ _5970_/A _5964_/Y _5970_/C _5955_/X vssd1 vssd1 vccd1 vccd1 _5966_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_75_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4917_ _4917_/A _4917_/B vssd1 vssd1 vccd1 vccd1 _4917_/X sky130_fd_sc_hd__and2_1
XFILLER_0_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5981__A1 _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5897_ _5898_/A _5898_/B _5898_/C vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__o21a_1
X_4848_ _6311_/A _4862_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4849_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ hold549/X _4580_/X _4785_/S vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6930__B1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7567_ _7579_/CLK _7567_/D vssd1 vssd1 vccd1 vccd1 _7567_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5733__A1 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7498_ _7498_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfxtp_1
X_6518_ _6518_/A _6518_/B vssd1 vssd1 vccd1 vccd1 _6575_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6449_ _5612_/B _6448_/Y _6463_/S vssd1 vssd1 vccd1 vccd1 _6471_/B sky130_fd_sc_hd__mux2_2
XANTENNA__4395__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7238__A1 hold213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6727__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold558_A _7570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4472__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4681__S _4721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5972__A1 _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4932__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6401__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3830__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5017__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7229__A1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6637__A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6356__B _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4157__A _4751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5820_ _5820_/A _5820_/B vssd1 vssd1 vccd1 vccd1 _5831_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5751_ _6690_/A _6807_/A _5774_/A vssd1 vssd1 vccd1 vccd1 _5751_/Y sky130_fd_sc_hd__a21oi_1
X_4702_ _4701_/B _4699_/Y _4658_/A vssd1 vssd1 vccd1 vccd1 _4702_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7421_ _7454_/CLK _7421_/D vssd1 vssd1 vccd1 vccd1 _7421_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5419__C _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5682_ _5682_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5684_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4633_ _6157_/A _4633_/B vssd1 vssd1 vccd1 vccd1 _4633_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4564_ _4562_/X _4563_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7352_ _7453_/CLK _7352_/D vssd1 vssd1 vccd1 vccd1 _7352_/Q sky130_fd_sc_hd__dfxtp_1
Xhold602 _4059_/X vssd1 vssd1 vccd1 vccd1 _7342_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3821__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7283_ _7597_/CLK _7283_/D vssd1 vssd1 vccd1 vccd1 _7283_/Q sky130_fd_sc_hd__dfxtp_1
Xhold624 _7351_/Q vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _6978_/A _6933_/B _6978_/B vssd1 vssd1 vccd1 vccd1 _6960_/B sky130_fd_sc_hd__a21o_1
Xhold635 _7588_/Q vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 _6209_/X vssd1 vssd1 vccd1 vccd1 _6210_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4495_ _4540_/B _4495_/B vssd1 vssd1 vccd1 vccd1 _4495_/Y sky130_fd_sc_hd__nand2_1
Xhold668 _7605_/Q vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _7192_/X vssd1 vssd1 vccd1 vccd1 _7607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _7585_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6235_/A _6827_/A vssd1 vssd1 vccd1 vccd1 _6234_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6140__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6140__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4151__A0 _7529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4766__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _3702_/Y _4699_/A _6164_/X _6022_/B _6157_/B vssd1 vssd1 vccd1 vccd1 _6165_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6547__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5116_ hold389/X _4849_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _7352_/D sky130_fd_sc_hd__mux2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6096_/A _6098_/B vssd1 vssd1 vccd1 vccd1 _6096_/Y sky130_fd_sc_hd__nor2_1
X_5047_ hold550/X _4912_/Y _5057_/S vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7489_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4206__A1 _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6998_ _6998_/A _6998_/B vssd1 vssd1 vccd1 vccd1 _6999_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4301__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5949_ _5931_/A _5932_/X _5948_/Y vssd1 vssd1 vccd1 vccd1 _5964_/B sky130_fd_sc_hd__o21a_1
X_7619_ _7623_/CLK _7619_/D vssd1 vssd1 vccd1 vccd1 _7619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4368__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6131__A1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4693__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6457__A _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4996__A2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5300__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7147__B1 _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7227__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4440__A _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4280_ _7043_/S _4280_/B _4290_/D vssd1 vssd1 vccd1 vccd1 _4986_/S sky130_fd_sc_hd__or3_4
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4684__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6921_ _6220_/B _6918_/X _4010_/Y _4113_/B vssd1 vssd1 vccd1 vccd1 _6927_/B sky130_fd_sc_hd__a2bb2o_1
X_6852_ _6882_/A _6882_/B vssd1 vssd1 vccd1 vccd1 _6852_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5210__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5803_ _5879_/A _5803_/A2 _5802_/X vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4295__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3995_ _4001_/D _7473_/Q hold56/X _3994_/X vssd1 vssd1 vccd1 vccd1 _3995_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5936__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6783_ _6722_/B _6775_/Y _6782_/X vssd1 vssd1 vccd1 vccd1 _6784_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5734_ _5763_/B _5734_/B vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__nor2_1
XANTENNA__7138__B1 _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5665_ _6683_/A _6962_/A _5854_/C _6793_/A vssd1 vssd1 vccd1 vccd1 _5665_/X sky130_fd_sc_hd__and4_1
X_7404_ _7439_/CLK _7404_/D vssd1 vssd1 vccd1 vccd1 _7404_/Q sky130_fd_sc_hd__dfxtp_1
X_4616_ _4614_/X _4615_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4616_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6041__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 _7458_/Q vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
X_7335_ _4004_/A _7335_/D vssd1 vssd1 vccd1 vccd1 _7335_/Q sky130_fd_sc_hd__dfxtp_1
X_5596_ _5598_/B _5598_/C _5818_/B vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__a21oi_1
Xhold454 _7591_/Q vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _7250_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _7384_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _7255_/Q vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _7272_/Q _7612_/Q _7604_/Q _7620_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4547_/X sky130_fd_sc_hd__mux4_1
X_7266_ _7479_/CLK _7266_/D vssd1 vssd1 vccd1 vccd1 _7266_/Q sky130_fd_sc_hd__dfxtp_1
Xhold465 _5145_/X vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _7377_/Q vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _7420_/Q vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4478_/A _4478_/B vssd1 vssd1 vccd1 vccd1 _4479_/B sky130_fd_sc_hd__and2_1
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold498 _7409_/Q vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7197_ hold200/X _4434_/Y _7209_/S vssd1 vssd1 vccd1 vccd1 _7197_/X sky130_fd_sc_hd__mux2_1
X_6217_ _6207_/S _6008_/B _6216_/X hold636/X vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6148_ _6148_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6148_/Y sky130_fd_sc_hd__nor2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6079_/A vssd1 vssd1 vccd1 vccd1 _6079_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5120__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4210__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7080__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5091__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3780_ _3780_/A _3780_/B vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__and2_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5450_ _5428_/X _5434_/S _5422_/Y vssd1 vssd1 vccd1 vccd1 _5479_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4401_ _4399_/X _4400_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4401_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4601__C _4601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6343__A1 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5381_ hold449/X _4483_/X _5391_/S vssd1 vssd1 vccd1 vccd1 _5381_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _7437_/Q _7429_/Q _7413_/Q _7405_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4332_/X sky130_fd_sc_hd__mux4_1
X_7120_ _7137_/A _6309_/Y _7119_/Y vssd1 vssd1 vccd1 vccd1 _7120_/X sky130_fd_sc_hd__o21a_1
X_4263_ _5024_/S _4263_/B vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__nor2_1
Xfanout208 _6015_/A vssd1 vssd1 vccd1 vccd1 _7245_/C1 sky130_fd_sc_hd__clkbuf_2
X_7051_ _7072_/B _7051_/B vssd1 vssd1 vccd1 vccd1 _7051_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5205__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6002_ _3650_/A _3651_/Y _3652_/A _3653_/Y _5998_/X vssd1 vssd1 vccd1 vccd1 _6004_/C
+ sky130_fd_sc_hd__a221o_1
X_4194_ _7422_/Q _7354_/Q _7346_/Q _7326_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4194_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5082__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6904_ _6311_/A _6872_/B _4037_/X _4030_/Y vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout161_A _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6835_ _6760_/X _6834_/X _6764_/X vssd1 vssd1 vccd1 vccd1 _6835_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4999__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3978_ _6223_/A _4007_/A vssd1 vssd1 vccd1 vccd1 _3978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6766_ _6766_/A _6781_/A _6786_/A _6789_/B vssd1 vssd1 vccd1 vccd1 _6766_/Y sky130_fd_sc_hd__nor4b_4
XANTENNA__6560__A _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5717_ _5682_/A _5683_/X _5814_/B _5716_/Y vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__o211ai_4
XFILLER_0_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6697_ _6869_/A _6697_/B vssd1 vssd1 vccd1 vccd1 _6698_/B sky130_fd_sc_hd__nor2_1
X_5648_ _6581_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5579_ _5524_/B _5578_/Y _5579_/S vssd1 vssd1 vccd1 vccd1 _5580_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold240 _5310_/X vssd1 vssd1 vccd1 vccd1 _7438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _7279_/Q vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _5054_/X vssd1 vssd1 vccd1 vccd1 _7321_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7318_ _7446_/CLK _7318_/D vssd1 vssd1 vccd1 vccd1 _7318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold284 _7433_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _5289_/X vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _4833_/X vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _4079_/X hold92/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7571_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4648__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5115__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6735__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5073__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4820__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4149__B _4728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 custom_settings[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XANTENNA_output55_A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5064__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4811__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4950_ _4955_/B _4922_/Y _4949_/X vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__a21bo_1
X_3901_ _6111_/A _3901_/B vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__and2_1
X_4881_ _6807_/A _4976_/B _5008_/A vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__a21o_1
XANTENNA_split27_A _6718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3832_ _7425_/Q _7357_/Q _7349_/Q _7329_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3832_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6620_ _6578_/Y _6619_/X split9/A vssd1 vssd1 vccd1 vccd1 _6637_/B sky130_fd_sc_hd__mux2_2
X_6551_ _6529_/B _6504_/Y _6558_/A _7090_/B vssd1 vssd1 vccd1 vccd1 _6551_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5502_ _5469_/Y _5495_/S _5500_/X vssd1 vssd1 vccd1 vccd1 _5504_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3763_ _3763_/A _4723_/A _4724_/S vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__or3_1
XFILLER_0_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _7553_/Q _5988_/A vssd1 vssd1 vccd1 vccd1 _4007_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6482_ _6710_/A _6484_/B vssd1 vssd1 vccd1 vccd1 _6482_/Y sky130_fd_sc_hd__nor2_1
X_5433_ _5437_/A _5433_/B vssd1 vssd1 vccd1 vccd1 _5433_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5364_ _4443_/X hold438/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7466_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4878__A1 _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5724__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _7319_/Q _7335_/Q _7311_/Q _7447_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4315_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5443__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7103_ _5879_/A _7090_/X _7093_/X _7102_/Y vssd1 vssd1 vccd1 vccd1 _7103_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3970__A_N _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5295_ hold484/X _4964_/X _5301_/S vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__mux2_1
X_4246_ _7454_/Q _4242_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4246_/Y sky130_fd_sc_hd__a21oi_1
X_7034_ _5970_/A _6709_/S _7033_/Y _6989_/A vssd1 vssd1 vccd1 vccd1 _7034_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4774__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4177_ _4175_/X _4176_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4326__A_N _4325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5055__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4075__A _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6290__A _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6818_ _6851_/A _6784_/B _6817_/X vssd1 vssd1 vccd1 vccd1 _6838_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6749_ _6748_/X _6747_/Y split7/X _6669_/B vssd1 vssd1 vccd1 vccd1 _6773_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5294__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5046__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6794__B2 _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6794__A1 _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5080_ hold360/X _4849_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _7332_/D sky130_fd_sc_hd__mux2_1
X_4100_ _6075_/A _4942_/A vssd1 vssd1 vccd1 vccd1 _4993_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4594__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6375__A _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _5811_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__nand2_1
XANTENNA__7026__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5982_ _6374_/A _4119_/A _6013_/B _7169_/B _6020_/C vssd1 vssd1 vccd1 vccd1 _5982_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4796__A0 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4933_ _4933_/A _4933_/B vssd1 vssd1 vccd1 vccd1 _4933_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4864_ _3663_/Y _4964_/S _4860_/X _4863_/X vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__o22a_4
XANTENNA__4623__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3815_ _7477_/Q _7465_/Q _7457_/Q _7251_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3815_/X sky130_fd_sc_hd__mux4_1
X_4795_ hold472/X _4483_/X _4805_/S vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6603_ _6603_/A _6603_/B vssd1 vssd1 vccd1 vccd1 _6603_/X sky130_fd_sc_hd__xor2_1
X_7583_ _7590_/CLK _7583_/D vssd1 vssd1 vccd1 vccd1 _7583_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_59_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7590_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6534_ _6535_/A _6534_/B vssd1 vssd1 vccd1 vccd1 _6534_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout124_A _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3746_ _6216_/B _6216_/C vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6465_ _6742_/A _6467_/B _6461_/A vssd1 vssd1 vccd1 vccd1 _6466_/B sky130_fd_sc_hd__o21ba_1
X_3677_ input7/X vssd1 vssd1 vccd1 vccd1 _3677_/Y sky130_fd_sc_hd__inv_2
X_5416_ _7499_/Q _5415_/Y _6875_/A vssd1 vssd1 vccd1 vccd1 _5955_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6396_ _6962_/A _6383_/Y _6395_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6396_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5347_ hold510/X _4529_/X _5355_/S vssd1 vssd1 vccd1 vccd1 _5347_/X sky130_fd_sc_hd__mux2_1
X_5278_ hold429/X _4947_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _7424_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5276__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4229_ _4977_/A _4977_/B vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__nor2_1
X_7017_ input34/X _4021_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _7017_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7017__A2 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4533__A _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6528__A1 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4003__A2 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5751__A2 _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5811__B _5811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4146__C _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5975__C1 _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7192__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__B _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput22 custom_settings[29] vssd1 vssd1 vccd1 vccd1 _7631_/A sky130_fd_sc_hd__buf_2
XFILLER_0_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput11 custom_settings[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4580_ _4529_/S _4561_/X _4579_/Y _4541_/Y vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__a31o_4
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput44 rst_n vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
Xinput33 io_in[13] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6250_ _6962_/A _6869_/A vssd1 vssd1 vccd1 vccd1 _6279_/B sky130_fd_sc_hd__nor2_2
XANTENNA__5705__C _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5201_ hold257/X _4912_/Y _5211_/S vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__mux2_1
X_6181_ hold80/X hold44/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6181_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5132_ _5132_/A _5132_/B _6920_/D vssd1 vssd1 vccd1 vccd1 _6225_/B sky130_fd_sc_hd__or3_4
XANTENNA__5258__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5063_ hold377/X _4887_/X _5075_/S vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__mux2_1
X_4014_ _4007_/X _4012_/Y _7244_/A vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5449__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5965_ _5964_/A _5964_/B _5964_/C vssd1 vssd1 vccd1 vccd1 _5970_/C sky130_fd_sc_hd__o21a_1
X_4916_ _6057_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _4917_/B sky130_fd_sc_hd__nand2_1
X_5896_ _5923_/B _5896_/B vssd1 vssd1 vccd1 vccd1 _5898_/C sky130_fd_sc_hd__nor2_1
X_4847_ _7175_/B _5159_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5040_/S sky130_fd_sc_hd__and3_4
XANTENNA__7183__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5194__A0 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ hold263/X _4492_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7279_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7566_ _7577_/CLK _7566_/D vssd1 vssd1 vccd1 vccd1 _7566_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5733__A2 _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7497_ _7538_/CLK _7497_/D vssd1 vssd1 vccd1 vccd1 _7497_/Q sky130_fd_sc_hd__dfxtp_1
X_6517_ _6518_/A _6518_/B vssd1 vssd1 vccd1 vccd1 _6575_/A sky130_fd_sc_hd__or2_1
X_3729_ _6223_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _6022_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6448_ _6448_/A _6448_/B vssd1 vssd1 vccd1 vccd1 _6448_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6379_ hold58/X _3762_/B _3762_/D _4139_/Y vssd1 vssd1 vccd1 vccd1 _6379_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5631__B _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5123__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3830__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7475_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4160__A1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4438__A _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3996__B _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4173__A _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5750_ _6808_/A _5788_/B _6799_/A _6864_/A vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__and4_1
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4701_ _5008_/A _4701_/B _4701_/C _4701_/D vssd1 vssd1 vccd1 vccd1 _4701_/X sky130_fd_sc_hd__or4_1
XFILLER_0_17_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5681_ _5681_/A _5681_/B vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__and2_1
XANTENNA__7165__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7420_ _7454_/CLK _7420_/D vssd1 vssd1 vccd1 vccd1 _7420_/Q sky130_fd_sc_hd__dfxtp_1
X_4632_ _6157_/A _6148_/A _4632_/C vssd1 vssd1 vccd1 vccd1 _4682_/B sky130_fd_sc_hd__or3_1
X_4563_ _7480_/Q _7468_/Q _7460_/Q _7254_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4563_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5208__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7351_ _7427_/CLK _7351_/D vssd1 vssd1 vccd1 vccd1 _7351_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold603 _7550_/Q vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__buf_1
XANTENNA__3821__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7282_ _7597_/CLK _7282_/D vssd1 vssd1 vccd1 vccd1 _7282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4494_ _7602_/Q _4493_/C hold626/X vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__o21ai_1
Xhold636 _7542_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6302_ _6948_/B _6932_/C _6949_/A vssd1 vssd1 vccd1 vccd1 _6933_/B sky130_fd_sc_hd__a21bo_1
Xhold614 _6210_/X vssd1 vssd1 vccd1 vccd1 _7539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _7501_/Q vssd1 vssd1 vccd1 vccd1 _3683_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 _7550_/Q vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold658 _6793_/A vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _7556_/Q vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6298_/A _6827_/A vssd1 vssd1 vccd1 vccd1 _6233_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5732__A _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6025_/Y _6161_/Y _6163_/X vssd1 vssd1 vccd1 vccd1 _6164_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6428__B1 _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5115_ hold388/X _4864_/X _5129_/S vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout191_A _7360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6094_/X hold42/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__mux2_1
XANTENNA__6979__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5046_ hold597/X _4871_/Y _5058_/S vssd1 vssd1 vccd1 vccd1 _7317_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6979__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4782__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5403__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6997_ _6968_/A _6968_/B _6868_/Y vssd1 vssd1 vccd1 vccd1 _6998_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4083__A _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5948_ _5964_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5948_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7156__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5879_ _5879_/A _5879_/B vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7618_ _7618_/CLK _7618_/D vssd1 vssd1 vccd1 vccd1 _7618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5706__A2 _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7549_ _7579_/CLK _7549_/D vssd1 vssd1 vccd1 vccd1 _7549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5118__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4678__C1 _4144_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6738__A _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4692__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5158__A0 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5817__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5552__A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5330__A0 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6920_ _6920_/A _7599_/Q hold58/A _6920_/D vssd1 vssd1 vccd1 vccd1 _6920_/X sky130_fd_sc_hd__or4_1
X_6851_ _6851_/A _6882_/B vssd1 vssd1 vccd1 vccd1 _6884_/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ _5955_/A _5802_/B _5802_/C vssd1 vssd1 vccd1 vccd1 _5802_/X sky130_fd_sc_hd__and3_1
XANTENNA__4295__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3994_ _5990_/A _3985_/X _3989_/X _5804_/B _3993_/Y vssd1 vssd1 vccd1 vccd1 _3994_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6782_ _6782_/A _6790_/S _6782_/C vssd1 vssd1 vccd1 vccd1 _6782_/X sky130_fd_sc_hd__and3_1
XFILLER_0_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5733_ _6273_/A _6802_/B _5732_/C vssd1 vssd1 vccd1 vccd1 _5734_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__7138__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5664_ _5666_/D vssd1 vssd1 vccd1 vccd1 _5664_/Y sky130_fd_sc_hd__inv_2
X_7403_ _7403_/CLK _7403_/D vssd1 vssd1 vccd1 vccd1 _7403_/Q sky130_fd_sc_hd__dfxtp_1
X_4615_ _7481_/Q _7469_/Q _7461_/Q _7255_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4615_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6897__A0 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5595_ _5598_/B _5598_/C vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__and2_1
Xhold400 _5305_/X vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _5345_/X vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
X_7334_ _7446_/CLK _7334_/D vssd1 vssd1 vccd1 vccd1 _7334_/Q sky130_fd_sc_hd__dfxtp_1
X_4546_ _7376_/Q _7304_/Q _7296_/Q _7288_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4546_/X sky130_fd_sc_hd__mux4_1
Xhold422 _4386_/X vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _5187_/X vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _4630_/X vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold455 _7152_/X vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7153__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 _7596_/Q vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7265_ _7489_/CLK _7265_/D vssd1 vssd1 vccd1 vccd1 _7265_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4777__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold477 _5171_/X vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _4477_/A _4477_/B _4477_/C _4383_/A vssd1 vssd1 vccd1 vccd1 _4478_/B sky130_fd_sc_hd__or4b_1
Xhold499 _5244_/X vssd1 vssd1 vccd1 vccd1 _7409_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _5269_/X vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
X_7196_ hold205/X _4111_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7608_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6216_ _6216_/A _6216_/B _6216_/C vssd1 vssd1 vccd1 vccd1 _6216_/X sky130_fd_sc_hd__or3_1
XFILLER_0_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6147_ _3702_/Y _4600_/Y _6146_/X _6375_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6147_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _4238_/A _6080_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4427__A2 _4320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5624__A1 _6718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5401__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _6840_/A _4976_/B _5028_/X _5008_/A vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3710__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4060__A0 hold92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4260__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3797__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4210__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6040__A1 _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6040__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4051__A0 _7569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6142__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4400_ _7269_/Q _7609_/Q _7601_/Q _7617_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4400_/X sky130_fd_sc_hd__mux4_1
X_5380_ _5379_/X _4394_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7477_/D sky130_fd_sc_hd__mux2_1
X_4331_ _4474_/A _6044_/B vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__xor2_1
X_4262_ _4180_/Y _4261_/Y _4260_/X vssd1 vssd1 vccd1 vccd1 _4262_/X sky130_fd_sc_hd__o21a_1
Xfanout209 _6345_/A vssd1 vssd1 vccd1 vccd1 _6015_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7050_ _6244_/A _6926_/Y _7048_/X _7049_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7587_/D
+ sky130_fd_sc_hd__o221a_1
X_6001_ _3646_/Y hold80/X _3648_/Y hold64/X _6000_/X vssd1 vssd1 vccd1 vccd1 _6004_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4193_ _7318_/Q _7334_/Q _7310_/Q _7446_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4193_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5221__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6803__B1 _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6903_ _3949_/Y _6897_/X _6898_/X _6901_/Y _6902_/X vssd1 vssd1 vccd1 vccd1 _6905_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout154_A _7574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6834_ _6750_/Y _6755_/Y _6822_/A _6774_/Y vssd1 vssd1 vccd1 vccd1 _6834_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_107_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3977_ _7473_/Q hold56/X _6375_/A vssd1 vssd1 vccd1 vccd1 _3985_/C sky130_fd_sc_hd__o21a_1
X_6765_ _6750_/Y _6755_/Y _6760_/X _6764_/X vssd1 vssd1 vccd1 vccd1 _6765_/X sky130_fd_sc_hd__a211o_4
X_5716_ _5715_/B _5715_/C _5715_/A vssd1 vssd1 vccd1 vccd1 _5716_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6696_ _6869_/A _6697_/B vssd1 vssd1 vccd1 vccd1 _6698_/A sky130_fd_sc_hd__and2_1
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5647_ _5736_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__or2_1
XFILLER_0_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5578_ _5578_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5578_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold230 _7594_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
X_7317_ _7446_/CLK _7317_/D vssd1 vssd1 vccd1 vccd1 _7317_/Q sky130_fd_sc_hd__dfxtp_1
Xhold252 _7328_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _7298_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4495_/Y _4528_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4529_/X sky130_fd_sc_hd__mux2_8
Xhold285 _5298_/X vssd1 vssd1 vccd1 vccd1 _7433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _7406_/Q vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _4777_/X vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _7479_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
X_7248_ _4076_/X hold558/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7570_/D sky130_fd_sc_hd__mux2_1
X_7179_ hold649/X _4434_/Y _7191_/S vssd1 vssd1 vccd1 vccd1 _7179_/X sky130_fd_sc_hd__mux2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__A _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4271__A _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6198__A _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 custom_settings[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output48_A _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3900_ _4103_/A _3937_/A vssd1 vssd1 vccd1 vccd1 _3901_/B sky130_fd_sc_hd__nor2_1
X_4880_ _4875_/Y _5001_/A _4879_/X _4123_/A vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__o211a_1
X_3831_ _7321_/Q _7337_/Q _7313_/Q _7449_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3831_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6550_ _6529_/B _6558_/A _6504_/Y vssd1 vssd1 vccd1 vccd1 _6550_/Y sky130_fd_sc_hd__o21ai_1
X_3762_ _3762_/A _3762_/B _3762_/C _3762_/D vssd1 vssd1 vccd1 vccd1 _4724_/S sky130_fd_sc_hd__or4_2
XFILLER_0_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5501_ _5469_/Y _5495_/S _5500_/X vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5772__B1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3693_ _6204_/A _3693_/B vssd1 vssd1 vccd1 vccd1 _3693_/Y sky130_fd_sc_hd__nor2_1
X_6481_ _6476_/B _6480_/X _6481_/S vssd1 vssd1 vccd1 vccd1 _6484_/B sky130_fd_sc_hd__mux2_1
X_5432_ _5432_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5433_/B sky130_fd_sc_hd__nor2_1
X_5363_ hold437/X _4483_/X _5373_/S vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5216__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4314_ _4312_/X _4313_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7102_ _7102_/A _7102_/B _7102_/C _7102_/D vssd1 vssd1 vccd1 vccd1 _7102_/Y sky130_fd_sc_hd__nand4_1
X_5294_ _5293_/X _4921_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _7431_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4245_ _4243_/X _4244_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4245_/X sky130_fd_sc_hd__mux2_1
X_7033_ _7033_/A _7033_/B vssd1 vssd1 vccd1 vccd1 _7033_/Y sky130_fd_sc_hd__xnor2_1
X_4176_ _7268_/Q _7608_/Q _7600_/Q _7616_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4176_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4075__B _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6817_ _6841_/A _6817_/B _6817_/C vssd1 vssd1 vccd1 vccd1 _6817_/X sky130_fd_sc_hd__or3_1
XFILLER_0_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6748_ _6747_/A _6747_/B split7/X vssd1 vssd1 vccd1 vccd1 _6748_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679_ _6681_/B vssd1 vssd1 vccd1 vccd1 _6679_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5915__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5126__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4205__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6703__C1 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _5988_/A _4030_/B vssd1 vssd1 vccd1 vccd1 _4030_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5690__C1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5981_ _7230_/A _3962_/D _5980_/B _4034_/B _6374_/A vssd1 vssd1 vccd1 vccd1 _6020_/C
+ sky130_fd_sc_hd__o2111a_1
X_4932_ _5031_/S _4930_/X _4931_/Y _4963_/S vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4863_ _4963_/S _4861_/X _4862_/Y _4989_/A vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__a31o_1
X_6602_ _6651_/A _6651_/B _6544_/Y _6548_/Y vssd1 vssd1 vccd1 vccd1 split9/A sky130_fd_sc_hd__a211o_4
X_3814_ _3931_/S _3814_/B vssd1 vssd1 vccd1 vccd1 _3814_/Y sky130_fd_sc_hd__nand2_1
X_4794_ _4394_/X _4793_/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7285_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7582_ _7582_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6533_ _6545_/A _6545_/B _6490_/X vssd1 vssd1 vccd1 vccd1 _6534_/B sky130_fd_sc_hd__a21o_1
X_3745_ _3741_/X _6357_/A _5990_/A vssd1 vssd1 vccd1 vccd1 _3762_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6464_ _6742_/A _6467_/B vssd1 vssd1 vccd1 vccd1 _6506_/A sky130_fd_sc_hd__nor2_1
X_5415_ hold78/A _6802_/B vssd1 vssd1 vccd1 vccd1 _5415_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _6827_/A vssd1 vssd1 vccd1 vccd1 _6840_/A sky130_fd_sc_hd__inv_6
XANTENNA_fanout117_A _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7618_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6395_ hold124/X _6415_/A _6356_/B hold92/X vssd1 vssd1 vccd1 vccd1 _6395_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4720__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5346_ _4443_/X hold411/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7458_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4785__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5277_ hold428/X _4964_/X _5283_/S vssd1 vssd1 vccd1 vccd1 _5277_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6566__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7161__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3906__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4228_ _4977_/B vssd1 vssd1 vccd1 vccd1 _4228_/Y sky130_fd_sc_hd__inv_2
X_7016_ _6996_/X _7015_/Y _4723_/A vssd1 vssd1 vccd1 vccd1 _7016_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4159_ _7527_/Q _4162_/B vssd1 vssd1 vccd1 vccd1 _4159_/X sky130_fd_sc_hd__or2_1
XANTENNA__4236__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6476__A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4778__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5975__B1 _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4162__C _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 custom_settings[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
XANTENNA__4950__A1 _4955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6150__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 io_in[14] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
Xinput23 custom_settings[2] vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5200_ _4871_/Y hold538/X _5212_/S vssd1 vssd1 vccd1 vccd1 _7389_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6180_ _3751_/Y _6178_/X _6179_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6180_/X sky130_fd_sc_hd__o211a_1
X_5131_ _5132_/A _5132_/B _6920_/D vssd1 vssd1 vccd1 vccd1 _6229_/S sky130_fd_sc_hd__nor3_2
X_5062_ hold556/X _4849_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _7324_/D sky130_fd_sc_hd__mux2_1
X_4013_ _5952_/A _4267_/D vssd1 vssd1 vccd1 vccd1 _4013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4313__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5964_ _5964_/A _5964_/B _5964_/C vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4915_ _6057_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _4915_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5895_ _6516_/A _6702_/A _5894_/C vssd1 vssd1 vccd1 vccd1 _5896_/B sky130_fd_sc_hd__a21oi_1
X_4846_ _4846_/A _4945_/B _4846_/C vssd1 vssd1 vccd1 vccd1 _5303_/C sky130_fd_sc_hd__nand3_4
XFILLER_0_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7565_ _7577_/CLK _7565_/D vssd1 vssd1 vccd1 vccd1 _7565_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6391__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7156__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4777_ hold262/X _4529_/X _4785_/S vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6060__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5465__A _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6516_ _6516_/A _6516_/B vssd1 vssd1 vccd1 vccd1 _6518_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7496_ _7498_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
X_3728_ _3728_/A _7230_/B vssd1 vssd1 vccd1 vccd1 _6383_/A sky130_fd_sc_hd__and2_4
XFILLER_0_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3659_ hold82/A vssd1 vssd1 vccd1 vccd1 _3659_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6447_ _5615_/B _6451_/B _5597_/X vssd1 vssd1 vccd1 vccd1 _6448_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6378_ _5980_/Y _6377_/X _6416_/A vssd1 vssd1 vccd1 vccd1 _6378_/Y sky130_fd_sc_hd__o21ai_1
X_5329_ hold605/X _4937_/Y _5337_/S vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5404__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3713__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__C _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5078__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6906__C1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5185__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6382__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4932__A1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4696__B1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4543__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _6827_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4701_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5680_ _5681_/A _5681_/B vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__nor2_2
X_4631_ _4589_/X hold433/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7255_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5176__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4562_ _7280_/Q _7595_/Q _7264_/Q _7488_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4562_/X sky130_fd_sc_hd__mux4_1
X_7350_ _7427_/CLK _7350_/D vssd1 vssd1 vccd1 vccd1 _7350_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4384__C1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7281_ _7593_/CLK _7281_/D vssd1 vssd1 vccd1 vccd1 _7281_/Q sky130_fd_sc_hd__dfxtp_1
Xhold626 _7603_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _7602_/Q _7603_/Q _4493_/C vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__or3_1
Xhold604 _4058_/X vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6301_ _6301_/A _6909_/B vssd1 vssd1 vccd1 vccd1 _6932_/C sky130_fd_sc_hd__nand2_1
Xhold615 _7559_/Q vssd1 vssd1 vccd1 vccd1 _3744_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold659 _6402_/X vssd1 vssd1 vccd1 vccd1 _7576_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold637 _6872_/B vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _7244_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _7556_/D sky130_fd_sc_hd__nor2_1
Xhold648 _6231_/X vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5732__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5224__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _7607_/Q _6162_/A _6162_/Y _3975_/X vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__a211o_1
X_5114_ _7212_/C _7194_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5129_/S sky130_fd_sc_hd__and3_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6427_/B _6092_/X _6093_/Y _4248_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6094_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5045_ hold596/X _4887_/X _5057_/S vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5100__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6844__A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout184_A _7452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6996_ _6990_/X _6992_/Y _6995_/X _6220_/C vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5947_ _5947_/A _5947_/B vssd1 vssd1 vccd1 vccd1 _5948_/B sky130_fd_sc_hd__and2_1
XFILLER_0_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7617_ _7617_/CLK _7617_/D vssd1 vssd1 vccd1 vccd1 _7617_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5167__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6364__A0 hold92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5878_ _5877_/A _5877_/B _5877_/C vssd1 vssd1 vccd1 vccd1 _5879_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4829_ hold578/X _4385_/X _4843_/S vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7306_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3708__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4303__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4914__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7548_ _7579_/CLK _7548_/D vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_2
X_7479_ _7479_/CLK _7479_/D vssd1 vssd1 vccd1 vccd1 _7479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6738__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6754__A _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5817__B _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7006__A2_N _7040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4516__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4883__S _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7083__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6850_ _6793_/B _6891_/B _6849_/X vssd1 vssd1 vccd1 vccd1 _6882_/B sky130_fd_sc_hd__o21a_1
XANTENNA__5397__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6781_ _6781_/A _6781_/B _6781_/C vssd1 vssd1 vccd1 vccd1 _6782_/C sky130_fd_sc_hd__nand3_1
X_5801_ _5800_/B _5800_/C _5800_/A vssd1 vssd1 vccd1 vccd1 _5802_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3993_ _4122_/D _4065_/C vssd1 vssd1 vccd1 vccd1 _3993_/Y sky130_fd_sc_hd__nor2_1
X_5732_ _6273_/A _6802_/B _5732_/C vssd1 vssd1 vccd1 vccd1 _5763_/B sky130_fd_sc_hd__and3_1
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7138__A2 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5149__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5219__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5663_ _6683_/A _6637_/A _6793_/A _6690_/A vssd1 vssd1 vccd1 vccd1 _5666_/D sky130_fd_sc_hd__a22o_1
X_7402_ _7434_/CLK _7402_/D vssd1 vssd1 vccd1 vccd1 _7402_/Q sky130_fd_sc_hd__dfxtp_1
X_4614_ _7281_/Q _7596_/Q _7265_/Q _7489_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4614_/X sky130_fd_sc_hd__mux4_1
X_5594_ _5594_/A _5605_/B _5594_/C vssd1 vssd1 vccd1 vccd1 _5598_/C sky130_fd_sc_hd__nand3_2
Xhold401 _5306_/X vssd1 vssd1 vccd1 vccd1 _7436_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4545_ _4689_/A _4545_/B vssd1 vssd1 vccd1 vccd1 _4545_/X sky130_fd_sc_hd__and2_1
X_7333_ _7446_/CLK _7333_/D vssd1 vssd1 vccd1 vccd1 _7333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold434 _7254_/Q vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _7272_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _7314_/Q vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _7326_/Q vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7264_ _7483_/CLK _7264_/D vssd1 vssd1 vccd1 vccd1 _7264_/Q sky130_fd_sc_hd__dfxtp_1
Xhold467 _7162_/X vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _7397_/Q vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _6098_/B _6107_/B _4474_/A vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__a21o_1
Xhold456 _7291_/Q vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold489 _7374_/Q vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
X_7195_ hold204/X _4385_/X _7209_/S vssd1 vssd1 vccd1 vccd1 _7195_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6215_ hold52/X _3754_/B _6214_/Y vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__a21o_1
X_6146_ _6025_/Y _6143_/Y _6145_/X vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__o21a_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__B _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6076_/X hold38/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__mux2_1
X_5028_ _5001_/A _5023_/X _5027_/Y _4957_/X _5025_/X vssd1 vssd1 vccd1 vccd1 _5028_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4094__A _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3710__B _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5388__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold144_A _7525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6979_ _6989_/A _7009_/C _6978_/Y _6977_/Y _5879_/A vssd1 vssd1 vccd1 vccd1 _6979_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5129__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4899__B1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3797__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5312__A1 _4921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3901__A _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6484__A _6840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5379__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4051__A1 _6882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5039__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4360_/B _4329_/X _4326_/Y vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__o21ai_2
X_4261_ _5027_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6000_ _3644_/Y hold88/X _3648_/A _3649_/Y vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__a22o_1
X_4192_ _4688_/S _4192_/B vssd1 vssd1 vccd1 vccd1 _4192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6902_ _6872_/A _6911_/A _7098_/A _7078_/A _6899_/Y vssd1 vssd1 vccd1 vccd1 _6902_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6833_ _6773_/B _6832_/A _6831_/X _6832_/Y vssd1 vssd1 vccd1 vccd1 _6836_/C sky130_fd_sc_hd__o22a_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6031__A2 _6022_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3976_ _4084_/A _5811_/A vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_A _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6764_ _6764_/A _6764_/B _6764_/C _6763_/Y vssd1 vssd1 vccd1 vccd1 _6764_/X sky130_fd_sc_hd__or4b_4
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6695_ _6625_/B _6694_/X _6709_/S vssd1 vssd1 vccd1 vccd1 _6697_/B sky130_fd_sc_hd__mux2_4
X_5715_ _5715_/A _5715_/B _5715_/C vssd1 vssd1 vccd1 vccd1 _5814_/B sky130_fd_sc_hd__or3_2
XFILLER_0_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5646_ _5681_/A _5646_/B vssd1 vssd1 vccd1 vccd1 _5653_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7164__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 _7199_/X vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_5577_ _5577_/A _5577_/B vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold242 _7597_/Q vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _7158_/X vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _5069_/X vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
X_7316_ _7423_/CLK _7316_/D vssd1 vssd1 vccd1 vccd1 _7316_/Q sky130_fd_sc_hd__dfxtp_1
X_4528_ _4515_/X _4527_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__mux2_1
Xhold275 _5237_/X vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _7260_/Q vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _7413_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
X_7247_ _4073_/X hold524/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7569_/D sky130_fd_sc_hd__mux2_1
X_4459_ _6799_/A _4458_/X _4700_/B vssd1 vssd1 vccd1 vccd1 _4459_/X sky130_fd_sc_hd__mux2_1
Xhold297 _5383_/X vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_7178_ _7177_/X _4111_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7600_/D sky130_fd_sc_hd__mux2_1
XANTENNA__7047__A1 _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6129_ _5810_/A _6123_/B _6128_/Y _4122_/C _6027_/Y vssd1 vssd1 vccd1 vccd1 _6129_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3721__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5648__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4552__A _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3920__A1_N _3665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3631__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _7401_/Q _7393_/Q _7369_/Q _7385_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3830_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7210__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5772__A1 _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3761_ _6345_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3762_/D sky130_fd_sc_hd__nand2_1
X_5500_ split8/A _5500_/B _5500_/C vssd1 vssd1 vccd1 vccd1 _5500_/X sky130_fd_sc_hd__or3_4
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5772__B2 _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3692_ _4084_/A _5952_/A _4723_/A vssd1 vssd1 vccd1 vccd1 _3693_/B sky130_fd_sc_hd__a21oi_1
X_6480_ _6480_/A _6480_/B vssd1 vssd1 vccd1 vccd1 _6480_/X sky130_fd_sc_hd__xor2_1
X_5431_ _5438_/A _5438_/B _5438_/C vssd1 vssd1 vccd1 vccd1 _5434_/S sky130_fd_sc_hd__or3_4
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3806__A _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5362_ _4394_/X _5361_/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7465_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4401__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5724__C _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4313_ _7399_/Q _7391_/Q _7367_/Q _7383_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4313_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7101_ _7101_/A _7101_/B _7101_/C vssd1 vssd1 vccd1 vccd1 _7102_/D sky130_fd_sc_hd__or3_1
X_5293_ hold442/X _4937_/Y _5301_/S vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__mux2_1
X_7032_ _6900_/A _7019_/A _7029_/X _7031_/Y _3949_/Y vssd1 vssd1 vccd1 vccd1 _7032_/X
+ sky130_fd_sc_hd__o221a_1
X_4244_ _7427_/Q _7359_/Q _7351_/Q _7331_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4244_/X sky130_fd_sc_hd__mux4_1
X_4175_ _7372_/Q _7300_/Q _7292_/Q _7284_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4175_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4637__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6852__A _6882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7159__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5212__A0 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7201__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6816_ _6817_/B _6817_/C vssd1 vssd1 vccd1 vccd1 _6841_/B sky130_fd_sc_hd__nor2_1
X_6747_ _6747_/A _6747_/B vssd1 vssd1 vccd1 vccd1 _6747_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _5977_/B _7554_/Q _7553_/Q _5988_/A vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__and4_1
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6678_ _6709_/S _6676_/Y _6677_/X vssd1 vssd1 vccd1 vccd1 _6681_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5629_ _5631_/D vssd1 vssd1 vccd1 vccd1 _5629_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5915__B _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5407__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6123__A_N _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5754__A1 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3860__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5825__B _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output60_A _7542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5052__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6219__C1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5690__B1 _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5442__B1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6672__A _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_split32_A _5556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5980_ _6374_/A _5980_/B vssd1 vssd1 vccd1 vccd1 _5980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A _5031_/S vssd1 vssd1 vccd1 vccd1 _4931_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4192__A _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4862_ _4862_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _4862_/Y sky130_fd_sc_hd__nand2_1
X_3813_ _7277_/Q _7592_/Q _7261_/Q _7485_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3814_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6601_ _6601_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _6601_/Y sky130_fd_sc_hd__nand2_1
X_4793_ hold328/X _4434_/Y _4805_/S vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3812__A1_N _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7581_ _7581_/CLK _7581_/D vssd1 vssd1 vccd1 vccd1 _7581_/Q sky130_fd_sc_hd__dfxtp_2
X_6532_ _6532_/A _6532_/B vssd1 vssd1 vccd1 vccd1 _6545_/B sky130_fd_sc_hd__xnor2_1
X_3744_ _3744_/A _6015_/C vssd1 vssd1 vccd1 vccd1 _6357_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3675_ _6532_/A vssd1 vssd1 vccd1 vccd1 _6754_/A sky130_fd_sc_hd__inv_2
X_6463_ _5601_/X _6462_/X _6463_/S vssd1 vssd1 vccd1 vccd1 _6467_/B sky130_fd_sc_hd__mux2_4
XANTENNA__5227__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5414_ _6683_/B _6518_/A _5818_/B _5438_/A _7499_/Q vssd1 vssd1 vccd1 vccd1 _5417_/B
+ sky130_fd_sc_hd__o41ai_2
XFILLER_0_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6394_ _6393_/X hold660/X _6414_/S vssd1 vssd1 vccd1 vccd1 _7574_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5345_ hold410/X _4483_/X _5355_/S vssd1 vssd1 vccd1 vccd1 _5345_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5276_ _5275_/X _4921_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _7423_/D sky130_fd_sc_hd__mux2_1
X_4227_ _4689_/A _4225_/X _4226_/Y _4221_/Y vssd1 vssd1 vccd1 vccd1 _4977_/B sky130_fd_sc_hd__a2bb2o_2
XANTENNA__3906__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7015_ _4030_/B _7013_/X _7014_/X vssd1 vssd1 vccd1 vccd1 _7015_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__4484__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4086__B _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4158_ hold66/A input13/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4236__A1 _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4089_ _4747_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _5357_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 custom_settings[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XANTENNA__4935__C1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 io_in[15] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_2
Xinput24 custom_settings[3] vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__buf_1
XANTENNA__5047__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6688__C1 _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5130_ hold569/X _5022_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _7359_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ hold555/X _4864_/X _5075_/S vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4012_ _5977_/B _4007_/B _4010_/Y _3733_/B vssd1 vssd1 vccd1 vccd1 _4012_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5663__B1 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4915__A _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4313__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5966__A1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5963_ _5970_/B _5963_/B vssd1 vssd1 vccd1 vccd1 _5964_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4914_ _4913_/X _4897_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _7310_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3977__B1 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _6516_/A _6702_/A _5894_/C vssd1 vssd1 vccd1 vccd1 _5923_/B sky130_fd_sc_hd__and3_1
X_4845_ _4846_/A _4945_/B _4846_/C vssd1 vssd1 vccd1 vccd1 _5321_/B sky130_fd_sc_hd__and3_2
XFILLER_0_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4776_ hold226/X _4443_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7278_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7564_ _7577_/CLK _7564_/D vssd1 vssd1 vccd1 vccd1 _7564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3824__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3727_ _6225_/A _5988_/A _3960_/C vssd1 vssd1 vccd1 vccd1 _7230_/B sky130_fd_sc_hd__or3_4
XANTENNA__6391__B2 hold558/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6515_ _6521_/A _6521_/D _6683_/B vssd1 vssd1 vccd1 vccd1 _6516_/B sky130_fd_sc_hd__a21oi_1
X_7495_ _7498_/CLK hold87/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4154__A0 _7569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ _7494_/Q vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__inv_2
XFILLER_0_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6446_ _6474_/A _6446_/B vssd1 vssd1 vccd1 vccd1 _6485_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4796__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6377_ _3716_/B _3780_/B _6383_/B vssd1 vssd1 vccd1 vccd1 _6377_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5328_ _4897_/X _5327_/X _5338_/S vssd1 vssd1 vccd1 vccd1 _5328_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3713__B hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5259_ hold318/X _4964_/X _5265_/S vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4457__A1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold174_A _7520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5406__A0 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5656__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3815__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6382__B2 hold66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4240__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__A1 _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4543__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout190 _3896_/S0 vssd1 vssd1 vccd1 vccd1 _3883_/S0 sky130_fd_sc_hd__buf_8
XANTENNA__5330__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4454__B _4460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4481__A1_N _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4630_ hold432/X _4629_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5566__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5285__B _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4561_ _5031_/S _4557_/X _4559_/X _4560_/X vssd1 vssd1 vccd1 vccd1 _4561_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6300_ _6311_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _6948_/B sky130_fd_sc_hd__nand2_2
X_7280_ _7598_/CLK _7280_/D vssd1 vssd1 vccd1 vccd1 _7280_/Q sky130_fd_sc_hd__dfxtp_1
Xhold605 _7447_/Q vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 _7183_/X vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _5022_/A _4492_/B vssd1 vssd1 vccd1 vccd1 _4492_/X sky130_fd_sc_hd__or2_4
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold616 _6352_/X vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold649 _7601_/Q vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _6386_/X vssd1 vssd1 vccd1 vccd1 _7572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ hold647/X _5994_/D _5988_/X _6220_/B vssd1 vssd1 vccd1 vccd1 _6231_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4231__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3814__A _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6162_/A _6162_/B vssd1 vssd1 vccd1 vccd1 _6162_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5113_ _7211_/C _7193_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5130_/S sky130_fd_sc_hd__and3_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6093_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6093_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5044_ hold321/X _4849_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _7316_/D sky130_fd_sc_hd__mux2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5240__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6995_ _3716_/Y _6988_/Y _6993_/Y _6994_/X vssd1 vssd1 vccd1 vccd1 _6995_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5946_ _5947_/A _5947_/B vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__nor2_1
X_5877_ _5877_/A _5877_/B _5877_/C vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__and3_1
XANTENNA__7167__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4828_ _7212_/B _5322_/B _7194_/C vssd1 vssd1 vccd1 vccd1 _4843_/S sky130_fd_sc_hd__and3_4
X_7616_ _7617_/CLK _7616_/D vssd1 vssd1 vccd1 vccd1 _7616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4470__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4759_ hold469/X _4529_/X _4767_/S vssd1 vssd1 vccd1 vccd1 _4759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7547_ _7547_/CLK _7547_/D vssd1 vssd1 vccd1 vccd1 _7547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7478_ _7596_/CLK _7478_/D vssd1 vssd1 vccd1 vccd1 _7478_/Q sky130_fd_sc_hd__dfxtp_1
X_6429_ _6223_/A _4103_/A _4030_/B vssd1 vssd1 vccd1 vccd1 _6429_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4222__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4004_/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4678__A1 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5150__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5817__C _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4213__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5325__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3634__A _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7068__C1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4516__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7083__A2 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5094__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4841__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3992_ _7553_/Q _6223_/A _3992_/C vssd1 vssd1 vccd1 vccd1 _4065_/C sky130_fd_sc_hd__or3_2
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6680__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6780_ _6844_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6780_/X sky130_fd_sc_hd__or2_1
X_5800_ _5800_/A _5800_/B _5800_/C vssd1 vssd1 vccd1 vccd1 _5802_/B sky130_fd_sc_hd__or3_1
X_5731_ _5763_/A _5731_/B vssd1 vssd1 vccd1 vccd1 _5732_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5662_ _5662_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__nor2_1
XANTENNA__6346__A1 _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6346__B2 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7401_ _7449_/CLK _7401_/D vssd1 vssd1 vccd1 vccd1 _7401_/Q sky130_fd_sc_hd__dfxtp_1
X_4613_ _4982_/A _4611_/X _4612_/X _4162_/B vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__o211a_1
X_5593_ _5605_/B _5594_/C _5594_/A vssd1 vssd1 vccd1 vccd1 _5598_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_4_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold402 _7391_/Q vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
X_4544_ _4542_/X _4543_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__mux2_1
X_7332_ _7448_/CLK _7332_/D vssd1 vssd1 vccd1 vccd1 _7332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold435 _7489_/Q vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
X_7263_ _7487_/CLK _7263_/D vssd1 vssd1 vccd1 vccd1 _7263_/Q sky130_fd_sc_hd__dfxtp_1
Xhold424 _5016_/X vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _5066_/X vssd1 vssd1 vccd1 vccd1 _7326_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold457 _7261_/Q vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _7462_/Q vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4204__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 _7426_/Q vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4475_/A _4525_/A vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__nand2_1
X_6214_ _6345_/A _6920_/D vssd1 vssd1 vccd1 vccd1 _6214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold479 _5217_/X vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_7194_ _7212_/B _7212_/C _7194_/C vssd1 vssd1 vccd1 vccd1 _7209_/S sky130_fd_sc_hd__and3_4
XFILLER_0_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6145_ _7605_/Q _6153_/A _6144_/Y _3975_/X vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__a211o_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6427_/B _6074_/X _6075_/Y _4228_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6076_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__C1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5085__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5027_ _5027_/A _5027_/B vssd1 vssd1 vccd1 vccd1 _5027_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4832__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4094__B _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6978_ _6978_/A _6978_/B _6978_/C vssd1 vssd1 vccd1 vccd1 _6978_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__4691__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5929_ _5930_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3719__A _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4314__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6337__A1 _7040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5145__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4269__B _4879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4823__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4587__B1 _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6931__C _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5000__A1 _4238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5055__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4260_ _4407_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4191_ _7398_/Q _7390_/Q _7366_/Q _7382_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4192_/B sky130_fd_sc_hd__mux4_1
XANTENNA__5067__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4814__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4275__C1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6901_ _7070_/A _7095_/A _6948_/B vssd1 vssd1 vccd1 vccd1 _6901_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6832_ _6832_/A _6832_/B vssd1 vssd1 vccd1 vccd1 _6832_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6016__B1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6763_ _6653_/Y _6763_/B vssd1 vssd1 vccd1 vccd1 _6763_/Y sky130_fd_sc_hd__nand2b_1
X_3975_ _6220_/C _4140_/B vssd1 vssd1 vccd1 vccd1 _3975_/X sky130_fd_sc_hd__or2_4
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6694_ _6694_/A _6694_/B vssd1 vssd1 vccd1 vccd1 _6694_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_18_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5714_ _5714_/A _5714_/B _5714_/C vssd1 vssd1 vccd1 vccd1 _5715_/C sky130_fd_sc_hd__and3_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5645_ _5644_/A _5675_/A _5640_/Y vssd1 vssd1 vccd1 vccd1 _5646_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 _7356_/Q vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5473__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5576_ _6793_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _6442_/A sky130_fd_sc_hd__xnor2_2
Xhold232 _7442_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _7301_/Q vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
X_7315_ _7451_/CLK _7315_/D vssd1 vssd1 vccd1 vccd1 _7315_/Q sky130_fd_sc_hd__dfxtp_1
X_4527_ _4487_/A _4526_/Y _4986_/S vssd1 vssd1 vccd1 vccd1 _4527_/X sky130_fd_sc_hd__mux2_1
Xhold243 _7533_/Q vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _5238_/X vssd1 vssd1 vccd1 vccd1 _7406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _4731_/X vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _5253_/X vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
X_7246_ hold99/X hold66/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7246_/X sky130_fd_sc_hd__mux2_1
X_4458_ _4455_/X _4457_/X _4701_/B vssd1 vssd1 vccd1 vccd1 _4458_/X sky130_fd_sc_hd__mux2_1
Xhold254 _7530_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__buf_1
Xhold298 _7335_/Q vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_7177_ _4170_/A _4385_/X _7191_/S vssd1 vssd1 vccd1 vccd1 _7177_/X sky130_fd_sc_hd__mux2_1
X_6128_ _6025_/Y _6125_/Y _6127_/X vssd1 vssd1 vccd1 vccd1 _6128_/Y sky130_fd_sc_hd__o21ai_2
X_4389_ _6111_/A _4389_/B vssd1 vssd1 vccd1 vccd1 _4390_/C sky130_fd_sc_hd__nand2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4805__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6059_ _6058_/X hold46/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__mux2_1
XFILLER_0_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5230__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4664__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5648__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4416__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5297__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3912__A _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4257__C1 _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5221__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _6216_/B _3758_/Y _6211_/B _5132_/B _3749_/Y vssd1 vssd1 vccd1 vccd1 _3761_/B
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4889__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5772__A2 _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5430_ _5428_/B _5428_/C _6871_/A vssd1 vssd1 vccd1 vccd1 _5438_/C sky130_fd_sc_hd__a21oi_4
XFILLER_0_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3691_ _6223_/A _5808_/A vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ hold571/X _4434_/Y _5373_/S vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5724__D _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5292_ hold269/X _4897_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__mux2_1
X_4312_ _7439_/Q _7431_/Q _7415_/Q _7407_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4312_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7100_ _7109_/A _7109_/B _7100_/C vssd1 vssd1 vccd1 vccd1 _7101_/C sky130_fd_sc_hd__and3_1
XANTENNA__5288__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4243_ _7323_/Q _7339_/Q _7315_/Q _7451_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4243_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7031_ split4/X _7030_/Y _6900_/A vssd1 vssd1 vccd1 vccd1 _7031_/Y sky130_fd_sc_hd__o21ai_1
X_4174_ _7476_/Q _7464_/Q _7456_/Q _7250_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4174_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6815_ _6817_/B _6815_/B vssd1 vssd1 vccd1 vccd1 _6848_/C sky130_fd_sc_hd__or2_1
XFILLER_0_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4646__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6746_ _6751_/A _6751_/B _6674_/A vssd1 vssd1 vccd1 vccd1 _6747_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4799__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3958_ _7098_/A _7230_/C _3973_/B _6920_/A vssd1 vssd1 vccd1 vccd1 _4113_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3889_ _6084_/A vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__inv_2
XFILLER_0_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6677_ _6629_/B _6629_/C _6670_/A _6648_/X _6658_/X vssd1 vssd1 vccd1 vccd1 _6677_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5628_ _6802_/A _6637_/A _6702_/A _6808_/A vssd1 vssd1 vccd1 vccd1 _5631_/D sky130_fd_sc_hd__a22o_1
X_5559_ _6532_/A _5566_/B _5558_/X vssd1 vssd1 vccd1 vccd1 _5559_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__5279__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4828__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7229_ _6417_/B _3728_/A _6015_/B _4033_/X _6015_/A vssd1 vssd1 vccd1 vccd1 _7231_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_hold636_A _7542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5203__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__C1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5754__A2 _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3860__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4502__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6703__A1 _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5825__C _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5911__C1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5333__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3642__A hold97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output53_A _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4473__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _4926_/X _4929_/X _4930_/S vssd1 vssd1 vccd1 vccd1 _4930_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7195__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4861_ _5034_/B _4861_/B vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3812_ _7363_/Q _3810_/X _3811_/Y _3806_/Y vssd1 vssd1 vccd1 vccd1 _6139_/A sky130_fd_sc_hd__a2bb2o_4
X_6600_ _6600_/A _6600_/B vssd1 vssd1 vccd1 vccd1 _6651_/B sky130_fd_sc_hd__and2_1
X_4792_ _4111_/X hold426/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7284_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6942__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7580_ _7582_/CLK _7580_/D vssd1 vssd1 vccd1 vccd1 _7580_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6531_ _6531_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _6545_/A sky130_fd_sc_hd__nand2_1
X_3743_ _6922_/A _3763_/A vssd1 vssd1 vccd1 vccd1 _6015_/C sky130_fd_sc_hd__nand2_2
X_3674_ _6611_/A vssd1 vssd1 vccd1 vccd1 _6673_/A sky130_fd_sc_hd__inv_4
X_6462_ _6462_/A _6462_/B vssd1 vssd1 vccd1 vccd1 _6462_/X sky130_fd_sc_hd__xor2_1
X_5413_ _3656_/Y _6802_/B _5788_/D _5818_/B _5438_/A vssd1 vssd1 vccd1 vccd1 _5413_/X
+ sky130_fd_sc_hd__a2111o_1
X_6393_ input33/X _6392_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__mux2_1
X_5344_ _4394_/X _5343_/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7457_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6458__B1 _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5275_ hold462/X _4937_/Y _5283_/S vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _4688_/S _4222_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4226_/Y sky130_fd_sc_hd__a21oi_1
X_7014_ _6057_/A _5804_/C _4029_/Y _6130_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _7014_/X
+ sky130_fd_sc_hd__a221o_1
X_4157_ _4751_/A vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__inv_2
XANTENNA__4086__C _4846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3692__B1 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4088_ hold669/X input10/X _5022_/A vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5479__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7483_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7186__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6729_ _6729_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6729_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5153__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4992__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5672__A1 _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A0 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7177__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5328__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 custom_settings[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XANTENNA__3637__A _7558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput36 io_in[16] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_2
Xinput25 custom_settings[4] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5360__A0 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5063__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6159__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ _7212_/A _7212_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5075_/S sky130_fd_sc_hd__and3_4
XFILLER_0_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5663__B2 _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__A1 _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4011_ _4033_/B _6331_/B vssd1 vssd1 vccd1 vccd1 _4011_/X sky130_fd_sc_hd__or2_1
XANTENNA__6683__A _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5962_ _5961_/A _5961_/B _5961_/C vssd1 vssd1 vccd1 vccd1 _5963_/B sky130_fd_sc_hd__a21oi_1
X_4913_ hold331/X _4912_/Y _5039_/S vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__mux2_1
X_5893_ _5923_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5894_/C sky130_fd_sc_hd__nor2_1
X_4844_ _4843_/X _4685_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7307_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4931__A _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6915__A1 _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6376__C1 _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4775_ hold225/X _4483_/X _4785_/S vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4650__B _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7563_ _7577_/CLK _7563_/D vssd1 vssd1 vccd1 vccd1 _7563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5238__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3824__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3726_ _7553_/Q _6223_/A _3960_/C vssd1 vssd1 vccd1 vccd1 _3728_/A sky130_fd_sc_hd__or3_4
X_6514_ _6512_/Y _6514_/B vssd1 vssd1 vccd1 vccd1 _6563_/A sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout122_A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7494_ _7498_/CLK _7494_/D vssd1 vssd1 vccd1 vccd1 _7494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3657_ hold90/A vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__inv_2
XFILLER_0_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6445_ _6445_/A _6487_/B vssd1 vssd1 vccd1 vccd1 _6446_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6376_ _5990_/A _6375_/X _6229_/S _6207_/S _3757_/A vssd1 vssd1 vccd1 vccd1 _6927_/A
+ sky130_fd_sc_hd__a2111o_2
X_5327_ hold451/X _4912_/Y _5337_/S vssd1 vssd1 vccd1 vccd1 _5327_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6069__S _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5481__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _5257_/X _4921_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _7415_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ hold520/X _4990_/Y _5193_/S vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__mux2_1
X_4209_ _4209_/A _4209_/B vssd1 vssd1 vccd1 vccd1 _4955_/A sky130_fd_sc_hd__and2_2
XFILLER_0_97_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4317__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3968__A1 _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7159__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4090__A0 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6906__A1 _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5656__B _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3815__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5148__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6119__C1 _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4052__S _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5342__A0 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3888__A1_N _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4145__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4240__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__A2 _4694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout180 _7453_/Q vssd1 vssd1 vccd1 vccd1 _4686_/S1 sky130_fd_sc_hd__buf_6
Xfanout191 _7360_/Q vssd1 vssd1 vccd1 vccd1 _3896_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4751__A _4751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5058__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4384__A1 _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4560_ input4/X _4850_/A _4700_/B _4963_/S vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4491_ _4083_/X _4489_/X _4490_/X _4536_/B vssd1 vssd1 vccd1 vccd1 _4492_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold617 _6353_/X vssd1 vssd1 vccd1 vccd1 _7559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold606 _7473_/Q vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold639 _7347_/Q vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _7184_/X vssd1 vssd1 vccd1 vccd1 _7603_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6230_ _7244_/A _6230_/B vssd1 vssd1 vccd1 vccd1 _7555_/D sky130_fd_sc_hd__or2_1
XANTENNA__4231__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6161_ _6161_/A vssd1 vssd1 vccd1 vccd1 _6161_/Y sky130_fd_sc_hd__inv_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5884__A1 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5112_ _5111_/X _5022_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _7351_/D sky130_fd_sc_hd__mux2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6328_/A _4248_/Y _6091_/X _6375_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6092_/X
+ sky130_fd_sc_hd__o221a_1
X_5043_ hold320/X _4864_/X _5057_/S vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__mux2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6994_ _7009_/B _6993_/B _6913_/A vssd1 vssd1 vccd1 vccd1 _6994_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4072__A0 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5945_ _5961_/B _5945_/B vssd1 vssd1 vccd1 vccd1 _5947_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5876_ _5876_/A _5876_/B vssd1 vssd1 vccd1 vccd1 _5877_/C sky130_fd_sc_hd__xnor2_1
X_4827_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _7194_/C sky130_fd_sc_hd__and2_2
X_7615_ _7623_/CLK _7615_/D vssd1 vssd1 vccd1 vccd1 _7615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4375__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ hold308/X _4443_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7270_/D sky130_fd_sc_hd__mux2_1
X_7546_ _7547_/CLK _7546_/D vssd1 vssd1 vccd1 vccd1 _7546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7477_ _7477_/CLK _7477_/D vssd1 vssd1 vccd1 vccd1 _7477_/Q sky130_fd_sc_hd__dfxtp_1
X_4689_ _4689_/A _4689_/B vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__and2_1
XANTENNA__4470__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5492__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6588__A _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3709_ _6328_/A _5985_/B vssd1 vssd1 vccd1 vccd1 _3724_/A sky130_fd_sc_hd__or2_1
XANTENNA__5324__A0 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6428_ hold95/X _6427_/X _6204_/A vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__a21oi_1
XANTENNA__4222__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _6373_/A _6359_/B vssd1 vssd1 vccd1 vccd1 _7560_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_52_wb_clk_i _7544_/CLK vssd1 vssd1 vccd1 vccd1 _7547_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3740__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3886__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4063__B1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4571__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5817__D _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3915__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4213__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5341__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6291__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _7552_/Q _5808_/A vssd1 vssd1 vccd1 vccd1 _4280_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5730_ _6244_/A _6807_/A _5727_/A _5749_/A vssd1 vssd1 vccd1 vccd1 _5731_/B sky130_fd_sc_hd__a211oi_1
XFILLER_0_57_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7400_ _7400_/CLK _7400_/D vssd1 vssd1 vccd1 vccd1 _7400_/Q sky130_fd_sc_hd__dfxtp_1
X_5661_ _6235_/A _5660_/B _5660_/C vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__a21oi_1
X_4612_ input5/X _4612_/B vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__or2_1
X_5592_ _6840_/A _5561_/X _6875_/A vssd1 vssd1 vccd1 vccd1 _5594_/C sky130_fd_sc_hd__a21o_1
X_4543_ _7480_/Q _7468_/Q _7460_/Q _7254_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4543_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7331_ _7427_/CLK _7331_/D vssd1 vssd1 vccd1 vccd1 _7331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7262_ _7592_/CLK _7262_/D vssd1 vssd1 vccd1 vccd1 _7262_/Q sky130_fd_sc_hd__dfxtp_1
Xhold436 _5405_/X vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold414 _7288_/Q vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _7284_/Q vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 _7622_/Q vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4109__A1 _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold458 _7592_/Q vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 _7253_/Q vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4204__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold469 _7271_/Q vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _4474_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__or2_1
X_6213_ _6345_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _7540_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7193_ _7211_/B _7211_/C _7193_/C vssd1 vssd1 vccd1 vccd1 _7210_/S sky130_fd_sc_hd__and3_4
XANTENNA__7059__B1 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6144_ _6153_/A _6144_/B vssd1 vssd1 vccd1 vccd1 _6144_/Y sky130_fd_sc_hd__nor2_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6075_/Y sky130_fd_sc_hd__nor2_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A _5026_/B vssd1 vssd1 vccd1 vccd1 _5027_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4094__C _4846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6871__A _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6977_ _6978_/B _6977_/B vssd1 vssd1 vccd1 vccd1 _6977_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4391__A _6874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5918__C _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _5947_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5930_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4691__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3719__B _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5859_ _5859_/A vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__inv_2
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4348__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7529_ _7569_/CLK _7529_/D vssd1 vssd1 vccd1 vccd1 _7529_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6111__A _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3735__A _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5848__A1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5161__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6025__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4587__A1 _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4339__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6733__C1 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5336__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5860__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4190_ _7438_/Q _7430_/Q _7414_/Q _7406_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4190_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5071__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6900_ _6900_/A _6989_/A vssd1 vssd1 vccd1 vccd1 _7095_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6831_ _6831_/A _6831_/B _6831_/C vssd1 vssd1 vccd1 vccd1 _6831_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3940__A_N _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6762_ split18/X _6648_/X _6658_/A _6658_/B vssd1 vssd1 vccd1 vccd1 _6763_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_18_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3974_ _6220_/C _4140_/B vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__nor2_2
X_6693_ _6723_/B _6724_/A _6680_/Y vssd1 vssd1 vccd1 vccd1 _6719_/A sky130_fd_sc_hd__a21o_1
X_5713_ _5714_/A _5714_/B _5714_/C vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5644_ _5644_/A _5675_/A _5640_/Y vssd1 vssd1 vccd1 vccd1 _5681_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5246__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold211 _7296_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
X_7314_ _7450_/CLK _7314_/D vssd1 vssd1 vccd1 vccd1 _7314_/Q sky130_fd_sc_hd__dfxtp_1
Xhold200 _7609_/Q vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4150__S _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5575_ _6568_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _5575_/X sky130_fd_sc_hd__or2_1
Xhold233 _5317_/X vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 _7375_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
X_4526_ _4526_/A _4526_/B vssd1 vssd1 vccd1 vccd1 _4526_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold244 _6197_/X vssd1 vssd1 vccd1 vccd1 _6198_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _7353_/Q vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _7623_/Q vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4698_/A _4508_/A _4456_/Y vssd1 vssd1 vccd1 vccd1 _4457_/X sky130_fd_sc_hd__o21a_1
Xhold255 _7241_/X vssd1 vssd1 vccd1 vccd1 _7530_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7245_ input34/X _6225_/B _5139_/Y _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7551_/D sky130_fd_sc_hd__o211a_1
Xhold288 _7419_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _7323_/Q vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_7176_ _7212_/B _7176_/B _7212_/C vssd1 vssd1 vccd1 vccd1 _7191_/S sky130_fd_sc_hd__and3_4
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5770__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6127_ _7603_/Q _6153_/A _6126_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6127_/X sky130_fd_sc_hd__a211o_1
X_4388_ _6111_/A _4389_/B vssd1 vssd1 vccd1 vccd1 _4438_/B sky130_fd_sc_hd__or2_1
XANTENNA__6077__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6922_/A _6056_/X _6057_/Y _4209_/B _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6058_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4361__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5009_ input27/X _4850_/A _4700_/B _4963_/S vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4325__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4018__B1 _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4664__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4416__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5156__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4741__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4235__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6954__C1 _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3690_ _5988_/A _3990_/B vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__nor2_4
XANTENNA__5066__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4732__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5360_ _4111_/X hold546/X _5374_/S vssd1 vssd1 vccd1 vccd1 _7464_/D sky130_fd_sc_hd__mux2_1
X_5291_ hold268/X _4912_/Y _5301_/S vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__mux2_1
X_4311_ _4311_/A _4311_/B vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4242_ _7403_/Q _7395_/Q _7371_/Q _7387_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4242_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5590__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7030_ _7030_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7030_/Y sky130_fd_sc_hd__xnor2_1
X_4173_ _4692_/S _4173_/B vssd1 vssd1 vccd1 vccd1 _4173_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4799__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4653__B _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4145__S _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6814_ _6813_/A _6813_/B _6813_/C _6794_/X vssd1 vssd1 vccd1 vccd1 _6817_/C sky130_fd_sc_hd__o31a_1
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout152_A _7574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4646__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3957_ _7553_/Q _7552_/Q _4128_/A vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__and3_1
X_6745_ _6721_/Y _6782_/A _6766_/A vssd1 vssd1 vccd1 vccd1 _6745_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3888_ _3827_/S _3886_/X _3887_/Y _3882_/Y vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_73_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6676_ _6685_/A _6676_/B vssd1 vssd1 vccd1 vccd1 _6676_/Y sky130_fd_sc_hd__xnor2_1
X_5627_ _5571_/X _6430_/A _5626_/X vssd1 vssd1 vccd1 vccd1 _6463_/S sky130_fd_sc_hd__o21ai_4
XFILLER_0_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5558_ _6532_/A _5566_/B _5556_/B _5556_/A vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4509_ _4876_/B _4601_/A _4509_/C vssd1 vssd1 vccd1 vccd1 _4509_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7228_ _7227_/X _4685_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7623_/D sky130_fd_sc_hd__mux2_1
X_5489_ _5489_/A _5489_/B vssd1 vssd1 vccd1 vccd1 _5489_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3732__B _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7159_ hold231/X _4492_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7594_/D sky130_fd_sc_hd__mux2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6400__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5394__B _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3923__A _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7454_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6219__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output46_A _7559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4860_ input1/X _5031_/S _4162_/B _4859_/X vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__o211a_1
X_3811_ _3915_/A _3807_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _3811_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4791_ hold425/X _4385_/X _4805_/S vssd1 vssd1 vccd1 vccd1 _4791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6530_ _6557_/A _6504_/Y _6557_/C _6529_/X _6505_/C vssd1 vssd1 vccd1 vccd1 _6531_/B
+ sky130_fd_sc_hd__a311oi_2
XFILLER_0_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _6374_/A _7539_/Q _3742_/C vssd1 vssd1 vccd1 vccd1 _6015_/B sky130_fd_sc_hd__or3_2
XFILLER_0_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ _6702_/A vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__inv_6
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6461_ _6461_/A _6461_/B _6522_/B vssd1 vssd1 vccd1 vccd1 _6507_/B sky130_fd_sc_hd__or3_4
XFILLER_0_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5412_ _5854_/C _6702_/A split8/A vssd1 vssd1 vccd1 vccd1 _5438_/A sky130_fd_sc_hd__or3_4
XFILLER_0_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6392_ _6935_/A _6383_/Y _6391_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6392_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5343_ hold463/X _4434_/Y _5355_/S vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5274_ _5273_/X _4897_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _7422_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4225_ _4223_/X _4224_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5130__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7013_ _6962_/A _6864_/A _4037_/X _7001_/X _7012_/X vssd1 vssd1 vccd1 vccd1 _7013_/X
+ sky130_fd_sc_hd__o32a_1
X_4156_ _4162_/B _4154_/X _4155_/X vssd1 vssd1 vccd1 vccd1 _4751_/A sky130_fd_sc_hd__a21o_2
XANTENNA__4316__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3692__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4087_ _6096_/A input11/X _5022_/A vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__mux2_2
XANTENNA__7040__A _7040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5197__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4989_ _4989_/A _4997_/B _4989_/C vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6728_ _6688_/X _6728_/B vssd1 vssd1 vccd1 vccd1 _6729_/B sky130_fd_sc_hd__nand2b_1
X_6659_ split18/X _6648_/X _6658_/X vssd1 vssd1 vccd1 vccd1 _6659_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__3727__B _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3743__A _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4217__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4558__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5121__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5672__A2 _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6385__A0 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4935__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4513__S _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 custom_settings[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput37 io_in[17] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
Xinput26 custom_settings[5] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XFILLER_0_107_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5344__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4468__B _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4546__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__A2 _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ _4033_/B _6331_/B vssd1 vssd1 vccd1 vccd1 _4010_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6683__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _5961_/A _5961_/B _5961_/C vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__and3_1
X_4912_ _4989_/A _4911_/X _4899_/X vssd1 vssd1 vccd1 vccd1 _4912_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__5179__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7631_ _7631_/A vssd1 vssd1 vccd1 vccd1 _7631_/X sky130_fd_sc_hd__buf_1
X_5892_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4843_ hold570/X _4719_/Y _4843_/S vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4931__B _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4774_ _4773_/X _4394_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7277_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6204__A _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7562_ _7587_/CLK _7562_/D vssd1 vssd1 vccd1 vccd1 _7562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3725_ _5977_/B _3733_/B vssd1 vssd1 vccd1 vccd1 _3960_/C sky130_fd_sc_hd__nand2_1
X_7493_ _7498_/CLK hold83/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfxtp_1
X_6513_ _6637_/A _6513_/B _6513_/C vssd1 vssd1 vccd1 vccd1 _6514_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6444_ _6611_/A _6487_/B vssd1 vssd1 vccd1 vccd1 _6474_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3656_ _3656_/A vssd1 vssd1 vccd1 vccd1 _3656_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5351__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ _6375_/A _7230_/D _6375_/C _4015_/B vssd1 vssd1 vccd1 vccd1 _6375_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_101_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_6__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5326_ _4871_/Y hold595/X _5338_/S vssd1 vssd1 vccd1 vccd1 _7445_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5257_ hold522/X _4937_/Y _5265_/S vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5103__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6874__A _6874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__inv_2
X_5188_ _4947_/X hold444/X _5194_/S vssd1 vssd1 vccd1 vccd1 _7384_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4394__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4139_ _6922_/D _4139_/B vssd1 vssd1 vccd1 vccd1 _4139_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__3968__A2 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4090__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6906__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5164__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6784__A _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 _3930_/S0 vssd1 vssd1 vccd1 vccd1 _3913_/S0 sky130_fd_sc_hd__buf_8
Xfanout181 _4244_/S0 vssd1 vssd1 vccd1 vccd1 _4255_/S0 sky130_fd_sc_hd__buf_8
Xfanout170 hold109/X vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__buf_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4751__B _4827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6358__A0 hold66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4384__A2 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold618 _7345_/Q vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4490_ _3935_/A _4487_/A _4106_/X vssd1 vssd1 vccd1 vccd1 _4490_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 _7171_/X vssd1 vssd1 vccd1 vccd1 _7174_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5333__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5074__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold629 _7349_/Q vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _4694_/A _6162_/B _6160_/S vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5884__A2 _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4519__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5111_ _5037_/A _5038_/X _5111_/S vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__mux2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6025_/Y _6088_/Y _6090_/X vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__o21a_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5042_ _5376_/C _5322_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5057_/S sky130_fd_sc_hd__and3_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4418__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6993_ _7009_/B _6993_/B vssd1 vssd1 vccd1 vccd1 _6993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4072__A1 hold610/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5944_ _5956_/A _5961_/A vssd1 vssd1 vccd1 vccd1 _5945_/B sky130_fd_sc_hd__or2_1
XFILLER_0_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5875_ _5876_/A _5876_/B vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__and2_1
X_4826_ _7211_/B _5159_/C _7193_/C vssd1 vssd1 vccd1 vccd1 _4844_/S sky130_fd_sc_hd__and3_4
X_7614_ _7623_/CLK _7614_/D vssd1 vssd1 vccd1 vccd1 _7614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7010__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7010__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7545_ _7547_/CLK _7545_/D vssd1 vssd1 vccd1 vccd1 _7545_/Q sky130_fd_sc_hd__dfxtp_1
X_4757_ hold307/X _4483_/X _4767_/S vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6869__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ _4686_/X _4687_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4689_/B sky130_fd_sc_hd__mux2_1
X_7476_ _7476_/CLK _7476_/D vssd1 vssd1 vccd1 vccd1 _7476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6588__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3708_ _7230_/A _7101_/A vssd1 vssd1 vccd1 vccd1 _5985_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4389__A _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6427_ _6427_/A _6427_/B _4037_/A vssd1 vssd1 vccd1 vccd1 _6427_/X sky130_fd_sc_hd__or3b_1
X_3639_ _3983_/A vssd1 vssd1 vccd1 vccd1 _6225_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6358_ hold66/X hold136/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6358_/X sky130_fd_sc_hd__mux2_1
X_5309_ hold238/X _4912_/Y _5319_/S vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7077__A1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6289_ _6807_/A _6949_/B _6316_/B vssd1 vssd1 vccd1 vccd1 _6290_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7212__B _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7403_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4852__A _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4063__B2 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7001__A1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4290__C _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5315__A1 _4990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6512__B1 _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7068__A1 _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6028__C1 _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7240__A1 hold601/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4054__A1 hold60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ _6223_/A _3990_/B vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5069__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5660_ _6235_/A _5660_/B _5660_/C vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__and3_1
XFILLER_0_84_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4611_ _4113_/Y _4603_/Y _4608_/X _4610_/X vssd1 vssd1 vccd1 vccd1 _4611_/X sky130_fd_sc_hd__o22a_1
X_5591_ _6710_/A _5591_/B _5542_/Y vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4542_ _7280_/Q _7595_/Q _7264_/Q _7488_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4542_/X sky130_fd_sc_hd__mux4_1
X_7330_ _7427_/CLK _7330_/D vssd1 vssd1 vccd1 vccd1 _7330_/Q sky130_fd_sc_hd__dfxtp_1
X_7261_ _7485_/CLK _7261_/D vssd1 vssd1 vccd1 vccd1 _7261_/Q sky130_fd_sc_hd__dfxtp_1
Xhold415 _7393_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5306__A1 _4849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 _4791_/X vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 _7425_/Q vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4474_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__nand2_1
Xhold437 _7466_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold459 _7481_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _4530_/X vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6216_/A _7599_/Q _3685_/B _6211_/Y vssd1 vssd1 vccd1 vccd1 _6212_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_96_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7192_ _7191_/X _4685_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7192_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6143_ _6143_/A vssd1 vssd1 vccd1 vccd1 _6143_/Y sky130_fd_sc_hd__inv_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6328_/A _4228_/Y _6073_/X _6375_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6074_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _6840_/A _4123_/B _5026_/B _4953_/Y _4123_/A vssd1 vssd1 vccd1 vccd1 _5025_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4148__S _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout182_A _7452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5242__A0 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6976_ _6974_/B _6949_/B _6258_/A vssd1 vssd1 vccd1 vccd1 _6977_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4045__A1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4391__B _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5927_ _5927_/A _5927_/B _5927_/C vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__or3_1
XFILLER_0_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5918__D _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5858_ _6244_/A _6771_/A _6773_/A _6690_/A vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3719__C _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4809_ hold216/X _4385_/X _4823_/S vssd1 vssd1 vccd1 vccd1 _4809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5789_ _6972_/A vssd1 vssd1 vccd1 vccd1 _5789_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6599__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7528_ _7570_/CLK _7528_/D vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ _7481_/CLK _7459_/D vssd1 vssd1 vccd1 vccd1 _7459_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5008__A _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6111__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3859__A1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout95_A _3702_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3897__S _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7222__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6025__A2 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit20 split20/A vssd1 vssd1 vccd1 vccd1 _6882_/A sky130_fd_sc_hd__buf_4
XANTENNA__5784__A1 _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3795__B1 _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4521__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5352__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__B _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output76_A _7525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4275__A1 _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6691__B _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7213__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4492__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6830_ _6831_/A _6831_/C _6831_/B vssd1 vssd1 vccd1 vccd1 _6832_/B sky130_fd_sc_hd__a21o_1
X_6761_ _6756_/B _6758_/X _6709_/X vssd1 vssd1 vccd1 vccd1 _6764_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5712_ _5834_/B _5712_/B vssd1 vssd1 vccd1 vccd1 _5714_/C sky130_fd_sc_hd__nand2_1
X_3973_ _7230_/C _3973_/B vssd1 vssd1 vccd1 vccd1 _6328_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3881__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6692_ _6728_/B _6729_/A _6688_/X vssd1 vssd1 vccd1 vccd1 _6724_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5643_ _6808_/A _6311_/A _6611_/A _6771_/A vssd1 vssd1 vccd1 vccd1 _5675_/A sky130_fd_sc_hd__and4_1
XFILLER_0_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5574_ _5546_/B _5573_/Y _5579_/S vssd1 vssd1 vccd1 vccd1 _5576_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 _7598_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
X_7313_ _7450_/CLK _7313_/D vssd1 vssd1 vccd1 vccd1 _7313_/Q sky130_fd_sc_hd__dfxtp_1
X_4525_ _4525_/A _4525_/B vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold234 _7412_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _7306_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _5167_/X vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold245 _7595_/Q vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _7491_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _7319_/Q vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _5117_/X vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4698_/A _4454_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4456_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7244_ _7244_/A _7244_/B vssd1 vssd1 vccd1 vccd1 _7550_/D sky130_fd_sc_hd__or2_1
Xhold289 _5265_/X vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_4387_ _4111_/X hold422/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7250_/D sky130_fd_sc_hd__mux2_1
X_7175_ _7211_/B _7175_/B _7211_/C vssd1 vssd1 vccd1 vccd1 _7192_/S sky130_fd_sc_hd__and3_4
XFILLER_0_0_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5770__B _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6126_ _6153_/A _6126_/B vssd1 vssd1 vccd1 vccd1 _6126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6057_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6882__A _6882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4361__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5008_ _5008_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _5008_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7204__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4018__A1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6959_ _6974_/A _6959_/B vssd1 vssd1 vccd1 vccd1 _6959_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__6963__B1 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3872__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7140__B1 _7558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5172__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4257__A1 _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6792__A _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5206__A0 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6954__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3863__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5347__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5290_ hold295/X _4871_/Y _5302_/S vssd1 vssd1 vccd1 vccd1 _7429_/D sky130_fd_sc_hd__mux2_1
X_4310_ _4474_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _4311_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7131__B1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4241_ _4401_/S _4241_/B vssd1 vssd1 vccd1 vccd1 _4241_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5082__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4172_ _7276_/Q _7591_/Q _7260_/Q _7484_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4173_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6813_ _6813_/A _6813_/B _6813_/C vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_92_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _4846_/A _5990_/A vssd1 vssd1 vccd1 vccd1 _4122_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6744_ _6781_/B _6781_/C _6781_/A vssd1 vssd1 vccd1 vccd1 _6782_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6675_ _6747_/A _6751_/A vssd1 vssd1 vccd1 vccd1 _6675_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3887_ _3886_/S _3883_/X _7363_/Q vssd1 vssd1 vccd1 vccd1 _3887_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5626_ _5571_/A _5571_/B _6430_/B _5625_/X vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__o31a_2
XFILLER_0_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5557_ _5557_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5557_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__5781__A _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4508_ _4508_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _4509_/C sky130_fd_sc_hd__nand2_1
X_5488_ _5556_/A _5488_/B vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__or2_2
XFILLER_0_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7227_ hold266/X _4719_/Y _7227_/S vssd1 vssd1 vccd1 vccd1 _7227_/X sky130_fd_sc_hd__mux2_1
X_4439_ _4487_/B _4439_/B vssd1 vssd1 vccd1 vccd1 _4439_/Y sky130_fd_sc_hd__nor2_1
X_7158_ hold230/X _4529_/X _7166_/S vssd1 vssd1 vccd1 vccd1 _7158_/X sky130_fd_sc_hd__mux2_1
X_6109_ _6025_/Y _6106_/Y _6108_/X vssd1 vssd1 vccd1 vccd1 _6109_/X sky130_fd_sc_hd__o21a_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _6900_/A _7110_/A _7088_/Y _3949_/Y vssd1 vssd1 vccd1 vccd1 _7089_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5987__A1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold524_A _7569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6936__B1 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4947__C1 _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A1 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5167__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5394__C _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6164__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5911__B2 _5811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5911__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7113__B1 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3923__B _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4100__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6219__A2 hold97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7015__B1_N _7014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6027__A _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4770__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3810_ _3808_/X _3809_/X _3931_/S vssd1 vssd1 vccd1 vccd1 _3810_/X sky130_fd_sc_hd__mux2_1
X_4790_ _7212_/A _7212_/B _5322_/B vssd1 vssd1 vccd1 vccd1 _4805_/S sky130_fd_sc_hd__and3_4
XANTENNA__3836__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4402__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3741_ _3742_/C _3741_/B vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__and2b_1
XANTENNA__5667__A2_N _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6155__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3672_ _6864_/A vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__inv_2
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6460_ _6516_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _6522_/B sky130_fd_sc_hd__nor2_1
X_5411_ _5556_/A _6532_/A _6710_/A vssd1 vssd1 vccd1 vccd1 split8/A sky130_fd_sc_hd__or3_4
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6391_ hold132/X _6415_/A _6356_/B hold558/X vssd1 vssd1 vccd1 vccd1 _6391_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6697__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5342_ _4111_/X hold339/X _5356_/S vssd1 vssd1 vccd1 vccd1 _7456_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5273_ hold577/X _4912_/Y _5283_/S vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__mux2_1
X_7012_ _7078_/A _7012_/B _7012_/C _7012_/D vssd1 vssd1 vccd1 vccd1 _7012_/X sky130_fd_sc_hd__or4_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4224_ _7425_/Q _7357_/Q _7349_/Q _7329_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4224_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4945__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4155_ hold60/A _4963_/S _4989_/A vssd1 vssd1 vccd1 vccd1 _4155_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3692__A2 _5952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4316__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4086_ _4945_/B _4440_/A _4846_/C vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__and3_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4988_ _7348_/Q _4948_/B _7349_/Q vssd1 vssd1 vccd1 vccd1 _4989_/C sky130_fd_sc_hd__o21ai_1
X_3939_ _3939_/A _3939_/B vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__or2_1
X_6727_ _6869_/A _6735_/B vssd1 vssd1 vccd1 vccd1 _6734_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6146__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6658_ _6658_/A _6658_/B _6658_/C vssd1 vssd1 vccd1 vccd1 _6658_/X sky130_fd_sc_hd__or3_4
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7623_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5609_ _5609_/A _5609_/B vssd1 vssd1 vccd1 vccd1 _6462_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4252__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6589_ _6621_/B _6622_/A _6621_/A vssd1 vssd1 vccd1 vccd1 _6619_/A sky130_fd_sc_hd__o21bai_4
XANTENNA_hold641_A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 custom_settings[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6137__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput27 custom_settings[6] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_109_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 io_in[18] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4243__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4546__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__A1 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5960_ _5960_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5961_/C sky130_fd_sc_hd__xnor2_1
X_4911_ _4162_/B _4907_/X _4908_/Y _4910_/X vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__a31o_1
X_5891_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__and2_1
X_7630_ _7630_/A vssd1 vssd1 vccd1 vccd1 _7630_/X sky130_fd_sc_hd__buf_1
XFILLER_0_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4387__A0 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4842_ _4841_/X _4637_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7306_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3809__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6376__A1 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4773_ hold385/X _4434_/Y _4785_/S vssd1 vssd1 vccd1 vccd1 _4773_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7561_ _7577_/CLK _7561_/D vssd1 vssd1 vccd1 vccd1 _7561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6128__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7492_ _7498_/CLK hold77/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
X_6512_ _6513_/B _6513_/C _6637_/A vssd1 vssd1 vccd1 vccd1 _6512_/Y sky130_fd_sc_hd__a21oi_1
X_3724_ _3724_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _5977_/D sky130_fd_sc_hd__or2_1
X_6443_ _5576_/B _6442_/Y _6463_/S vssd1 vssd1 vccd1 vccd1 _6487_/B sky130_fd_sc_hd__mux2_1
X_3655_ _3683_/A vssd1 vssd1 vccd1 vccd1 _6216_/B sky130_fd_sc_hd__inv_2
XANTENNA__4234__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6374_ _6374_/A _6374_/B vssd1 vssd1 vccd1 vccd1 _7230_/D sky130_fd_sc_hd__nand2_1
X_5325_ hold594/X _4887_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__mux2_1
X_5256_ hold335/X _4897_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _5256_/X sky130_fd_sc_hd__mux2_1
X_4207_ _4689_/A _4205_/X _4206_/Y _4201_/Y vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__a2bb2o_2
X_5187_ hold443/X _4964_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5270__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4138_ _5811_/B _6415_/B vssd1 vssd1 vccd1 vccd1 _4139_/B sky130_fd_sc_hd__nand2_1
X_4069_ hold97/X _6872_/B _6329_/A vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7197__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3738__B _7559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6119__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6119__B2 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6130__A _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold591_A _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5180__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 _7452_/Q vssd1 vssd1 vccd1 vccd1 _4244_/S0 sky130_fd_sc_hd__buf_8
Xfanout160 _7572_/Q vssd1 vssd1 vccd1 vccd1 _6872_/B sky130_fd_sc_hd__buf_6
Xfanout171 _4001_/D vssd1 vssd1 vccd1 vccd1 _6920_/A sky130_fd_sc_hd__buf_4
Xfanout193 _7360_/Q vssd1 vssd1 vccd1 vccd1 _3930_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4605__A1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5030__A1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3664__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5355__S _5355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 _7174_/X vssd1 vssd1 vccd1 vccd1 _7599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold619 _5099_/X vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4541__B1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5110_ _5109_/X _4996_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _7350_/D sky130_fd_sc_hd__mux2_1
X_6090_ _7351_/Q _6153_/A _6089_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__a211o_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5041_ _5375_/C _5159_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5058_/S sky130_fd_sc_hd__and3_4
XANTENNA__4519__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5097__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5090__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4844__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_6992_ _6235_/A _6922_/B _6991_/X _7098_/A vssd1 vssd1 vccd1 vccd1 _6992_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5943_ _5943_/A _5958_/B vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__and2_1
XFILLER_0_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5874_ _5905_/A _5874_/B vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7613_ _7621_/CLK _7613_/D vssd1 vssd1 vccd1 vccd1 _7613_/Q sky130_fd_sc_hd__dfxtp_1
X_4825_ _4748_/A _4825_/B vssd1 vssd1 vccd1 vccd1 _7193_/C sky130_fd_sc_hd__and2b_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5021__B2 _4083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7544_ _7544_/CLK _7544_/D vssd1 vssd1 vccd1 vccd1 _7544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4756_ _4755_/X _4394_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7269_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4687_ _7483_/Q _7471_/Q _7463_/Q _7257_/Q _7452_/Q _7453_/Q vssd1 vssd1 vccd1 vccd1
+ _4687_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7475_ _7475_/CLK hold57/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3707_ _7043_/S _6989_/A vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3638_ _3733_/A vssd1 vssd1 vccd1 vccd1 _5977_/B sky130_fd_sc_hd__inv_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6426_ hold94/X _6427_/A vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__nand2_1
X_6357_ _6357_/A _7231_/B _6357_/C _6351_/A vssd1 vssd1 vccd1 vccd1 _6372_/S sky130_fd_sc_hd__or4b_4
XFILLER_0_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5308_ hold341/X _4871_/Y _5320_/S vssd1 vssd1 vccd1 vccd1 _7437_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5088__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6288_ _6949_/B _6316_/B _6807_/A vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__a21o_1
X_5239_ hold584/X _4937_/Y _5247_/S vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4835__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5260__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4852__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7577_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4446__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5175__S _5175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6795__A _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5079__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6028__B1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6035__A _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4610_ _5008_/A _4609_/X _4118_/B vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__a21o_1
X_5590_ _6875_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5085__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4541_ _4539_/Y _4638_/C _4529_/S vssd1 vssd1 vccd1 vccd1 _4541_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold427 _7480_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _5208_/X vssd1 vssd1 vccd1 vccd1 _7393_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7260_ _7592_/CLK _7260_/D vssd1 vssd1 vccd1 vccd1 _7260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4472_ _4667_/B _4471_/X _4468_/Y vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__o21ai_2
Xhold405 _5280_/X vssd1 vssd1 vccd1 vccd1 _7425_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold438 _5363_/X vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _7478_/Q vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_7191_ hold645/X _4719_/Y _7191_/S vssd1 vssd1 vccd1 vccd1 _7191_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6211_ _7540_/Q _6211_/B vssd1 vssd1 vccd1 vccd1 _6211_/Y sky130_fd_sc_hd__nor2_1
X_6142_ _4601_/C _6144_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__mux2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6073_ _6025_/Y _6070_/Y _6072_/X vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__o21a_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5026_/B _5023_/X _5024_/S vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout175_A _7455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4953__A _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4672__B _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4045__A2 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6975_ _3716_/Y _6264_/B _6974_/X _7070_/A _7009_/A vssd1 vssd1 vccd1 vccd1 _6975_/X
+ sky130_fd_sc_hd__o32a_1
X_5926_ _5927_/A _5927_/B _5927_/C vssd1 vssd1 vccd1 vccd1 _5947_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _6273_/A _6851_/A vssd1 vssd1 vccd1 vccd1 _7109_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4808_ _7212_/B _7176_/B _5322_/B vssd1 vssd1 vccd1 vccd1 _4823_/S sky130_fd_sc_hd__and3_4
X_5788_ _6808_/A _5788_/B _6802_/B _5788_/D vssd1 vssd1 vccd1 vccd1 _6972_/A sky130_fd_sc_hd__and4_1
X_4739_ hold218/X _4580_/X _4745_/S vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__mux2_1
X_7527_ _7570_/CLK _7527_/D vssd1 vssd1 vccd1 vccd1 _7527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7458_ _7592_/CLK _7458_/D vssd1 vssd1 vccd1 vccd1 _7458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6409_ input37/X _6408_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6409_/X sky130_fd_sc_hd__mux2_1
X_7389_ _4004_/A _7389_/D vssd1 vssd1 vccd1 vccd1 _7389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout88_A _6022_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4108__A1_N _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5233__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3795__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5784__A2 _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit32 _5556_/A vssd1 vssd1 vccd1 vccd1 _6445_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4419__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5694__A _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4802__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6733__A1 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4103__A _4103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5224__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ _6710_/B split7/X _6758_/X _6759_/Y vssd1 vssd1 vccd1 vccd1 _6760_/X sky130_fd_sc_hd__a2bb2o_1
X_5711_ _5711_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5712_/B sky130_fd_sc_hd__or2_1
X_3972_ _7230_/C _3972_/B vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__or2_2
XFILLER_0_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4983__B1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6691_ _6691_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6729_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3881__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5642_ _5642_/A vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__inv_2
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5573_ _5573_/A _5573_/B vssd1 vssd1 vccd1 vccd1 _5573_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold202 _7418_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
X_7312_ _7413_/CLK _7312_/D vssd1 vssd1 vccd1 vccd1 _7312_/Q sky130_fd_sc_hd__dfxtp_1
X_4524_ _4672_/B _6126_/B vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4013__A _5952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 _5251_/X vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _7293_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _7527_/Q vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold268 _7430_/Q vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _7390_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _7297_/Q vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ _4405_/X _4460_/B _4508_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7243_ input32/X _6225_/B _5135_/X _6373_/A vssd1 vssd1 vccd1 vccd1 _7549_/D sky130_fd_sc_hd__o211a_1
X_4386_ hold421/X _4385_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4386_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4667__B _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold279 _7330_/Q vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5770__C _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7174_ _7173_/Y _5132_/B _7174_/S vssd1 vssd1 vccd1 vccd1 _7174_/X sky130_fd_sc_hd__mux2_1
X_6125_ _6125_/A vssd1 vssd1 vccd1 vccd1 _6125_/Y sky130_fd_sc_hd__inv_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6328_/A _4209_/B _6055_/X _6375_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6056_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _4238_/A _5001_/B _5024_/S vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5215__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6963__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6958_ _6872_/A _6926_/Y _6956_/X _6957_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7584_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6889_ _6836_/B _6888_/A _6836_/C vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__a21oi_1
X_5909_ _5875_/X _5879_/B _5907_/Y _5955_/A vssd1 vssd1 vccd1 vccd1 _5909_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3872__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4069__S _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6403__B1 _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6954__B2 _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3863__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5363__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3672__A _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4240_ _7443_/Q _7435_/Q _7419_/Q _7411_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4241_/B sky130_fd_sc_hd__mux4_1
X_4171_ _4529_/S _4171_/B vssd1 vssd1 vccd1 vccd1 _4171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4707__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7198__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6812_ _6806_/X _6809_/A _6859_/B _6811_/A vssd1 vssd1 vccd1 vccd1 _6813_/C sky130_fd_sc_hd__o211a_1
XANTENNA__4008__A _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4956__A0 _4955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6743_ _6786_/A _6789_/A _6789_/B vssd1 vssd1 vccd1 vccd1 _6781_/C sky130_fd_sc_hd__nand3b_1
X_3955_ _6911_/A _3955_/B vssd1 vssd1 vccd1 vccd1 _3965_/D sky130_fd_sc_hd__xnor2_1
X_6674_ _6674_/A _6674_/B vssd1 vssd1 vccd1 vccd1 _6751_/A sky130_fd_sc_hd__nor2_2
XANTENNA__6223__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3886_ _3884_/X _3885_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout138_A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5625_ _6532_/A _5565_/B _5571_/A _5568_/B _6710_/A vssd1 vssd1 vccd1 vccd1 _5625_/X
+ sky130_fd_sc_hd__o32a_1
X_5556_ _5556_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5273__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4507_ _4554_/A _4507_/B vssd1 vssd1 vccd1 vccd1 _4507_/X sky130_fd_sc_hd__or2_1
X_5487_ _5486_/C _5495_/S _6656_/A vssd1 vssd1 vccd1 vccd1 _5488_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5781__B _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7226_ _7225_/X _4637_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7622_/D sky130_fd_sc_hd__mux2_1
X_4438_ _6120_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4439_/B sky130_fd_sc_hd__and2_1
XANTENNA__6330__C1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7157_ hold312/X _4443_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7593_/D sky130_fd_sc_hd__mux2_1
X_4369_ _7403_/Q _7395_/Q _7371_/Q _7387_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4369_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3790__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6108_ _7601_/Q _6162_/A _6107_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6108_/X sky130_fd_sc_hd__a211o_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7086_/Y _7087_/X _6900_/A vssd1 vssd1 vccd1 vccd1 _7088_/Y sky130_fd_sc_hd__o21ai_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _6039_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6039_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7189__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6936__A1 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5372__A0 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5183__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4527__S _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4770__B _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3667__A _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3836__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ _6374_/A _3763_/A vssd1 vssd1 vccd1 vccd1 _3741_/B sky130_fd_sc_hd__nor2_2
X_3671_ _6742_/A vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__inv_2
X_5410_ _4685_/X _5409_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7491_/D sky130_fd_sc_hd__mux2_1
X_6390_ _6389_/X hold610/X _6414_/S vssd1 vssd1 vccd1 vccd1 _7573_/D sky130_fd_sc_hd__mux2_1
X_5341_ hold338/X _4385_/X _5355_/S vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7104__A1 _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5093__S _5093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5272_ hold395/X _4871_/Y _5284_/S vssd1 vssd1 vccd1 vccd1 _7421_/D sky130_fd_sc_hd__mux2_1
X_7011_ _7003_/X _7010_/X _7043_/S vssd1 vssd1 vccd1 vccd1 _7012_/D sky130_fd_sc_hd__mux2_1
X_4223_ _7321_/Q _7337_/Q _7313_/Q _7449_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4223_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4154_ _7569_/Q input14/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4085_ _4015_/B _4290_/D _4946_/A vssd1 vssd1 vccd1 vccd1 _4846_/C sky130_fd_sc_hd__o21a_4
XANTENNA__6218__A _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6091__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6918__A1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4987_ _4982_/X _4983_/X _4986_/X _4162_/B vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__o2bb2a_1
X_6726_ _6735_/B vssd1 vssd1 vccd1 vccd1 _6726_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3938_ _4972_/A _6084_/A vssd1 vssd1 vccd1 vccd1 _3939_/B sky130_fd_sc_hd__nor2_1
X_3869_ _7397_/Q _7389_/Q _7365_/Q _7381_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3869_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6657_ _6764_/B _6764_/A _6653_/Y vssd1 vssd1 vccd1 vccd1 _6658_/C sky130_fd_sc_hd__or3b_4
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5354__A0 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6588_ _6628_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _6622_/A sky130_fd_sc_hd__nor2_1
X_5608_ _5608_/A vssd1 vssd1 vccd1 vccd1 _5621_/C sky130_fd_sc_hd__inv_2
XANTENNA__4252__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5539_ _5488_/X _5493_/A _5554_/A _5517_/X _5537_/Y vssd1 vssd1 vccd1 vccd1 _5539_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4201__A _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5657__A1 _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7209_ hold306/X _4719_/Y _7209_/S vssd1 vssd1 vccd1 vccd1 _7209_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5409__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4347__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6082__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7031__B1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 custom_settings[24] vssd1 vssd1 vccd1 vccd1 _4004_/B sky130_fd_sc_hd__buf_1
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 custom_settings[7] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XANTENNA__4810__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput39 io_in[25] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4243__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3934__B _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4111__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output51_A _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6073__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4608__C1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4910_ _6048_/A _4986_/S _4351_/X _4909_/Y _4963_/S vssd1 vssd1 vccd1 vccd1 _4910_/X
+ sky130_fd_sc_hd__o221a_1
X_5890_ _5913_/B _5890_/B vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4841_ hold212/X _4679_/X _4843_/S vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5088__S _5094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3809__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772_ hold387/X _4111_/X _4786_/S vssd1 vssd1 vccd1 vccd1 _7276_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7560_ _7579_/CLK _7560_/D vssd1 vssd1 vccd1 vccd1 _7560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7491_ _7598_/CLK _7491_/D vssd1 vssd1 vccd1 vccd1 _7491_/Q sky130_fd_sc_hd__dfxtp_1
X_3723_ _3724_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _4267_/C sky130_fd_sc_hd__nor2_4
X_6511_ _6513_/B _6513_/C vssd1 vssd1 vccd1 vccd1 _6511_/X sky130_fd_sc_hd__and2_1
XANTENNA__4720__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5336__A0 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6442_ _6442_/A _6442_/B vssd1 vssd1 vccd1 vccd1 _6442_/Y sky130_fd_sc_hd__xnor2_1
X_3654_ _6216_/A vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__inv_2
XANTENNA__4234__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6373_ _6373_/A _6373_/B vssd1 vssd1 vccd1 vccd1 _7567_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5324_ _4849_/X hold355/X _5338_/S vssd1 vssd1 vccd1 vccd1 _7444_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4021__A _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5255_ hold334/X _4912_/Y _5265_/S vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__mux2_1
X_4206_ _4688_/S _4202_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _4206_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5186_ _4921_/X _5185_/X _5194_/S vssd1 vssd1 vccd1 vccd1 _7383_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6064__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4137_ _6417_/B _7230_/B vssd1 vssd1 vccd1 vccd1 _6415_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _4068_/A _4068_/B vssd1 vssd1 vccd1 vccd1 _7249_/S sky130_fd_sc_hd__or2_4
XANTENNA__5787__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6709_ _6647_/B _6708_/Y _6709_/S vssd1 vssd1 vccd1 vccd1 _6709_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4630__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6130__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 _4686_/S0 vssd1 vssd1 vccd1 vccd1 _4691_/S0 sky130_fd_sc_hd__buf_8
Xfanout150 _6864_/A vssd1 vssd1 vccd1 vccd1 _6637_/A sky130_fd_sc_hd__buf_6
Xfanout161 _6900_/A vssd1 vssd1 vccd1 vccd1 _4084_/A sky130_fd_sc_hd__buf_6
Xfanout172 _6922_/A vssd1 vssd1 vccd1 vccd1 _6417_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout194 _4360_/B vssd1 vssd1 vccd1 vccd1 _4667_/B sky130_fd_sc_hd__buf_6
XANTENNA__6055__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4805__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7004__B1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold609 _7555_/Q vssd1 vssd1 vccd1 vccd1 _3733_/A sky130_fd_sc_hd__buf_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5371__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5040_ hold567/X _5022_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _7315_/D sky130_fd_sc_hd__mux2_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6046__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6991_ _6244_/A _6935_/A _7551_/Q vssd1 vssd1 vccd1 vccd1 _6991_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4715__S _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5942_ _5941_/A _5941_/B _5941_/C vssd1 vssd1 vccd1 vccd1 _5958_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5873_ _5904_/B _5872_/C _5872_/A vssd1 vssd1 vccd1 vccd1 _5874_/B sky130_fd_sc_hd__a21oi_1
X_7612_ _7620_/CLK _7612_/D vssd1 vssd1 vccd1 vccd1 _7612_/Q sky130_fd_sc_hd__dfxtp_1
X_4824_ _4823_/X _4685_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7299_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4755_ hold228/X _4434_/Y _4767_/S vssd1 vssd1 vccd1 vccd1 _4755_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7543_ _7590_/CLK _7543_/D vssd1 vssd1 vccd1 vccd1 _7543_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4780__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3706_ _4036_/A _3780_/A vssd1 vssd1 vccd1 vccd1 _6910_/A sky130_fd_sc_hd__nand2_2
X_4686_ _7283_/Q _7598_/Q _7267_/Q _7491_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4686_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7474_ _7541_/CLK _7474_/D vssd1 vssd1 vccd1 vccd1 _7474_/Q sky130_fd_sc_hd__dfxtp_1
X_3637_ _7558_/Q vssd1 vssd1 vccd1 vccd1 _7090_/A sky130_fd_sc_hd__inv_2
X_6425_ hold107/X _6424_/X _6204_/A vssd1 vssd1 vccd1 vccd1 _6425_/Y sky130_fd_sc_hd__a21oi_1
X_6356_ _6417_/B _6356_/B vssd1 vssd1 vccd1 vccd1 _6357_/C sky130_fd_sc_hd__nor2_1
X_5307_ hold340/X _4887_/X _5319_/S vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5281__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _7557_/Q _6287_/B vssd1 vssd1 vccd1 vccd1 _6316_/B sky130_fd_sc_hd__nand2_1
X_5238_ _4897_/X hold275/X _5248_/S vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__mux2_1
X_5169_ hold325/X _4580_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6037__A1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4048__A0 hold97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4599__A1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4446__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3765__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4771__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7477_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4523__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5980__A _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5191__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6028__A1 _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5366__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3675__A _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4762__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4540_ _7604_/Q _4540_/B vssd1 vssd1 vccd1 vccd1 _4638_/C sky130_fd_sc_hd__or2_2
Xhold417 _7449_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ _4470_/X _4469_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4471_/X sky130_fd_sc_hd__mux2_1
Xhold406 _7290_/Q vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold439 _7486_/Q vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold428 _7424_/Q vssd1 vssd1 vccd1 vccd1 hold428/X sky130_fd_sc_hd__dlygate4sd3_1
X_7190_ _7189_/X _4637_/X _7192_/S vssd1 vssd1 vccd1 vccd1 _7190_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4514__A1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6210_ _4723_/Y _6210_/B _6345_/A vssd1 vssd1 vccd1 vccd1 _6210_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6141_ _6140_/X hold80/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6197__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6072_ _7349_/Q _6162_/A _6071_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4278__B1 _4143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5026_/B _4999_/X _4261_/Y vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6974_ _6974_/A _6974_/B _6974_/C vssd1 vssd1 vccd1 vccd1 _6974_/X sky130_fd_sc_hd__and3_1
XFILLER_0_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5925_ _5925_/A _5961_/A vssd1 vssd1 vccd1 vccd1 _5927_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5856_ _5856_/A _5856_/B vssd1 vssd1 vccd1 vccd1 _5864_/A sky130_fd_sc_hd__or2_1
X_4807_ _7211_/B _7175_/B _5159_/C vssd1 vssd1 vccd1 vccd1 _4824_/S sky130_fd_sc_hd__and3_4
XFILLER_0_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5276__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5787_ _6808_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _5787_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4738_ hold345/X _4492_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7263_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4753__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5950__B1 _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7526_ _7538_/CLK _7526_/D vssd1 vssd1 vccd1 vccd1 _7526_/Q sky130_fd_sc_hd__dfxtp_1
X_7457_ _7485_/CLK _7457_/D vssd1 vssd1 vccd1 vccd1 _7457_/Q sky130_fd_sc_hd__dfxtp_1
X_4669_ _7274_/Q _7614_/Q _7606_/Q _7622_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4669_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6408_ _7123_/A _6383_/Y _6407_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6408_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7388_ _7396_/CLK _7388_/D vssd1 vssd1 vccd1 vccd1 _7388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6339_ _6339_/A _7074_/B vssd1 vssd1 vccd1 vccd1 _7100_/C sky130_fd_sc_hd__or2_1
XFILLER_0_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5694__B _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5186__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4744__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4090__S _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3942__B _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3971_ _5132_/A _7098_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _3972_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4983__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5710_ _5711_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5834_/B sky130_fd_sc_hd__nand2_1
X_6690_ _6690_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6690_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5641_ _6808_/A _6611_/A _6532_/A _6311_/A vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4735__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5572_ _5529_/Y _5572_/B vssd1 vssd1 vccd1 vccd1 _5573_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7311_ _4004_/A _7311_/D vssd1 vssd1 vccd1 vccd1 _7311_/Q sky130_fd_sc_hd__dfxtp_1
X_4523_ _4667_/B _4518_/X _4522_/X vssd1 vssd1 vccd1 vccd1 _6126_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 _7278_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _7266_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold214 _4050_/X vssd1 vssd1 vccd1 vccd1 _7340_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6488__A1 _6481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7242_ input31/X _6225_/B _5133_/Y _6373_/A vssd1 vssd1 vccd1 vccd1 _7548_/D sky130_fd_sc_hd__o211a_1
Xhold269 _5291_/X vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _5201_/X vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _4819_/X vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _7611_/Q vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _4454_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4508_/A sky130_fd_sc_hd__or2_1
X_4385_ _4529_/S _4278_/X _4384_/X _4171_/Y vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__a31o_4
XANTENNA__5770__D _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7173_ _3728_/A _7172_/X _6417_/B vssd1 vssd1 vccd1 vccd1 _7173_/Y sky130_fd_sc_hd__a21oi_1
X_6124_ _6123_/B _6126_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__mux2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4346__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6055_ _6025_/Y _6052_/Y _6054_/X vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__o21a_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _6844_/A _4905_/B _5005_/Y _4116_/Y vssd1 vssd1 vccd1 vccd1 _5006_/X sky130_fd_sc_hd__a211o_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ input32/X _4021_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _6957_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6412__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6963__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5908_ _5875_/X _5879_/B _5907_/Y vssd1 vssd1 vccd1 vccd1 _5933_/B sky130_fd_sc_hd__o21a_1
X_6888_ _6888_/A _6891_/B vssd1 vssd1 vccd1 vccd1 _6888_/Y sky130_fd_sc_hd__nand2_1
X_5839_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__or2_1
XFILLER_0_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7509_ _7537_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5151__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4337__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4662__B1 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6403__B2 hold60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6954__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4414__B1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4965__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5390__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4170_ _4170_/A _4170_/B vssd1 vssd1 vccd1 vccd1 _4171_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4328__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5850__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6811_ _6811_/A _6811_/B vssd1 vssd1 vccd1 vccd1 _6860_/A sky130_fd_sc_hd__and2_1
XFILLER_0_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4008__B _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4500__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6742_ _6742_/A _6742_/B vssd1 vssd1 vccd1 vccd1 _6789_/B sky130_fd_sc_hd__xnor2_2
X_3954_ _3954_/A _3954_/B _3954_/C _3953_/X vssd1 vssd1 vccd1 vccd1 _3955_/B sky130_fd_sc_hd__or4b_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3885_ _7426_/Q _7358_/Q _7350_/Q _7330_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3885_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6673_ _6673_/A _6673_/B vssd1 vssd1 vccd1 vccd1 _6674_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5624_ _6718_/A _5580_/B _5623_/X vssd1 vssd1 vccd1 vccd1 _6430_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5381__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _5492_/B _5554_/Y _5555_/S vssd1 vssd1 vccd1 vccd1 _5556_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7107__C1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4506_ _4999_/B _4508_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _4507_/B sky130_fd_sc_hd__o21a_1
X_5486_ _6568_/A split8/X _5486_/C _5477_/X vssd1 vssd1 vccd1 vccd1 _6656_/A sky130_fd_sc_hd__or4b_4
X_7225_ hold403/X _4679_/X _7227_/S vssd1 vssd1 vccd1 vccd1 _7225_/X sky130_fd_sc_hd__mux2_1
X_4437_ _6120_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6424__C_N _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7156_ hold311/X _4483_/X _7166_/S vssd1 vssd1 vccd1 vccd1 _7156_/X sky130_fd_sc_hd__mux2_1
X_4368_ _7443_/Q _7435_/Q _7419_/Q _7411_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4368_/X sky130_fd_sc_hd__mux4_1
X_6107_ _6162_/A _6107_/B vssd1 vssd1 vccd1 vccd1 _6107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3790__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4299_ _4360_/B _4294_/X _4298_/X vssd1 vssd1 vccd1 vccd1 _6071_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__3802__S _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4694__A _4694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7087_ _7129_/A _7085_/A _7085_/B _6893_/Y _6844_/B vssd1 vssd1 vccd1 vccd1 _7087_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7070__A _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6038_ _6328_/A _4902_/A _6037_/X _6375_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6038_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6397__A0 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6936__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4947__A1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3757__B _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3773__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5124__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4883__A0 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4938__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _6518_/A vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5363__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5374__S _5374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5340_ _5376_/A _7212_/B _7176_/B vssd1 vssd1 vccd1 vccd1 _5355_/S sky130_fd_sc_hd__and3_4
XFILLER_0_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7104__A2 _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5115__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5271_ hold394/X _4887_/X _5283_/S vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6312__B1 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4222_ _7401_/Q _7393_/Q _7369_/Q _7385_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4222_/X sky130_fd_sc_hd__mux4_1
X_7010_ _6989_/A _7040_/C _7009_/Y _7008_/X _5879_/A vssd1 vssd1 vccd1 vccd1 _7010_/X
+ sky130_fd_sc_hd__a32o_1
X_4153_ _4789_/B _4750_/B vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__nor2_4
X_4084_ _4084_/A _5985_/A _4121_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4019__A _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ _6075_/A _4985_/Y _4986_/S vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout150_A _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6234__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3937_ _3937_/A _3937_/B vssd1 vssd1 vccd1 vccd1 _3937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6725_ _6679_/Y _6724_/Y split7/A vssd1 vssd1 vccd1 vccd1 _6735_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3868_ _7437_/Q _7429_/Q _7413_/Q _7405_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3868_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6656_ _6656_/A _6656_/B vssd1 vssd1 vccd1 vccd1 _6764_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3799_ _7481_/Q _7469_/Q _7461_/Q _7255_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3799_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4689__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5284__S _5284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6587_ _6586_/B _6586_/C _6629_/A vssd1 vssd1 vccd1 vccd1 _6621_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5607_ _6462_/A _5607_/B vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__nand2_1
X_5538_ _5488_/X _5493_/A _5554_/A _5517_/X _5537_/A vssd1 vssd1 vccd1 vccd1 _5538_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5106__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7208_ _7207_/X _4637_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7614_/D sky130_fd_sc_hd__mux2_1
X_5469_ _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5469_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5657__A2 _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7139_ _7020_/A _6270_/Y _7137_/X _7138_/X vssd1 vssd1 vccd1 vccd1 _7139_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_55_wb_clk_i _7544_/CLK vssd1 vssd1 vccd1 vccd1 _7582_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4363__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6144__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3768__A _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 custom_settings[25] vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__buf_1
XFILLER_0_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5194__S _5194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5345__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput29 custom_settings[8] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4856__B1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5369__S _5373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ hold494/X _4589_/X _4844_/S vssd1 vssd1 vccd1 vccd1 _7305_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ hold386/X _4385_/X _4785_/S vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6989__A _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6510_ _6521_/A _6509_/B _6508_/X vssd1 vssd1 vccd1 vccd1 _6513_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7490_ _7597_/CLK _7490_/D vssd1 vssd1 vccd1 vccd1 _7490_/Q sky130_fd_sc_hd__dfxtp_1
X_3722_ _6333_/A _3721_/Y _4084_/A vssd1 vssd1 vccd1 vccd1 _4124_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3653_ hold72/X vssd1 vssd1 vccd1 vccd1 _3653_/Y sky130_fd_sc_hd__inv_2
X_6441_ _6441_/A vssd1 vssd1 vccd1 vccd1 _6441_/Y sky130_fd_sc_hd__inv_2
X_6372_ _7530_/Q hold130/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6372_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3898__A1 _3665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5323_ hold354/X _4864_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7089__A1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6220__C _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5254_ hold287/X _4871_/Y _5266_/S vssd1 vssd1 vccd1 vccd1 _7413_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5185_ hold409/X _4937_/Y _5193_/S vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__mux2_1
X_4205_ _4203_/X _4204_/X _4401_/S vssd1 vssd1 vccd1 vccd1 _4205_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout198_A _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4136_ _4850_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5133__A _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4067_ _4067_/A _4067_/B _4067_/C _4066_/X vssd1 vssd1 vccd1 vccd1 _4068_/B sky130_fd_sc_hd__or4b_1
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5787__B _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5279__S _5283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5024__A0 _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7013__A1 _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4969_ _6075_/A _4968_/B _4945_/B vssd1 vssd1 vccd1 vccd1 _4969_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6708_ _6708_/A _6708_/B vssd1 vssd1 vccd1 vccd1 _6708_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5327__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6639_ _6857_/A _6639_/B vssd1 vssd1 vccd1 vccd1 _6640_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4212__A _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6139__A _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 _6844_/A vssd1 vssd1 vccd1 vccd1 _6771_/A sky130_fd_sc_hd__buf_4
Xfanout173 _6427_/B vssd1 vssd1 vccd1 vccd1 _6922_/A sky130_fd_sc_hd__buf_4
Xfanout151 _7575_/Q vssd1 vssd1 vccd1 vccd1 _6864_/A sky130_fd_sc_hd__clkbuf_8
Xfanout162 _7558_/Q vssd1 vssd1 vccd1 vccd1 _6900_/A sky130_fd_sc_hd__clkbuf_8
Xfanout184 _7452_/Q vssd1 vssd1 vccd1 vccd1 _4686_/S0 sky130_fd_sc_hd__buf_8
Xfanout195 _7343_/Q vssd1 vssd1 vccd1 vccd1 _4360_/B sky130_fd_sc_hd__buf_8
XANTENNA__5189__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4821__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5318__A1 _4996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6515__B1 _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4122__A _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6818__A1 _6851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6990_ _7009_/A _7009_/B _6960_/B _6989_/Y vssd1 vssd1 vccd1 vccd1 _6990_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7243__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5888__A _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _5941_/A _5941_/B _5941_/C vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__or3_1
XFILLER_0_48_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7557_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5872_ _5872_/A _5904_/B _5872_/C vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__and3_1
X_4823_ hold486/X _4719_/Y _4823_/S vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__mux2_1
X_7611_ _7623_/CLK _7611_/D vssd1 vssd1 vccd1 vccd1 _7611_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4731__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ hold353/X _4111_/X _4768_/S vssd1 vssd1 vccd1 vccd1 _7268_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7542_ _7581_/CLK _7542_/D vssd1 vssd1 vccd1 vccd1 _7542_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5309__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3705_ _4036_/A _3780_/A vssd1 vssd1 vccd1 vccd1 _3705_/X sky130_fd_sc_hd__and2_2
X_7473_ _7475_/CLK _7473_/D vssd1 vssd1 vccd1 vccd1 _7473_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4685_ _4685_/A _4685_/B vssd1 vssd1 vccd1 vccd1 _4685_/X sky130_fd_sc_hd__or2_4
X_3636_ _5788_/B vssd1 vssd1 vccd1 vccd1 _6261_/A sky130_fd_sc_hd__inv_2
X_6424_ _6427_/A _6427_/B _6326_/B vssd1 vssd1 vccd1 vccd1 _6424_/X sky130_fd_sc_hd__or3b_1
XANTENNA__4032__A _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6355_ _5980_/Y _6354_/Y _6015_/C vssd1 vssd1 vccd1 vccd1 _7231_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5306_ hold400/X _4849_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3871__A _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6286_ _6939_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6909_/B sky130_fd_sc_hd__nand2_1
X_5237_ hold274/X _4912_/Y _5247_/S vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__mux2_1
X_5168_ hold223/X _4492_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7375_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3810__S _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5099_ _4872_/B _4887_/X _5111_/S vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__mux2_1
X_4119_ _4119_/A _4290_/D vssd1 vssd1 vccd1 vccd1 _4134_/D sky130_fd_sc_hd__nor2_2
XANTENNA__6393__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3781__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4088__S _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5236__A0 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7225__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4816__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6028__A2 _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6736__A0 _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3956__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold407 _7487_/Q vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _5334_/X vssd1 vssd1 vccd1 vccd1 _7449_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4470_ _7270_/Q _7610_/Q _7602_/Q _7618_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4470_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold429 _5277_/X vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5382__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6140_ _6427_/B _6138_/X _6139_/Y _4553_/B _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6140_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3691__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3722__B1 _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6071_ _6356_/B _6071_/B vssd1 vssd1 vccd1 vccd1 _6071_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4278__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5114__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5022_ _5022_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__or2_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7216__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5411__A _5556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6975__B1 _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6973_ _6989_/A _7002_/A _6972_/X _6832_/A _5879_/A vssd1 vssd1 vccd1 vccd1 _6973_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5924_ _5923_/A _5923_/B _5923_/C vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3884__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5855_ _5855_/A _5901_/A vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__nor2_1
X_4806_ _4685_/X _4805_/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7291_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6242__A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5786_ _5788_/B _6799_/A _5785_/B _5782_/X vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4737_ hold344/X _4529_/X _4745_/S vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7525_ _7534_/CLK _7525_/D vssd1 vssd1 vccd1 vccd1 _7525_/Q sky130_fd_sc_hd__dfxtp_2
X_7456_ _7477_/CLK _7456_/D vssd1 vssd1 vccd1 vccd1 _7456_/Q sky130_fd_sc_hd__dfxtp_1
X_4668_ _7378_/Q _7306_/Q _7298_/Q _7290_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4668_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6896__B _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6407_ hold140/X _6415_/A _6356_/B hold601/X vssd1 vssd1 vccd1 vccd1 _6407_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5702__A1 _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5292__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7387_ _7403_/CLK _7387_/D vssd1 vssd1 vccd1 vccd1 _7387_/Q sky130_fd_sc_hd__dfxtp_1
X_4599_ _3668_/Y _4598_/X _4595_/X vssd1 vssd1 vccd1 vccd1 _4601_/C sky130_fd_sc_hd__a21oi_4
XANTENNA__5702__B2 _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4910__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6338_ _6338_/A _7041_/A vssd1 vssd1 vccd1 vccd1 _7074_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6269_ _6276_/B _7096_/A _6238_/X vssd1 vssd1 vccd1 vccd1 _7137_/B sky130_fd_sc_hd__a21o_1
XANTENNA__7207__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4441__A1 _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__B1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3942__C _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4680__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3970_ _5974_/C _3970_/B _4267_/C _4001_/D vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__and4b_1
XFILLER_0_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5377__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4983__A2 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6062__A _6356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5640_ _5640_/A _5640_/B vssd1 vssd1 vccd1 vccd1 _5640_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4196__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5571_ _5571_/A _5571_/B vssd1 vssd1 vccd1 vccd1 _5571_/X sky130_fd_sc_hd__or2_2
XFILLER_0_86_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7310_ _7446_/CLK _7310_/D vssd1 vssd1 vccd1 vccd1 _7310_/Q sky130_fd_sc_hd__dfxtp_1
X_4522_ _4667_/B _4522_/B vssd1 vssd1 vccd1 vccd1 _4522_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7134__B1 _7558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 _4775_/X vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _7267_/Q vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _7608_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4460_/B vssd1 vssd1 vccd1 vccd1 _4453_/Y sky130_fd_sc_hd__inv_2
X_7241_ _4063_/X hold254/X _7241_/S vssd1 vssd1 vccd1 vccd1 _7241_/X sky130_fd_sc_hd__mux2_1
Xhold259 _5202_/X vssd1 vssd1 vccd1 vccd1 _7390_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _7476_/Q vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _7201_/X vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ _4103_/A _5034_/B _4382_/X _4383_/Y _4162_/B vssd1 vssd1 vccd1 vccd1 _4384_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4310__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7172_ _6326_/C _6377_/X _7230_/A _7230_/B vssd1 vssd1 vccd1 vccd1 _7172_/X sky130_fd_sc_hd__o2bb2a_1
X_6123_ _7236_/B1 _6123_/B vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__and2b_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _7347_/Q _6356_/B _6053_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5448__B1 _5452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4346__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5005_ _5001_/X _5004_/X _4976_/B vssd1 vssd1 vccd1 vccd1 _5005_/Y sky130_fd_sc_hd__a21oi_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4671__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A _7453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6956_ _6938_/X _6955_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6956_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4423__A1 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5907_ _5933_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _5907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6887_ _6887_/A _6887_/B vssd1 vssd1 vccd1 vccd1 _6887_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5838_ _5838_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4187__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5769_ _5769_/A _5769_/B vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__and2_1
XANTENNA__4282__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7508_ _7536_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7439_ _7439_/CLK _7439_/D vssd1 vssd1 vccd1 vccd1 _7439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4337__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3848__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4414__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5611__B1 _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5197__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6167__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6167__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4178__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4130__A _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output74_A _7523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4328__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__A _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6810_ _6865_/A _6865_/B vssd1 vssd1 vccd1 vccd1 _6811_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3839__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4008__C _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5602__B1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4500__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6741_ _6796_/A _6740_/B _6737_/X vssd1 vssd1 vccd1 vccd1 _6789_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3953_ hold97/A _3643_/Y _4036_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__a211o_1
X_3884_ _7322_/Q _7338_/Q _7314_/Q _7450_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3884_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6158__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6158__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6672_ _6673_/A _6673_/B vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5623_ _6445_/A _5580_/B _5576_/B _6793_/A vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5554_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4505_ _4999_/B _4601_/A vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__nor2_1
X_5485_ split8/A _5500_/B vssd1 vssd1 vccd1 vccd1 _5495_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4436_ _4394_/X _4435_/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7251_/D sky130_fd_sc_hd__mux2_1
X_7224_ hold179/X _4589_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7621_/D sky130_fd_sc_hd__mux2_1
X_7155_ _7154_/X _4394_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7592_/D sky130_fd_sc_hd__mux2_1
X_4367_ _4367_/A _5032_/C vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6106_ _6106_/A vssd1 vssd1 vccd1 vccd1 _6106_/Y sky130_fd_sc_hd__inv_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4360_/B _4298_/B vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__and2b_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _6887_/Y _7085_/Y split4/X vssd1 vssd1 vccd1 vccd1 _7086_/Y sky130_fd_sc_hd__a21oi_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4186__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6037_ _6025_/Y _6034_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__o21a_1
Xrebuffer30 split1/A vssd1 vssd1 vccd1 vccd1 _5528_/S sky130_fd_sc_hd__buf_6
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4914__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _6939_/A _6939_/B vssd1 vssd1 vccd1 vccd1 _6940_/B sky130_fd_sc_hd__xnor2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6149__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6149__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4255__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold590 _5210_/X vssd1 vssd1 vccd1 vccd1 _7394_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4635__A1 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4824__S _4824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7200__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6388__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6605__A _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3948__B _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4125__A _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5270_ hold488/X _4849_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _7420_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6312__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4221_ _4401_/S _4221_/B vssd1 vssd1 vccd1 vccd1 _4221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5390__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4152_ _4964_/S _4789_/C vssd1 vssd1 vccd1 vccd1 _4750_/B sky130_fd_sc_hd__nand2_1
X_4083_ _4084_/A _5985_/A _4121_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__and4_4
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4019__B _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4734__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6918__A3 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5051__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4985_ _4985_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4985_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__6234__B _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3936_ _3939_/A _6093_/A vssd1 vssd1 vccd1 vccd1 _3937_/B sky130_fd_sc_hd__or2_1
X_6724_ _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6724_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout143_A _6718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3867_ _3827_/S _3865_/X _3866_/Y _3861_/Y vssd1 vssd1 vccd1 vccd1 _4862_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6655_ _6583_/B _6540_/B _6540_/C vssd1 vssd1 vccd1 vccd1 _6656_/B sky130_fd_sc_hd__a21o_1
X_3798_ _3931_/S _3798_/B vssd1 vssd1 vccd1 vccd1 _3798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5606_ hold76/A _6808_/B vssd1 vssd1 vccd1 vccd1 _5607_/B sky130_fd_sc_hd__nand2_1
X_6586_ _6629_/A _6586_/B _6586_/C vssd1 vssd1 vccd1 vccd1 _6621_/A sky130_fd_sc_hd__and3_1
XANTENNA__6250__A _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5537_ _5537_/A vssd1 vssd1 vccd1 vccd1 _5537_/Y sky130_fd_sc_hd__inv_2
X_7207_ hold188/X _4679_/X _7209_/S vssd1 vssd1 vccd1 vccd1 _7207_/X sky130_fd_sc_hd__mux2_1
X_5468_ _5454_/A _5454_/B _5454_/C _5466_/A vssd1 vssd1 vccd1 vccd1 _5471_/C sky130_fd_sc_hd__a31o_4
X_5399_ hold439/X _4483_/X _5409_/S vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__mux2_1
X_4419_ _7373_/Q _7301_/Q _7293_/Q _7285_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4419_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4865__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7138_ _6235_/A _6827_/A _3946_/Y _7078_/A _7123_/X vssd1 vssd1 vccd1 vccd1 _7138_/X
+ sky130_fd_sc_hd__a311o_1
X_7069_ _7069_/A _7069_/B _7069_/C vssd1 vssd1 vccd1 vccd1 _7073_/B sky130_fd_sc_hd__and3_1
XANTENNA__5290__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3768__B _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 custom_settings[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3784__A _5811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4819__S _4823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4400__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5504__A _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4856__A1 _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5281__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _7212_/B _7151_/B _5376_/C vssd1 vssd1 vccd1 vccd1 _4785_/S sky130_fd_sc_hd__and3_4
XANTENNA__4792__A0 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5385__S _5391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3721_ _7230_/A _3780_/A vssd1 vssd1 vccd1 vccd1 _3721_/Y sky130_fd_sc_hd__nand2_1
X_6440_ _6532_/A _6476_/B vssd1 vssd1 vccd1 vccd1 _6441_/A sky130_fd_sc_hd__nor2_1
X_3652_ _3652_/A vssd1 vssd1 vccd1 vccd1 _3652_/Y sky130_fd_sc_hd__inv_2
X_6371_ _6373_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _7566_/D sky130_fd_sc_hd__and2_1
X_5322_ _7212_/A _5322_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5337_/S sky130_fd_sc_hd__and3_4
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5253_ hold286/X _4887_/X _5265_/S vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5184_ _4897_/X hold357/X _5194_/S vssd1 vssd1 vccd1 vccd1 _5184_/X sky130_fd_sc_hd__mux2_1
X_4204_ _7423_/Q _7355_/Q _7347_/Q _7327_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4204_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4135_ _4850_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4982_/A sky130_fd_sc_hd__and2_4
XANTENNA__5272__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4066_ _5810_/A _5804_/B _5979_/B _4065_/X vssd1 vssd1 vccd1 vccd1 _4066_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6245__A _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7013__A2 _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6221__B1 _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4968_ _6075_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _4968_/X sky130_fd_sc_hd__and2_1
X_3919_ _3918_/X _3912_/X _3827_/S _3917_/Y vssd1 vssd1 vccd1 vccd1 _6130_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4899_ _4166_/B hold667/X _4964_/S vssd1 vssd1 vccd1 vccd1 _4899_/X sky130_fd_sc_hd__a21o_1
X_6707_ _6648_/A _6642_/B _6605_/X vssd1 vssd1 vccd1 vccd1 _6708_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_19_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6638_ _6694_/A _6694_/B _6699_/B _6636_/X vssd1 vssd1 vccd1 vccd1 _6670_/A sky130_fd_sc_hd__a31o_4
XFILLER_0_34_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold103_A _7580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6569_ _6575_/A _6569_/B _6569_/C vssd1 vssd1 vccd1 vccd1 _6570_/B sky130_fd_sc_hd__nand3_1
XANTENNA__6288__B1 _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4838__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 hold654/X vssd1 vssd1 vccd1 vccd1 _6962_/A sky130_fd_sc_hd__buf_6
XANTENNA__6139__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout163 hold664/X vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__buf_8
Xfanout141 _6844_/A vssd1 vssd1 vccd1 vccd1 _6532_/A sky130_fd_sc_hd__clkbuf_8
Xfanout152 _7574_/Q vssd1 vssd1 vccd1 vccd1 _5818_/B sky130_fd_sc_hd__clkbuf_8
Xfanout174 hold665/X vssd1 vssd1 vccd1 vccd1 _6427_/B sky130_fd_sc_hd__buf_6
Xfanout185 _7362_/Q vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__buf_6
Xfanout196 _4421_/S vssd1 vssd1 vccd1 vccd1 _4710_/S sky130_fd_sc_hd__buf_8
XANTENNA__5263__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4449__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__A1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4403__A _4407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4829__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3961__B _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5254__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5888__B _5918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _5940_/A _5940_/B vssd1 vssd1 vccd1 vccd1 _5941_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7610_ _7618_/CLK _7610_/D vssd1 vssd1 vccd1 vccd1 _7610_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5006__A1 _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5871_ _5904_/A _5869_/Y _5816_/X _5820_/A vssd1 vssd1 vccd1 vccd1 _5872_/C sky130_fd_sc_hd__a211o_1
X_4822_ _4821_/X _4637_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7298_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4753_ hold352/X _4385_/X _4767_/S vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__mux2_1
X_7541_ _7541_/CLK hold53/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7472_ _7475_/CLK _7472_/D vssd1 vssd1 vccd1 vccd1 _7472_/Q sky130_fd_sc_hd__dfxtp_1
X_3704_ _6326_/B _4035_/A vssd1 vssd1 vccd1 vccd1 _3780_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4684_ _3933_/Y _4107_/Y _4683_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _4685_/B sky130_fd_sc_hd__o2bb2a_1
X_6423_ _6423_/A _6427_/A vssd1 vssd1 vccd1 vccd1 _6423_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5190__A0 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3635_ _6872_/A vssd1 vssd1 vccd1 vccd1 _6874_/A sky130_fd_sc_hd__inv_2
XANTENNA_fanout106_A _5452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6354_ _7230_/A _7070_/A vssd1 vssd1 vccd1 vccd1 _6354_/Y sky130_fd_sc_hd__nor2_1
X_5305_ hold399/X _4864_/X _5319_/S vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__mux2_1
X_6285_ _6939_/A _6949_/B vssd1 vssd1 vccd1 vccd1 _6287_/B sky130_fd_sc_hd__and2_1
X_5236_ _4871_/Y hold540/X _5248_/S vssd1 vssd1 vccd1 vccd1 _7405_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ hold222/X _4529_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5245__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5098_ _5097_/X _4849_/X _5112_/S vssd1 vssd1 vccd1 vccd1 _7344_/D sky130_fd_sc_hd__mux2_1
X_4118_ _4953_/A _4118_/B _4118_/C _5008_/A vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__or4_2
X_4049_ _7244_/A input8/X _4039_/C _4048_/X vssd1 vssd1 vccd1 vccd1 _4049_/X sky130_fd_sc_hd__a22o_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6984__A1 _4030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4832__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3956__B _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7161__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 _5401_/X vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _7441_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5357__C_N _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A vssd1 vssd1 vccd1 vccd1 _6070_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5475__A1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4278__A2 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _3937_/Y _4106_/X _5020_/X _4083_/X vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__o22a_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5227__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5411__B _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4986__A0 _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6975__A1 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6972_ _6972_/A _6972_/B vssd1 vssd1 vccd1 vccd1 _6972_/X sky130_fd_sc_hd__or2_1
X_5923_ _5923_/A _5923_/B _5923_/C vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__nor3_1
XANTENNA__4742__S _4746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3884__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5854_ _6516_/A _7123_/A _5854_/C _6702_/A vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__and4_1
X_4805_ hold456/X _4719_/Y _4805_/S vssd1 vssd1 vccd1 vccd1 _4805_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5139__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5785_ _5782_/X _5785_/B vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__and2b_1
XANTENNA__6242__B _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7524_ _7534_/CLK _7524_/D vssd1 vssd1 vccd1 vccd1 _7524_/Q sky130_fd_sc_hd__dfxtp_2
X_4736_ hold372/X _4443_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7262_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7152__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3882__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4667_ _4666_/X _4667_/B vssd1 vssd1 vccd1 vccd1 _4667_/Y sky130_fd_sc_hd__nand2b_1
X_7455_ _7569_/CLK hold93/X vssd1 vssd1 vccd1 vccd1 _7455_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7386_ _7403_/CLK _7386_/D vssd1 vssd1 vccd1 vccd1 _7386_/Q sky130_fd_sc_hd__dfxtp_1
X_6406_ _6405_/X _6882_/A _6414_/S vssd1 vssd1 vccd1 vccd1 _7577_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4598_ _4596_/X _4597_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4598_/X sky130_fd_sc_hd__mux2_1
X_6337_ _7040_/A _7040_/C _7040_/B vssd1 vssd1 vccd1 vccd1 _7041_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6268_ _6242_/X _7072_/A _6240_/X vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__a21o_1
X_5219_ hold368/X _4912_/Y _5229_/S vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__mux2_1
X_6199_ _3648_/Y _3649_/Y _6207_/S vssd1 vssd1 vccd1 vccd1 _6199_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5218__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6417__B _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4218__A _4955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6966__B2 _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6966__A1 _3716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4441__A2 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit24 _6716_/A vssd1 vssd1 vccd1 vccd1 _5918_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__B2 _7547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7143__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__A0 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3942__D _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7203__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5209__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6957__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3686__B _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4196__A1 _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _6431_/A _5571_/A _5570_/C vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__nor3_1
X_4521_ _4520_/X _4519_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__mux2_1
X_4452_ _3668_/Y _4451_/X _4448_/X vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__a21oi_4
Xhold216 _7292_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _7195_/X vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
X_7240_ hold604/X hold601/X _7241_/S vssd1 vssd1 vccd1 vccd1 _7529_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold238 _7438_/Q vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _5377_/X vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _7620_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
X_4383_ _4383_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4383_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7171_ _7171_/A _7233_/B _7171_/C vssd1 vssd1 vccd1 vccd1 _7171_/X sky130_fd_sc_hd__or3_1
X_6122_ _6121_/X hold84/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__mux2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4737__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6053_ _6356_/B _6053_/B vssd1 vssd1 vccd1 vccd1 _6053_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6518__A _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _4238_/A _4953_/Y _4957_/X _5003_/Y vssd1 vssd1 vccd1 vccd1 _5004_/X sky130_fd_sc_hd__o22a_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4038__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6955_ _4030_/B _6953_/X _6954_/X vssd1 vssd1 vccd1 vccd1 _6955_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__6253__A _6738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _5930_/A _5905_/C _5905_/A vssd1 vssd1 vccd1 vccd1 _5907_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6886_ _7030_/A _7030_/B _7062_/A _6883_/X vssd1 vssd1 vccd1 vccd1 _7085_/B sky130_fd_sc_hd__a31oi_2
XFILLER_0_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5837_ _5852_/B _5837_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4187__A1 _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5768_ _5768_/A _5768_/B vssd1 vssd1 vccd1 vccd1 _5769_/B sky130_fd_sc_hd__or2_1
XANTENNA__4282__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4719_ _4719_/A _4719_/B vssd1 vssd1 vccd1 vccd1 _4719_/Y sky130_fd_sc_hd__nor2_8
X_7507_ _7538_/CLK hold45/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7438_ _7439_/CLK _7438_/D vssd1 vssd1 vccd1 vccd1 _7438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5699_ _6581_/A _6742_/A _5698_/C vssd1 vssd1 vccd1 vccd1 _5700_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_49_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7537_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7369_ _7418_/CLK _7369_/D vssd1 vssd1 vccd1 vccd1 _7369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4895__C1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3793__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_A _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4647__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3848__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4414__A2 _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4178__A1 _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7116__A1 _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4350__A1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output67_A _7556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6338__A _6338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7052__B1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5388__S _5392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3839__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ _6737_/X _6740_/B vssd1 vssd1 vccd1 vccd1 _6796_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3952_ _7545_/Q _5879_/A _7020_/A _7547_/Q vssd1 vssd1 vccd1 vccd1 _3954_/C sky130_fd_sc_hd__a22o_1
X_3883_ _7402_/Q _7394_/Q _7370_/Q _7386_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3883_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6671_ _6639_/B _6670_/X _6709_/S vssd1 vssd1 vccd1 vccd1 _6673_/B sky130_fd_sc_hd__mux2_2
XANTENNA__5366__A0 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5622_ _5622_/A _5622_/B _5621_/A vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5553_ _5553_/A _5553_/B _5553_/C vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__nand3_1
XANTENNA__7107__A1 _6084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4504_ _4508_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__or2_1
XFILLER_0_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4321__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5484_ _5477_/X _5479_/Y _5480_/Y vssd1 vssd1 vccd1 vccd1 _5500_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4435_ hold534/X _4434_/Y _4720_/S vssd1 vssd1 vccd1 vccd1 _4435_/X sky130_fd_sc_hd__mux2_1
X_7223_ hold178/X _4629_/X _7227_/S vssd1 vssd1 vccd1 vccd1 _7223_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6330__A2 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7154_ hold458/X _4434_/Y _7166_/S vssd1 vssd1 vccd1 vccd1 _7154_/X sky130_fd_sc_hd__mux2_1
X_4366_ _4474_/A _6080_/B vssd1 vssd1 vccd1 vccd1 _5032_/C sky130_fd_sc_hd__or2_1
XFILLER_0_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4467__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6105_ _4407_/B _6107_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__mux2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4296_/X _4295_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4298_/B sky130_fd_sc_hd__mux2_1
XANTENNA__6094__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6094__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6248__A _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _7085_/A _7085_/B vssd1 vssd1 vccd1 vccd1 _7085_/Y sky130_fd_sc_hd__nand2_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _7345_/Q _6162_/A _6035_/Y _6922_/C vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__a211o_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer31 _5585_/A vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__clkbuf_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5298__S _5302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _6931_/X _6933_/X _6937_/X _6326_/C vssd1 vssd1 vccd1 vccd1 _6938_/X sky130_fd_sc_hd__o31a_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6869_ _6869_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6880_/B sky130_fd_sc_hd__and2_1
XFILLER_0_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4930__S _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4255__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4580__A1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold580 _7333_/Q vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 _7554_/Q vssd1 vssd1 vccd1 vccd1 _3733_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6085__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6085__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4191__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5596__B1 _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5348__A0 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4840__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6312__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4220_ _7441_/Q _7433_/Q _7417_/Q _7409_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4221_/B sky130_fd_sc_hd__mux4_1
XANTENNA__6076__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4151_ _7529_/Q _4150_/X _4162_/B vssd1 vssd1 vccd1 vccd1 _4789_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4087__A0 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6076__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4082_ _4084_/A _4280_/B _4290_/D vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__or3_4
XANTENNA__3834__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5036__C1 _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4984_ _4311_/B _4984_/B vssd1 vssd1 vccd1 vccd1 _4985_/B sky130_fd_sc_hd__and2b_1
X_3935_ _3935_/A _3935_/B vssd1 vssd1 vccd1 vccd1 _3935_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6723_ _6680_/Y _6723_/B vssd1 vssd1 vccd1 vccd1 _6724_/B sky130_fd_sc_hd__nand2b_1
X_6654_ _6600_/A _6601_/Y _6544_/A vssd1 vssd1 vccd1 vccd1 _6764_/A sky130_fd_sc_hd__a21oi_1
X_3866_ _3886_/S _3862_/X _7363_/Q vssd1 vssd1 vccd1 vccd1 _3866_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5605_ _6518_/A _5605_/B _5605_/C vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3797_ _7281_/Q _7596_/Q _7265_/Q _7489_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3798_/B sky130_fd_sc_hd__mux4_1
XANTENNA__6250__B _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6585_ _6585_/A vssd1 vssd1 vccd1 vccd1 _6585_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5536_ _5536_/A _5536_/B vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__or2_1
X_5467_ _5460_/A _5466_/Y _5467_/B1 _5454_/B _5454_/A vssd1 vssd1 vccd1 vccd1 _5471_/B
+ sky130_fd_sc_hd__o2111ai_4
X_4418_ _4416_/X _4417_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__mux2_1
X_7206_ hold351/X _4589_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7613_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3890__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5398_ _4394_/X _5397_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7485_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4349_ _4349_/A _4861_/B vssd1 vssd1 vccd1 vccd1 _4349_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6067__A1 _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7137_ _7137_/A _7137_/B vssd1 vssd1 vccd1 vccd1 _7137_/X sky130_fd_sc_hd__or2_1
XANTENNA__6067__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7068_ _7090_/A split9/X _7067_/X _5970_/A vssd1 vssd1 vccd1 vccd1 _7068_/X sky130_fd_sc_hd__o211a_1
X_6019_ _7168_/A _6349_/A _7168_/B _7231_/A vssd1 vssd1 vccd1 vccd1 _6020_/B sky130_fd_sc_hd__or4b_1
XANTENNA__7016__B1 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3768__C _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4896__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4400__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6058__A1 _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6058__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4069__A0 hold97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3911__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3959__B _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _5805_/A _4035_/A _4036_/A vssd1 vssd1 vccd1 vccd1 _6333_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__3975__A _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3694__B _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ hold84/X vssd1 vssd1 vccd1 vccd1 _3651_/Y sky130_fd_sc_hd__inv_2
X_6370_ _7529_/Q hold140/X _6372_/S vssd1 vssd1 vccd1 vccd1 _6370_/X sky130_fd_sc_hd__mux2_1
X_5321_ _5393_/A _5321_/B _5159_/C vssd1 vssd1 vccd1 vccd1 _5338_/S sky130_fd_sc_hd__or3b_4
XFILLER_0_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5252_ hold235/X _4849_/X _5266_/S vssd1 vssd1 vccd1 vccd1 _7412_/D sky130_fd_sc_hd__mux2_1
X_5183_ hold356/X _4912_/Y _5193_/S vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__mux2_1
X_4203_ _7319_/Q _7335_/Q _7311_/Q _7447_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4203_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6049__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6049__A1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4134_ _5132_/A _7473_/Q _4267_/C _4134_/D vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__nand4_4
XANTENNA__4745__S _4745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ _7555_/Q _4846_/A _4065_/C vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3902__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__B1 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6245__B _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _4971_/B _4942_/B _4942_/Y vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4783__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3918_ _7362_/Q _3913_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _3918_/X sky130_fd_sc_hd__a21o_1
X_4898_ _7344_/Q hold666/X hold633/X vssd1 vssd1 vccd1 vccd1 _4898_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6261__A _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6706_ _6771_/A _6669_/B _6674_/A vssd1 vssd1 vccd1 vccd1 _6706_/X sky130_fd_sc_hd__o21ba_4
X_3849_ _3847_/X _3848_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6637_ _6637_/A _6637_/B vssd1 vssd1 vccd1 vccd1 _6699_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4535__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6568_ _6568_/A _6568_/B vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__and2_1
XFILLER_0_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5519_ _5553_/B _5520_/B _5520_/C vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__a21oi_1
X_6499_ _6471_/B _6521_/D _6521_/A vssd1 vssd1 vccd1 vccd1 _6503_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__5605__A _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout131 _6935_/A vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__clkbuf_8
Xfanout120 hold644/X vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__buf_6
Xfanout153 _6799_/A vssd1 vssd1 vccd1 vccd1 _6742_/A sky130_fd_sc_hd__buf_6
Xfanout142 _7578_/Q vssd1 vssd1 vccd1 vccd1 _6844_/A sky130_fd_sc_hd__buf_6
Xfanout164 _7551_/Q vssd1 vssd1 vccd1 vccd1 _7230_/A sky130_fd_sc_hd__buf_4
Xfanout186 _3896_/S1 vssd1 vssd1 vccd1 vccd1 _3883_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout175 _7455_/Q vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__clkbuf_8
Xfanout197 _7342_/Q vssd1 vssd1 vccd1 vccd1 _4421_/S sky130_fd_sc_hd__buf_8
XFILLER_0_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4449__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4774__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5971__B1 _5952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4122__C _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7206__S _7210_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5250__A _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5870_ _5816_/X _5820_/A _5904_/A _5869_/Y vssd1 vssd1 vccd1 vccd1 _5904_/B sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ hold241/X _4679_/X _4823_/S vssd1 vssd1 vccd1 vccd1 _4821_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5396__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4765__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4752_ _7212_/B _7212_/C _5376_/C vssd1 vssd1 vccd1 vccd1 _4767_/S sky130_fd_sc_hd__and3_4
X_7540_ _7581_/CLK _7540_/D vssd1 vssd1 vccd1 vccd1 _7540_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7471_ _7596_/CLK _7471_/D vssd1 vssd1 vccd1 vccd1 _7471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4683_ _6235_/A _4440_/A _4440_/Y _4682_/X vssd1 vssd1 vccd1 vccd1 _4683_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3703_ _4084_/A _4119_/A _5985_/A vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3634_ _6802_/A vssd1 vssd1 vccd1 vccd1 _6738_/A sky130_fd_sc_hd__clkinv_4
X_6422_ hold104/X _6421_/X _6204_/A vssd1 vssd1 vccd1 vccd1 _6422_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6353_ _6374_/A _5811_/B _6351_/A _6351_/B hold616/X vssd1 vssd1 vccd1 vccd1 _6353_/X
+ sky130_fd_sc_hd__a41o_1
X_5304_ _7151_/B _5376_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5319_/S sky130_fd_sc_hd__and3_4
XFILLER_0_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6284_ _7020_/A _6271_/X _6283_/Y _5879_/A vssd1 vssd1 vccd1 vccd1 _6333_/B sky130_fd_sc_hd__a22o_1
X_5235_ hold539/X _4887_/X _5247_/S vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ hold490/X _4443_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7374_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5160__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5097_ _3663_/A _4864_/X _5111_/S vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__mux2_1
X_4117_ _6328_/B _4290_/D vssd1 vssd1 vccd1 vccd1 _4930_/S sky130_fd_sc_hd__or2_4
XANTENNA__6256__A _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4048_ hold97/X _4047_/X _6329_/A vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5999_ _5999_/A hold68/X vssd1 vssd1 vccd1 vccd1 _5999_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4756__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5953__B1 _5810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold213_A _7527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5181__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6166__A _6166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6433__B2 _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6105__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold409 _7383_/Q vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5172__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4358__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5020_ _6235_/A _4945_/B _4918_/Y _5019_/Y vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__o22a_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5411__C _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6971_ _4084_/A _6974_/A _6970_/X _3949_/Y vssd1 vssd1 vccd1 vccd1 _6971_/X sky130_fd_sc_hd__o211a_1
X_5922_ _5922_/A _5922_/B vssd1 vssd1 vccd1 vccd1 _5923_/C sky130_fd_sc_hd__xnor2_1
X_5853_ _6516_/A _5854_/C _6702_/A _7123_/A vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__a22oi_1
XANTENNA__4738__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4804_ _4637_/X _4803_/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7290_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5935__B1 _5952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5784_ _6738_/A _6808_/B _6978_/A vssd1 vssd1 vccd1 vccd1 _5785_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4735_ hold371/X _4483_/X _4745_/S vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7523_ _7538_/CLK _7523_/D vssd1 vssd1 vccd1 vccd1 _7523_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4666_ _4664_/X _4665_/X _4710_/S vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__mux2_1
X_7454_ _7454_/CLK _7454_/D vssd1 vssd1 vccd1 vccd1 _7454_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7385_ _7418_/CLK _7385_/D vssd1 vssd1 vccd1 vccd1 _7385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5163__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4597__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4597_ _7273_/Q _7613_/Q _7605_/Q _7621_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4597_/X sky130_fd_sc_hd__mux4_1
X_6405_ input36/X _6404_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6405_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6360__A0 _7569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6427__C_N _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6336_ _7009_/A _7009_/C _7009_/B vssd1 vssd1 vccd1 vccd1 _7040_/C sky130_fd_sc_hd__a21o_1
X_6267_ _6295_/A _6267_/B vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__nand2_1
X_5218_ hold479/X _4871_/Y _5230_/S vssd1 vssd1 vccd1 vccd1 _7397_/D sky130_fd_sc_hd__mux2_1
X_6198_ _6198_/A _6198_/B vssd1 vssd1 vccd1 vccd1 _7533_/D sky130_fd_sc_hd__nand2_1
X_5149_ hold598/X _4937_/Y _5157_/S vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5623__C1 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xsplit25 _6790_/S vssd1 vssd1 vccd1 vccd1 _6832_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3952__A2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6406__A1 _6882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6957__A2 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4843__S _4843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6624__A _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _7271_/Q _7611_/Q _7603_/Q _7619_/Q _4709_/S0 _4709_/S1 vssd1 vssd1 vccd1
+ vccd1 _4520_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5145__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 _7467_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _4449_/X _4450_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__mux2_1
Xhold217 _4809_/X vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _5309_/X vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _7269_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
X_7170_ _6020_/C _7170_/B _7231_/A vssd1 vssd1 vccd1 vccd1 _7171_/C sky130_fd_sc_hd__nand3b_1
X_4382_ _4383_/A _4383_/B _4986_/S vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__o21a_1
X_6121_ _6427_/B _6119_/X _6120_/Y _4453_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6121_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6052_/A vssd1 vssd1 vccd1 vccd1 _6052_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5003_ _5026_/A _5003_/B vssd1 vssd1 vccd1 vccd1 _5003_/Y sky130_fd_sc_hd__nand2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4038__B _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4753__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6954_ _6039_/A _5804_/C _4029_/Y _6111_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _6954_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout166_A _7551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3877__B _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6253__B _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5905_ _5905_/A _5930_/A _5905_/C vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__and3_1
X_6885_ _7030_/A _7030_/B _7062_/A _6883_/X vssd1 vssd1 vccd1 vccd1 _6887_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5836_ _5852_/A _5834_/Y _5697_/B _5700_/A vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__a211o_1
XANTENNA__5384__A1 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4989__A _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5767_ _5797_/B _5767_/B vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__nand2_1
X_4718_ _4144_/Y _4715_/X _4704_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4719_/B sky130_fd_sc_hd__o211a_2
X_7506_ _7537_/CLK hold47/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7125__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5698_ _6581_/A _6742_/A _5698_/C vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__and3_1
X_7437_ _7449_/CLK _7437_/D vssd1 vssd1 vccd1 vccd1 _7437_/Q sky130_fd_sc_hd__dfxtp_1
X_4649_ _4698_/C vssd1 vssd1 vccd1 vccd1 _4649_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5136__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7368_ _4004_/A _7368_/D vssd1 vssd1 vccd1 vccd1 _7368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3793__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7299_ _7378_/CLK _7299_/D vssd1 vssd1 vccd1 vccd1 _7299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6319_ _6319_/A _6319_/B vssd1 vssd1 vccd1 vccd1 _6993_/B sky130_fd_sc_hd__or2_1
XFILLER_0_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6636__A1 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7418_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6444__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5127__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4130__C _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4838__S _4844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7214__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5523__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit1 split1/A vssd1 vssd1 vccd1 vccd1 split1/X sky130_fd_sc_hd__buf_6
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3978__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6354__A _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3697__B _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3951_ _7546_/Q _7098_/A _3950_/X vssd1 vssd1 vccd1 vccd1 _3954_/B sky130_fd_sc_hd__a21o_1
X_3882_ _3915_/A _3882_/B vssd1 vssd1 vccd1 vccd1 _3882_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6670_ _6670_/A _6670_/B vssd1 vssd1 vccd1 vccd1 _6670_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5621_ _5621_/A _5621_/B _5621_/C _5621_/D vssd1 vssd1 vccd1 vccd1 _5621_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__4602__A _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5552_ _6532_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _5557_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5118__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4503_ _3668_/Y _4502_/X _4499_/X vssd1 vssd1 vccd1 vccd1 _6123_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7107__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5483_ _5458_/Y _5483_/B vssd1 vssd1 vccd1 vccd1 _5489_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7222_ _7221_/X _4538_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7620_/D sky130_fd_sc_hd__mux2_1
X_4434_ _4989_/A _4493_/C _4433_/Y _4431_/X vssd1 vssd1 vccd1 vccd1 _4434_/Y sky130_fd_sc_hd__a31oi_4
X_7153_ hold455/X _4111_/X _7167_/S vssd1 vssd1 vccd1 vccd1 _7591_/D sky130_fd_sc_hd__mux2_1
X_4365_ _4474_/A _6080_/B vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _7025_/A _6926_/Y _7082_/Y _7083_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7588_/D
+ sky130_fd_sc_hd__o221a_1
X_6104_ _6103_/X hold74/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__mux2_1
X_4296_ _7425_/Q _7357_/Q _7349_/Q _7329_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4296_/X sky130_fd_sc_hd__mux4_1
X_6035_ _6162_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6035_/Y sky130_fd_sc_hd__nor2_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6248__B _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer21 _5605_/C vssd1 vssd1 vccd1 vccd1 _5601_/B sky130_fd_sc_hd__clkbuf_1
Xrebuffer10 _6463_/S vssd1 vssd1 vccd1 vccd1 _6432_/S sky130_fd_sc_hd__buf_1
XFILLER_0_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4483__S _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _7025_/A _6922_/B _7023_/A _6934_/Y _6952_/B vssd1 vssd1 vccd1 vccd1 _6937_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6868_ _6807_/B _6891_/B _6866_/X _6871_/A vssd1 vssd1 vccd1 vccd1 _6868_/Y sky130_fd_sc_hd__o211ai_2
X_5819_ _5818_/C _5818_/D _6298_/A _5504_/A vssd1 vssd1 vccd1 vccd1 _5820_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3827__S _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6203__S _6207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6799_ _6799_/A _6799_/B vssd1 vssd1 vccd1 vccd1 _6813_/B sky130_fd_sc_hd__and2_1
XANTENNA__5109__A1 _5015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold581 _5081_/X vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 _7307_/Q vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 hold97/A vssd1 vssd1 vccd1 vccd1 _4035_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4191__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3798__A _3931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7034__B2 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7034__A1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7209__S _7209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6113__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4859__B1 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _7570_/Q input15/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4150_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4706__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4087__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4081_ _4081_/A _4279_/C vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__nand2_8
XANTENNA__3834__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5399__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6084__A _6084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4673__A_N _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4983_ input26/X _5031_/S _4162_/B vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3934_ _3934_/A _6120_/A vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__or2_1
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6722_ _6857_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6781_/A sky130_fd_sc_hd__xnor2_4
X_3865_ _3863_/X _3864_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6653_ _6601_/Y split9/X _6651_/X _6652_/Y vssd1 vssd1 vccd1 vccd1 _6653_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5428__A _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5604_ _5604_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _6462_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3796_ _3827_/S _3794_/X _3795_/Y _3791_/Y vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout129_A _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6584_ _6586_/B _6586_/C vssd1 vssd1 vccd1 vccd1 _6585_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5535_ _5535_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _5536_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ _5466_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _5466_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _7477_/Q _7465_/Q _7457_/Q _7251_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4417_/X sky130_fd_sc_hd__mux4_1
X_7205_ hold350/X _4629_/X _7209_/S vssd1 vssd1 vccd1 vccd1 _7205_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5511__A1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5397_ hold441/X _4434_/Y _5409_/S vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__mux2_1
X_4348_ _4360_/B _4347_/X _4344_/Y vssd1 vssd1 vccd1 vccd1 _4861_/B sky130_fd_sc_hd__o21ai_2
X_7136_ _5800_/B _5747_/X _5798_/A _5798_/Y vssd1 vssd1 vccd1 vccd1 _7136_/X sky130_fd_sc_hd__o211a_1
X_4279_ _6900_/A _5804_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__and3_4
X_7067_ _7065_/X _7066_/X _6900_/A vssd1 vssd1 vccd1 vccd1 _7067_/X sky130_fd_sc_hd__a21o_1
X_6018_ _3988_/A _7230_/B _6417_/B vssd1 vssd1 vccd1 vccd1 _6349_/A sky130_fd_sc_hd__a21oi_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__D _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6722__A _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7593_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4069__A1 _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3911__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4152__A _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3650_ _3650_/A vssd1 vssd1 vccd1 vccd1 _3650_/Y sky130_fd_sc_hd__inv_2
Xrebuffer1 _5454_/C vssd1 vssd1 vccd1 vccd1 _5467_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5320_ hold187/X _5022_/X _5320_/S vssd1 vssd1 vccd1 vccd1 _7443_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5251_ hold234/X _4864_/X _5265_/S vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4202_ _7399_/Q _7391_/Q _7367_/Q _7383_/Q _4255_/S0 _4255_/S1 vssd1 vssd1 vccd1
+ vccd1 _4202_/X sky130_fd_sc_hd__mux4_1
X_5182_ _4871_/Y hold563/X _5194_/S vssd1 vssd1 vccd1 vccd1 _7381_/D sky130_fd_sc_hd__mux2_1
XANTENNA__7246__A1 hold66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4133_ _5132_/A _7473_/Q _4267_/C _4134_/D vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__and4_4
XANTENNA__6807__A _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4064_ _4063_/X hold254/X _7241_/S vssd1 vssd1 vccd1 vccd1 _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3902__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5009__B1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4761__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ hold170/X _4947_/X _5040_/S vssd1 vssd1 vccd1 vccd1 _7312_/D sky130_fd_sc_hd__mux2_1
X_6705_ _6719_/A _6719_/B _6714_/A _6704_/X vssd1 vssd1 vccd1 vccd1 _6751_/B sky130_fd_sc_hd__a31o_4
XFILLER_0_104_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3917_ _3931_/S _3916_/X _3915_/X vssd1 vssd1 vccd1 vccd1 _3917_/Y sky130_fd_sc_hd__a21oi_1
X_4897_ _5022_/A _4897_/B _4897_/C vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__or3_4
XANTENNA__6261__B _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3848_ _7423_/Q _7355_/Q _7347_/Q _7327_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3848_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4062__A _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6636_ _6869_/A _6637_/B _6635_/X vssd1 vssd1 vccd1 vccd1 _6636_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4535__A2 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6567_ _6567_/A vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__inv_2
X_3779_ _7559_/Q _3780_/A _7123_/C _4084_/A vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__a31o_1
X_5518_ _5488_/X _5493_/A _5554_/A _5517_/X vssd1 vssd1 vccd1 vccd1 split1/A sky130_fd_sc_hd__a31oi_4
XFILLER_0_42_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6498_ _6498_/A _6498_/B vssd1 vssd1 vccd1 vccd1 _6498_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4299__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5449_ _6568_/A split8/A vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout110 _6808_/B vssd1 vssd1 vccd1 vccd1 _6683_/B sky130_fd_sc_hd__clkbuf_8
Xfanout121 _7590_/Q vssd1 vssd1 vccd1 vccd1 _6516_/A sky130_fd_sc_hd__buf_4
XANTENNA__5248__A0 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _6096_/A vssd1 vssd1 vccd1 vccd1 _5024_/S sky130_fd_sc_hd__buf_4
Xfanout132 hold657/X vssd1 vssd1 vccd1 vccd1 _6935_/A sky130_fd_sc_hd__buf_4
XANTENNA__6717__A _6718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 _7574_/Q vssd1 vssd1 vccd1 vccd1 _6799_/A sky130_fd_sc_hd__buf_8
Xfanout143 _6718_/A vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__buf_8
X_7119_ _7137_/A _6309_/Y _6910_/A vssd1 vssd1 vccd1 vccd1 _7119_/Y sky130_fd_sc_hd__a21oi_1
Xfanout198 _4369_/S1 vssd1 vssd1 vccd1 vccd1 _4371_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout176 _7454_/Q vssd1 vssd1 vccd1 vccd1 _4688_/S sky130_fd_sc_hd__buf_6
Xfanout187 _7361_/Q vssd1 vssd1 vccd1 vccd1 _3896_/S1 sky130_fd_sc_hd__buf_6
XANTENNA__5340__B _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6996__B1 _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5971__A1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7173__B1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4700__A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7228__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7222__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4147__A _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3896__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4581__S _4720_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4820_ hold247/X _4589_/X _4824_/S vssd1 vssd1 vccd1 vccd1 _7297_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3986__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4751_ _4751_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _5376_/C sky130_fd_sc_hd__nor2_4
XFILLER_0_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7470_ _7596_/CLK _7470_/D vssd1 vssd1 vccd1 vccd1 _7470_/Q sky130_fd_sc_hd__dfxtp_1
X_4682_ _6166_/A _4682_/B vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4711__A_N _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3702_ _4084_/A _4119_/A _5985_/A vssd1 vssd1 vccd1 vccd1 _3702_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_71_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3633_ _6690_/A vssd1 vssd1 vccd1 vccd1 _6691_/A sky130_fd_sc_hd__inv_2
X_6421_ _6427_/B _6421_/B _6427_/A vssd1 vssd1 vccd1 vccd1 _6421_/X sky130_fd_sc_hd__or3_1
XFILLER_0_31_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6352_ _3744_/A _6351_/Y _7244_/A vssd1 vssd1 vccd1 vccd1 _6352_/X sky130_fd_sc_hd__a21o_1
X_5303_ _7150_/B _5375_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5320_/S sky130_fd_sc_hd__and3_4
XFILLER_0_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6283_ _6974_/C _6282_/X _6271_/X vssd1 vssd1 vccd1 vccd1 _6283_/Y sky130_fd_sc_hd__o21ai_1
X_5234_ _4849_/X hold544/X _5248_/S vssd1 vssd1 vccd1 vccd1 _7404_/D sky130_fd_sc_hd__mux2_1
X_5165_ hold489/X _4483_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4756__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7219__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4150__A0 _7570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5441__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4116_ _6328_/B _4290_/D vssd1 vssd1 vccd1 vccd1 _4116_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5096_ _7176_/B _7212_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5111_/S sky130_fd_sc_hd__and3_4
XANTENNA__6256__B _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4047_ hold66/X _6793_/A _6023_/S vssd1 vssd1 vccd1 vccd1 _4047_/X sky130_fd_sc_hd__mux2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5402__A0 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6272__A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5998_ _5998_/A hold74/X vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__xor2_1
X_4949_ _4977_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__or2_1
XANTENNA__4504__B _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5953__A1 _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6619_ _6619_/A _6619_/B vssd1 vssd1 vccd1 vccd1 _6619_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6902__B1 _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7599_ _7599_/CLK _7599_/D vssd1 vssd1 vccd1 vccd1 _7599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4666__S _4710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6166__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5641__B1 _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7217__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4380__B1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4227__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6121__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4358__S1 _4369_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6121__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4683__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6970_ _6871_/B split4/X _6969_/Y _7043_/S vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4435__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3869__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _5913_/A _5913_/B _5922_/B vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5200__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5852_ _5852_/A _5852_/B vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__nand2_1
X_4803_ hold406/X _4679_/X _4805_/S vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5935__A1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5783_ _5788_/B _6799_/A vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__nand2_1
X_4734_ _4733_/X _4394_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7261_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6820__A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7522_ _7534_/CLK _7522_/D vssd1 vssd1 vccd1 vccd1 _7522_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _7482_/Q _7470_/Q _7462_/Q _7256_/Q _7340_/Q _7341_/Q vssd1 vssd1 vccd1 vccd1
+ _4665_/X sky130_fd_sc_hd__mux4_1
X_7453_ _7453_/CLK _7453_/D vssd1 vssd1 vccd1 vccd1 _7453_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7384_ _4004_/A _7384_/D vssd1 vssd1 vccd1 vccd1 _7384_/Q sky130_fd_sc_hd__dfxtp_1
X_4596_ _7377_/Q _7305_/Q _7297_/Q _7289_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4596_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4597__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4340__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6404_ _7025_/A _6383_/Y _6403_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6404_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout209_A _6345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4910__A2 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6335_ _6978_/A _6978_/C _6978_/B vssd1 vssd1 vccd1 vccd1 _7009_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6112__A1 _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6112__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6266_ _6249_/A _6265_/Y _7019_/A vssd1 vssd1 vccd1 vccd1 _6267_/B sky130_fd_sc_hd__a21o_1
X_5217_ hold478/X _4887_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__mux2_1
X_6197_ _3650_/Y _3651_/Y _6207_/S vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__mux2_1
X_5148_ _4897_/X hold503/X _5158_/S vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__mux2_1
X_5079_ hold359/X _4864_/X _5093_/S vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7098__A _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xsplit26 _6445_/A vssd1 vssd1 vccd1 vccd1 _6611_/A sky130_fd_sc_hd__buf_4
Xsplit15 _6521_/D vssd1 vssd1 vccd1 vccd1 _6509_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4285__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4250__A _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4287__A_N _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6103__B2 _7236_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5090__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4425__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 _5365_/X vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4450_ _7270_/Q _7610_/Q _7602_/Q _7618_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4450_/X sky130_fd_sc_hd__mux4_1
Xhold218 _7264_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _7378_/Q vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ _5011_/A _5012_/A _4376_/Y _4380_/X _5032_/C vssd1 vssd1 vccd1 vccd1 _4477_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6120_ _6120_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4200__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6051_ _4208_/A _6053_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6052_/A sky130_fd_sc_hd__mux2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__B2 _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5002_ _5002_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _5003_/B sky130_fd_sc_hd__or2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__B1 _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6953_ _6872_/A hold610/X _4037_/X _6942_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _6953_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6884_ _6884_/A _6884_/B vssd1 vssd1 vccd1 vccd1 _7062_/A sky130_fd_sc_hd__nor2_1
X_5904_ _5904_/A _5904_/B _5904_/C vssd1 vssd1 vccd1 vccd1 _5905_/C sky130_fd_sc_hd__nand3_1
XANTENNA_fanout159_A _6872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5835_ _5697_/B _5700_/A _5852_/A _5834_/Y vssd1 vssd1 vccd1 vccd1 _5852_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3919__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5766_ _5766_/A _5766_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__or3_1
X_4717_ _7607_/Q _4638_/X _4716_/Y vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7505_ _7582_/CLK hold49/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5697_ _5697_/A _5697_/B vssd1 vssd1 vccd1 vccd1 _5698_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_102_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7436_ _7439_/CLK _7436_/D vssd1 vssd1 vccd1 vccd1 _7436_/Q sky130_fd_sc_hd__dfxtp_1
X_4648_ _3668_/Y _4647_/X _4644_/X vssd1 vssd1 vccd1 vccd1 _4698_/C sky130_fd_sc_hd__a21oi_4
XANTENNA__7125__A3 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7367_ _7396_/CLK _7367_/D vssd1 vssd1 vccd1 vccd1 _7367_/Q sky130_fd_sc_hd__dfxtp_1
X_4579_ _6139_/A _4986_/S _4578_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4579_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__4895__A1 _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5541__C1 _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7298_ _7306_/CLK _7298_/D vssd1 vssd1 vccd1 vccd1 _7298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6097__B1 _6025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6318_ _6264_/A _6318_/B vssd1 vssd1 vccd1 vccd1 _6319_/B sky130_fd_sc_hd__and2b_1
X_6249_ _6249_/A vssd1 vssd1 vccd1 vccd1 _7035_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7046__C1 _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4229__B _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5072__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7541_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6460__A _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4886__A1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5063__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6354__B _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4497__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3950_ _7544_/Q _3705_/X _3949_/Y _7557_/Q vssd1 vssd1 vccd1 vccd1 _3950_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4810__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ _7442_/Q _7434_/Q _7418_/Q _7410_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3882_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5620_ _5622_/B _5620_/B _5620_/C vssd1 vssd1 vccd1 vccd1 _6430_/A sky130_fd_sc_hd__or3_4
X_5551_ split1/X _5550_/X _5488_/B vssd1 vssd1 vccd1 vccd1 _5566_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4502_ _4500_/X _4501_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6315__A1 _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7221_ hold227/X _4580_/X _7227_/S vssd1 vssd1 vccd1 vccd1 _7221_/X sky130_fd_sc_hd__mux2_1
X_5482_ _5482_/A _5482_/B vssd1 vssd1 vccd1 vccd1 _5494_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6315__B2 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4433_ _7351_/Q _7600_/Q _5037_/B _7601_/Q vssd1 vssd1 vccd1 vccd1 _4433_/Y sky130_fd_sc_hd__o31ai_2
XANTENNA__4877__A1 _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7152_ hold454/X _4385_/X _7166_/S vssd1 vssd1 vccd1 vccd1 _7152_/X sky130_fd_sc_hd__mux2_1
X_4364_ _4360_/B _4363_/X _4360_/Y vssd1 vssd1 vccd1 vccd1 _6080_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__4877__B2 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4295_ _7321_/Q _7337_/Q _7313_/Q _7449_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4295_/X sky130_fd_sc_hd__mux4_1
X_6103_ _6101_/X _6102_/Y _4180_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ input36/X _4021_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__a21o_1
X_6034_ _6034_/A vssd1 vssd1 vccd1 vccd1 _6034_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4629__A1 _4989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4764__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer11 _6432_/S vssd1 vssd1 vccd1 vccd1 _5803_/A2 sky130_fd_sc_hd__clkbuf_1
Xrebuffer33 split1/A vssd1 vssd1 vccd1 vccd1 _5532_/S sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 _5561_/X vssd1 vssd1 vccd1 vccd1 _5586_/A2 sky130_fd_sc_hd__clkbuf_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5054__A1 _4973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _6311_/A _6911_/A _7098_/A _6935_/X vssd1 vssd1 vccd1 vccd1 _6952_/B sky130_fd_sc_hd__o211a_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4801__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _6807_/B _6891_/B _6866_/X vssd1 vssd1 vccd1 vccd1 _6871_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6798_ _6790_/S _6796_/Y _6797_/Y vssd1 vssd1 vccd1 vccd1 _6799_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5818_ _6516_/A _5818_/B _5818_/C _5818_/D vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__and4_1
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5749_ _5749_/A _5749_/B vssd1 vssd1 vccd1 vccd1 _5768_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7419_ _7441_/CLK _7419_/D vssd1 vssd1 vccd1 vccd1 _7419_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4939__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold571 _7465_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _7368_/Q vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout91_A _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 _7257_/Q vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _7238_/X vssd1 vssd1 vccd1 vccd1 _7527_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5293__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5045__A1 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4005__C1 _7540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3820__A1_N _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4556__A0 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3835__A1_N _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7225__S _7227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output72_A _7521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4706__S1 _4706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5284__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4080_ _4079_/X hold92/X _7249_/S vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__mux2_1
XANTENNA__5036__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6084__B _6157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4982_ _4982_/A _4982_/B _4982_/C _4976_/X vssd1 vssd1 vccd1 vccd1 _4982_/X sky130_fd_sc_hd__or4b_1
X_3933_ _3933_/A _6166_/A vssd1 vssd1 vccd1 vccd1 _3933_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7570_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6721_ _6857_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6721_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold97_A hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3864_ _7420_/Q _7352_/Q _7344_/Q _7324_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3864_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6652_ _6652_/A split9/X vssd1 vssd1 vccd1 vccd1 _6652_/Y sky130_fd_sc_hd__nor2_1
X_5603_ _5605_/B _5605_/C _6518_/A vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4642__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3795_ _3915_/A _3789_/X _7363_/Q vssd1 vssd1 vccd1 vccd1 _3795_/Y sky130_fd_sc_hd__o21ai_1
X_6583_ _6581_/A _6583_/B _6583_/C vssd1 vssd1 vccd1 vccd1 _6586_/C sky130_fd_sc_hd__nand3b_1
X_5534_ _5534_/A _5818_/B vssd1 vssd1 vccd1 vccd1 _5583_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4759__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5465_ _5504_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__nand2_1
X_4416_ _7277_/Q _7592_/Q _7261_/Q _7485_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4416_/X sky130_fd_sc_hd__mux4_1
X_7204_ _7203_/X _4538_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7612_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3890__C _6084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5444__A _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5396_ _4111_/X hold575/X _5410_/S vssd1 vssd1 vccd1 vccd1 _7484_/D sky130_fd_sc_hd__mux2_1
X_7135_ _7043_/S _6481_/S _7133_/Y _7134_/X _5879_/A vssd1 vssd1 vccd1 vccd1 _7135_/X
+ sky130_fd_sc_hd__o221a_1
X_4347_ _4346_/X _4345_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4347_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5275__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4278_ input29/X _4982_/A _4143_/X _4277_/X vssd1 vssd1 vccd1 vccd1 _4278_/X sky130_fd_sc_hd__a211o_1
X_7066_ _7066_/A _7072_/B _7039_/Y vssd1 vssd1 vccd1 vccd1 _7066_/X sky130_fd_sc_hd__or3b_1
X_6017_ _6417_/B _4007_/A _4007_/B _4033_/B _5985_/Y vssd1 vssd1 vccd1 vccd1 _7231_/A
+ sky130_fd_sc_hd__o32a_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6919_ _7555_/Q _6919_/B vssd1 vssd1 vccd1 vccd1 _6919_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold390 _7417_/Q vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5266__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3959__D _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6913__A _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6124__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5529__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4152__B _4789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7191__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer2 _5589_/X vssd1 vssd1 vccd1 vccd1 _5616_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5250_ _7151_/B _7176_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5265_/S sky130_fd_sc_hd__and3_4
XFILLER_0_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4201_ _4401_/S _4201_/B vssd1 vssd1 vccd1 vccd1 _4201_/Y sky130_fd_sc_hd__nand2_1
X_5181_ hold562/X _4887_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__mux2_1
X_4132_ _4163_/A _4905_/B _4163_/B vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__nor3_4
XANTENNA__5257__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4063_ _4039_/C _4061_/X _4062_/Y input11/X _7244_/A vssd1 vssd1 vccd1 vccd1 _4063_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5203__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5009__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4965_ hold169/X _4964_/X _5039_/S vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire79 wire79/A vssd1 vssd1 vccd1 vccd1 wire79/X sky130_fd_sc_hd__buf_2
XFILLER_0_74_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3916_ _7271_/Q _7611_/Q _7603_/Q _7619_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3916_/X sky130_fd_sc_hd__mux4_1
X_6704_ _6857_/A _6702_/B _6703_/X vssd1 vssd1 vccd1 vccd1 _6704_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4896_ _4946_/A _4896_/B vssd1 vssd1 vccd1 vccd1 _4897_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4615__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3847_ _7319_/Q _7335_/Q _7311_/Q _7447_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3847_/X sky130_fd_sc_hd__mux4_1
XANTENNA__7182__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4062__B _6220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6635_ _6869_/A _6637_/B _6625_/B _6871_/A vssd1 vssd1 vccd1 vccd1 _6635_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ _6568_/A _6568_/B vssd1 vssd1 vccd1 vccd1 _6567_/A sky130_fd_sc_hd__or2_2
X_3778_ _7543_/Q _3780_/B _7123_/C _3712_/B vssd1 vssd1 vccd1 vccd1 _3787_/D sky130_fd_sc_hd__or4b_1
X_5517_ _5556_/A _5488_/B _6710_/A _6532_/A vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6497_ _6529_/B _6505_/B vssd1 vssd1 vccd1 vccd1 _6557_/A sky130_fd_sc_hd__nor2_1
X_5448_ _5452_/B _5452_/C _5452_/A vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5379_ hold453/X _4434_/Y _5391_/S vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__mux2_1
Xfanout100 _3959_/X vssd1 vssd1 vccd1 vccd1 _6326_/C sky130_fd_sc_hd__buf_4
Xfanout111 _3669_/Y vssd1 vssd1 vccd1 vccd1 _6808_/B sky130_fd_sc_hd__clkbuf_8
Xfanout122 _7123_/A vssd1 vssd1 vccd1 vccd1 _6581_/A sky130_fd_sc_hd__buf_4
Xfanout155 _5788_/D vssd1 vssd1 vccd1 vccd1 _6518_/A sky130_fd_sc_hd__clkbuf_8
Xfanout144 _6851_/A vssd1 vssd1 vccd1 vccd1 _6718_/A sky130_fd_sc_hd__buf_8
Xfanout133 hold640/X vssd1 vssd1 vccd1 vccd1 _6872_/A sky130_fd_sc_hd__clkbuf_8
X_7118_ _7137_/A _6297_/X _7117_/Y vssd1 vssd1 vccd1 vccd1 _7118_/X sky130_fd_sc_hd__o21a_1
Xfanout188 _3930_/S1 vssd1 vssd1 vccd1 vccd1 _3913_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout177 _4244_/S1 vssd1 vssd1 vccd1 vccd1 _4255_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout199 _7341_/Q vssd1 vssd1 vccd1 vccd1 _4369_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout166 _7551_/Q vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__clkbuf_8
X_7049_ input35/X _4021_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _7049_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5420__A1 _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5184__A0 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5239__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6987__A1 _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5250__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4998__B1 _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3896__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4750_ _4789_/B _4750_/B vssd1 vssd1 vccd1 vccd1 _7212_/C sky130_fd_sc_hd__and2_2
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7164__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4681_ _4637_/X _4680_/X _4721_/S vssd1 vssd1 vccd1 vccd1 _7256_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3701_ _5988_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3988_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3632_ _6683_/A vssd1 vssd1 vccd1 vccd1 _6630_/A sky130_fd_sc_hd__inv_2
X_6420_ _6420_/A _6427_/A vssd1 vssd1 vccd1 vccd1 _6420_/Y sky130_fd_sc_hd__nand2_1
X_6351_ _6351_/A _6351_/B vssd1 vssd1 vccd1 vccd1 _6351_/Y sky130_fd_sc_hd__nand2_1
X_5302_ hold304/X _5022_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _7435_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6282_ _6282_/A _7110_/A _6282_/C _6949_/B vssd1 vssd1 vccd1 vccd1 _6282_/X sky130_fd_sc_hd__or4b_1
X_5233_ hold543/X _4864_/X _5247_/S vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__mux2_1
X_5164_ _5163_/X _4394_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7373_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4150__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4115_ _4846_/A _5990_/A _4115_/C vssd1 vssd1 vccd1 vccd1 _4118_/C sky130_fd_sc_hd__and3_1
XANTENNA_fanout189_A _7361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5095_ _7175_/B _7211_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5112_/S sky130_fd_sc_hd__and3_4
XANTENNA__4057__B _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ _4067_/A _4067_/B _4046_/C _4046_/D vssd1 vssd1 vccd1 vccd1 _7241_/S sky130_fd_sc_hd__or4_4
XANTENNA__4772__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5650__A1 _6273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _3644_/A _3645_/Y _3646_/A _3647_/Y _5996_/X vssd1 vssd1 vccd1 vccd1 _6004_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6272__B _6882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4948_ _4948_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _4948_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7155__A1 _4394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4879_ _4878_/X _4873_/A _4879_/S vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6618_ _6579_/Y _6618_/B vssd1 vssd1 vccd1 vccd1 _6619_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7598_ _7598_/CLK _7598_/D vssd1 vssd1 vccd1 vccd1 _7598_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6902__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6549_ _6557_/B _6557_/C _6557_/A vssd1 vssd1 vccd1 vccd1 _6558_/A sky130_fd_sc_hd__o21a_1
XANTENNA__4141__B2 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4248__A _5026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5641__B2 _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__A1 _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4683__A2 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6409__A0 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7082__B1 _4723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3869__S1 _3883_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5920_ _5941_/B _5920_/B vssd1 vssd1 vccd1 vccd1 _5922_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ _5838_/A _5838_/B _5841_/A vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__5396__A0 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4802_ _4589_/X hold393/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7289_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5782_ _6802_/A _6808_/A _6872_/B _6807_/A vssd1 vssd1 vccd1 vccd1 _5782_/X sky130_fd_sc_hd__and4_1
X_4733_ hold457/X _4434_/Y _4745_/S vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7521_ _7534_/CLK _7521_/D vssd1 vssd1 vccd1 vccd1 _7521_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5148__A0 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7452_ _7453_/CLK hold67/X vssd1 vssd1 vccd1 vccd1 _7452_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4664_ _7282_/Q _7597_/Q _7266_/Q _7490_/Q _4706_/S0 _4706_/S1 vssd1 vssd1 vccd1
+ vccd1 _4664_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5436__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6403_ hold142/X _6415_/A _6356_/B hold60/X vssd1 vssd1 vccd1 vccd1 _6403_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5699__A1 _6581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7383_ _7400_/CLK _7383_/D vssd1 vssd1 vccd1 vccd1 _7383_/Q sky130_fd_sc_hd__dfxtp_1
X_4595_ _4689_/A _4595_/B vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6334_ _6974_/B _6259_/B _6948_/B vssd1 vssd1 vccd1 vccd1 _6978_/C sky130_fd_sc_hd__a21o_1
XANTENNA_fanout104_A _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__S _4767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6265_ _6279_/B _6265_/B vssd1 vssd1 vccd1 vccd1 _6265_/Y sky130_fd_sc_hd__nand2b_1
X_5216_ hold398/X _4849_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _7396_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5452__A _5452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6196_ _6198_/A _6196_/B vssd1 vssd1 vccd1 vccd1 _7532_/D sky130_fd_sc_hd__nand2_1
X_5147_ hold502/X _4912_/Y _5157_/S vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _5322_/B _7194_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5093_/S sky130_fd_sc_hd__and3_4
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5623__A1 _6445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4029_ _6223_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _4029_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_79_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3700__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit27 _6718_/A vssd1 vssd1 vccd1 vccd1 _6716_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4285__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4114__A1 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7228__S _7228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold208 _7428_/Q vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold219 _7610_/Q vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_4380_ _6071_/B _6062_/B _6089_/B _4474_/A vssd1 vssd1 vccd1 vccd1 _4380_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6049_/X hold48/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__mux2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4200__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5001_ _5001_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5001_/X sky130_fd_sc_hd__or2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__B2 _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5853__A1 _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7055__B1 _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5211__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6952_ _7078_/A _6952_/B _6952_/C _6952_/D vssd1 vssd1 vccd1 vccd1 _6952_/X sky130_fd_sc_hd__or4_1
XANTENNA__4335__B _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6883_ _6852_/Y _6856_/X _6884_/B vssd1 vssd1 vccd1 vccd1 _6883_/X sky130_fd_sc_hd__a21o_1
X_5903_ _5904_/A _5904_/B _5904_/C vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _5834_/A _5834_/B _5834_/C vssd1 vssd1 vccd1 vccd1 _5834_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__6030__A1 _4862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5765_ _5797_/A _5797_/B _5797_/C vssd1 vssd1 vccd1 vccd1 _5798_/A sky130_fd_sc_hd__a21o_1
XANTENNA__4041__B1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6042__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4716_ _7607_/Q _4638_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4716_/Y sky130_fd_sc_hd__a21oi_1
X_7504_ _7581_/CLK hold51/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfxtp_1
X_5696_ _6628_/A _6637_/A _6338_/A vssd1 vssd1 vccd1 vccd1 _5697_/B sky130_fd_sc_hd__and3_1
X_7435_ _7443_/CLK _7435_/D vssd1 vssd1 vccd1 vccd1 _7435_/Q sky130_fd_sc_hd__dfxtp_1
X_4647_ _4645_/X _4646_/X _4692_/S vssd1 vssd1 vccd1 vccd1 _4647_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7366_ _7400_/CLK _7366_/D vssd1 vssd1 vccd1 vccd1 _7366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4578_ _5034_/B _4578_/B _4625_/B vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__or3_1
X_6317_ _6974_/B _6934_/B _6258_/A vssd1 vssd1 vccd1 vccd1 _6318_/B sky130_fd_sc_hd__a21o_1
X_7297_ _7618_/CLK _7297_/D vssd1 vssd1 vccd1 vccd1 _7297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6097__A1 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6278__A _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6248_ _6962_/A _6869_/A vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__nand2_2
X_6179_ _6179_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__or2_1
XANTENNA__7046__B1 _4029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5121__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4960__S _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7372_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6460__B _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4194__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__buf_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5031__S _5031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4497__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3880_ _6075_/A _4971_/B vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__and2_1
XFILLER_0_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4171__A _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__A1 _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5550_ _5493_/A _5554_/A split8/X vssd1 vssd1 vccd1 vccd1 _5550_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4501_ _7271_/Q _7611_/Q _7603_/Q _7619_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4501_/X sky130_fd_sc_hd__mux4_1
X_5481_ hold86/A _6683_/B vssd1 vssd1 vccd1 vccd1 _5481_/Y sky130_fd_sc_hd__nand2_1
X_4432_ _7351_/Q _7600_/Q _7601_/Q _5037_/B vssd1 vssd1 vccd1 vccd1 _4493_/C sky130_fd_sc_hd__or4_4
X_7220_ hold367/X _4492_/X _7228_/S vssd1 vssd1 vccd1 vccd1 _7619_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5206__S _5212_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7151_ _7212_/B _7151_/B _7194_/C vssd1 vssd1 vccd1 vccd1 _7166_/S sky130_fd_sc_hd__and3_4
X_4363_ _4362_/X _4361_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4363_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6098__A _6153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4294_ _4292_/X _4293_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__mux2_1
X_6102_ _4103_/A _6027_/Y _6427_/B vssd1 vssd1 vccd1 vccd1 _6102_/Y sky130_fd_sc_hd__a21oi_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7082_ _7059_/X _7081_/X _4723_/A vssd1 vssd1 vccd1 vccd1 _7082_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4185__S0 _4255_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6033_ _4873_/A _6035_/B _6142_/S vssd1 vssd1 vccd1 vccd1 _6034_/A sky130_fd_sc_hd__mux2_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5826__A1 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7028__B1 _6326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6826__A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer12 rebuffer16/X vssd1 vssd1 vccd1 vccd1 _6601_/A sky130_fd_sc_hd__clkbuf_1
Xrebuffer34 rebuffer4/X vssd1 vssd1 vccd1 vccd1 rebuffer5/A sky130_fd_sc_hd__clkbuf_1
Xrebuffer23 _5589_/C vssd1 vssd1 vccd1 vccd1 _5611_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4065__B _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ _6935_/A _7230_/A vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__or2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4780__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6866_ _6862_/B _6874_/C _6865_/X _6811_/B vssd1 vssd1 vccd1 vccd1 _6866_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6561__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4014__B1 _7244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6797_ _6803_/A1 _6774_/Y _6739_/B _6765_/X vssd1 vssd1 vccd1 vccd1 _6797_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5817_ _6581_/A _6628_/A _5854_/C _6702_/A vssd1 vssd1 vccd1 vccd1 _5818_/D sky130_fd_sc_hd__nand4_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5748_ _7009_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _5749_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5679_ _5714_/B _5679_/B vssd1 vssd1 vccd1 vccd1 _5681_/B sky130_fd_sc_hd__nand2_1
X_7418_ _7418_/CLK _7418_/D vssd1 vssd1 vccd1 vccd1 _7418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold572 _7461_/Q vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _5151_/X vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _7318_/Q vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5116__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7349_ _7424_/CLK _7349_/D vssd1 vssd1 vccd1 vccd1 _7349_/Q sky130_fd_sc_hd__dfxtp_1
Xhold594 _7445_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _7355_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4176__S0 _4686_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A _4147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6471__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4308__A1 _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5534__B _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 _7519_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XANTENNA_output65_A _7581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4865__S _5039_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3819__B1 _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3914__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4981_ _5024_/S _4228_/Y _4980_/Y _5008_/A vssd1 vssd1 vccd1 vccd1 _4982_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4795__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _3827_/S _3931_/X _3928_/X vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__a21oi_4
X_6720_ _6697_/B _6719_/X split7/A vssd1 vssd1 vccd1 vccd1 _6722_/B sky130_fd_sc_hd__mux2_2
XANTENNA__5992__B1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3863_ _7316_/Q _7332_/Q _7308_/Q _7444_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3863_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6651_ _6651_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _6651_/X sky130_fd_sc_hd__or2_1
X_5602_ _5605_/B _5601_/B _6518_/A vssd1 vssd1 vccd1 vccd1 _5609_/A sky130_fd_sc_hd__a21oi_1
X_6582_ _6583_/B _6583_/C _6581_/X _6576_/A vssd1 vssd1 vccd1 vccd1 _6586_/B sky130_fd_sc_hd__a211o_1
XANTENNA__4642__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3794_ _3792_/X _3793_/X _3886_/S vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5533_ _5818_/B _5534_/A vssd1 vssd1 vccd1 vccd1 _5533_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5725__A _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5464_ _5818_/B _5464_/B vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__nand2_1
X_5395_ hold574/X _4385_/X _5409_/S vssd1 vssd1 vccd1 vccd1 _5395_/X sky130_fd_sc_hd__mux2_1
X_7203_ hold173/X _4580_/X _7209_/S vssd1 vssd1 vccd1 vccd1 _7203_/X sky130_fd_sc_hd__mux2_1
X_4415_ _5031_/S _4411_/X _4413_/X _4414_/Y vssd1 vssd1 vccd1 vccd1 _4431_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4346_ _7420_/Q _7352_/Q _7344_/Q _7324_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4346_/X sky130_fd_sc_hd__mux4_1
X_7134_ _7137_/A _6276_/B _7091_/X _7558_/Q vssd1 vssd1 vccd1 vccd1 _7134_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4775__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4277_ _4930_/S _4276_/X _4275_/X _5031_/S vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__o211a_1
X_7065_ _6247_/B _7039_/Y _7074_/A vssd1 vssd1 vccd1 vccd1 _7065_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6556__A _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3905__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3899__B _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6016_ _3988_/C _5988_/X _6417_/B vssd1 vssd1 vccd1 vccd1 _7168_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6224__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4786__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6918_ _4084_/A _3775_/Y _6922_/C _3728_/A vssd1 vssd1 vccd1 vccd1 _6918_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5983__B1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6849_ _6862_/B _6874_/C _6847_/Y _6848_/X vssd1 vssd1 vccd1 vccd1 _6849_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5635__A _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6160__A0 _4694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 _7617_/Q vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold391 _5262_/X vssd1 vssd1 vccd1 vccd1 _7417_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7620_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4226__B1 _3668_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4777__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6405__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5726__B1 _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer3 _5589_/X vssd1 vssd1 vccd1 vccd1 _5620_/B sky130_fd_sc_hd__buf_1
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6151__A0 _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4200_ _7439_/Q _7431_/Q _7415_/Q _7407_/Q _4244_/S0 _4244_/S1 vssd1 vssd1 vccd1
+ vccd1 _4201_/B sky130_fd_sc_hd__mux4_1
X_5180_ _4849_/X hold532/X _5194_/S vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4131_ _4007_/B _3960_/C _4039_/C _4128_/C _4007_/A vssd1 vssd1 vccd1 vccd1 _4131_/X
+ sky130_fd_sc_hd__o2111a_1
X_4062_ _6142_/S _6220_/C vssd1 vssd1 vccd1 vccd1 _4062_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4312__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _4948_/Y _4963_/X _4964_/S vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__mux2_8
XANTENNA__4768__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3915_ _3915_/A _3915_/B vssd1 vssd1 vccd1 vccd1 _3915_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6703_ _6857_/A _6702_/B _6697_/B _6869_/A vssd1 vssd1 vccd1 vccd1 _6703_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4895_ _6935_/A _4945_/B _4893_/Y _4894_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4897_/B
+ sky130_fd_sc_hd__o221a_1
X_3846_ _7399_/Q _7391_/Q _7367_/Q _7383_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3846_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6634_ _6694_/A _6694_/B _6624_/Y vssd1 vssd1 vccd1 vccd1 _6699_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5193__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4615__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6565_ _6568_/B vssd1 vssd1 vccd1 vccd1 _6565_/Y sky130_fd_sc_hd__inv_2
X_3777_ _7557_/Q _3777_/B vssd1 vssd1 vccd1 vccd1 _3777_/X sky130_fd_sc_hd__or2_1
X_5516_ _5553_/B _5553_/C _5553_/A vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__a21o_4
XANTENNA__5455__A _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6050__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6496_ _6568_/A _6496_/B _6496_/C vssd1 vssd1 vccd1 vccd1 _6505_/B sky130_fd_sc_hd__and3_1
XANTENNA__6142__A0 _4601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5447_ _5818_/B _5455_/B _5460_/A _5445_/B _5442_/X vssd1 vssd1 vccd1 vccd1 _5452_/C
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout112 _3667_/Y vssd1 vssd1 vccd1 vccd1 _4401_/S sky130_fd_sc_hd__clkbuf_8
X_5378_ hold249/X _4111_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7476_/D sky130_fd_sc_hd__mux2_1
Xfanout101 _3705_/X vssd1 vssd1 vccd1 vccd1 _6989_/A sky130_fd_sc_hd__clkbuf_8
X_4329_ _4328_/X _4327_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__mux2_1
Xfanout156 _6807_/A vssd1 vssd1 vccd1 vccd1 _5788_/D sky130_fd_sc_hd__buf_6
Xfanout145 _7577_/Q vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__buf_8
Xfanout134 _7584_/Q vssd1 vssd1 vccd1 vccd1 _6808_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout123 hold643/X vssd1 vssd1 vccd1 vccd1 _7123_/A sky130_fd_sc_hd__clkbuf_8
X_7117_ _7137_/A _6297_/X _3716_/Y vssd1 vssd1 vccd1 vccd1 _7117_/Y sky130_fd_sc_hd__a21oi_1
Xfanout189 _7361_/Q vssd1 vssd1 vccd1 vccd1 _3930_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout178 _7453_/Q vssd1 vssd1 vccd1 vccd1 _4244_/S1 sky130_fd_sc_hd__buf_6
X_7048_ _7028_/X _7047_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _7048_/X sky130_fd_sc_hd__o21a_1
Xfanout167 _4037_/A vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__buf_6
XANTENNA__4456__B1 _4460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3849__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4759__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6133__A0 _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6196__A _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4542__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3700_ _5988_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__nor2_4
X_4680_ hold471/X _4679_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4680_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5175__A1 _4719_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ _6235_/A vssd1 vssd1 vccd1 vccd1 _6298_/A sky130_fd_sc_hd__inv_2
XANTENNA__7193__C _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6350_ _4039_/D _5980_/Y _6015_/C vssd1 vssd1 vccd1 vccd1 _6351_/B sky130_fd_sc_hd__o21ai_1
X_5301_ hold303/X _5038_/X _5301_/S vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6124__A0 _6123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6281_ _7019_/A _6974_/A _7074_/A _6988_/A vssd1 vssd1 vccd1 vccd1 _6282_/C sky130_fd_sc_hd__or4_1
X_5232_ _7212_/A _7151_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5247_/S sky130_fd_sc_hd__and3_4
XFILLER_0_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5163_ hold271/X _4434_/Y _5175_/S vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5883__C1 _6198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4114_ _6374_/A _6920_/A _6375_/A _3742_/C _3741_/B vssd1 vssd1 vccd1 vccd1 _4115_/C
+ sky130_fd_sc_hd__a32o_1
X_5094_ hold199/X _5022_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _7339_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4045_ _4846_/A _6328_/A _4042_/Y _4044_/Y _4068_/A vssd1 vssd1 vccd1 vccd1 _4046_/D
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5650__A2 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5996_ _5996_/A hold62/X vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__xor2_1
X_4947_ _4946_/A _4944_/Y _4945_/X _4946_/Y _5022_/A vssd1 vssd1 vccd1 vccd1 _4947_/X
+ sky130_fd_sc_hd__a311o_4
XFILLER_0_47_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4878_ _6807_/A _4123_/B _4877_/Y _4263_/B vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__o22a_1
X_3829_ _3886_/S _3829_/B vssd1 vssd1 vccd1 vccd1 _3829_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5166__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6617_ _6617_/A _6617_/B vssd1 vssd1 vccd1 vccd1 _6666_/A sky130_fd_sc_hd__nor2_1
X_7597_ _7597_/CLK _7597_/D vssd1 vssd1 vccd1 vccd1 _7597_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4913__A1 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6902__A2 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6548_ _6600_/A vssd1 vssd1 vccd1 vccd1 _6548_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6479_ _6521_/A _6509_/B vssd1 vssd1 vccd1 vccd1 _6481_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_30_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4141__A2 _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5124__S _5130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6418__A1 _6417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4429__B1 _4986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4963__S _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__A2 _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5157__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5542__B _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5632__A2 _6871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5850_ hold82/X wire79/X _5849_/X _6198_/A vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__o211a_1
X_4801_ hold392/X _4629_/X _4805_/S vssd1 vssd1 vccd1 vccd1 _4801_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5781_ _6872_/A _6807_/A vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4732_ hold265/X _4111_/X _4746_/S vssd1 vssd1 vccd1 vccd1 _7260_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7520_ _7534_/CLK _7520_/D vssd1 vssd1 vccd1 vccd1 _7520_/Q sky130_fd_sc_hd__dfxtp_2
X_7451_ _7451_/CLK _7451_/D vssd1 vssd1 vccd1 vccd1 _7451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ input6/X _4982_/A _4661_/X _4662_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4663_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5209__S _5211_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6402_ _6401_/X hold658/X _6414_/S vssd1 vssd1 vccd1 vccd1 _6402_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5699__A2 _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7382_ _7396_/CLK _7382_/D vssd1 vssd1 vccd1 vccd1 _7382_/Q sky130_fd_sc_hd__dfxtp_1
X_4594_ _4592_/X _4593_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4595_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6333_ _6333_/A _6333_/B _6333_/C vssd1 vssd1 vccd1 vccd1 _6333_/X sky130_fd_sc_hd__or3_1
X_6264_ _6264_/A _6264_/B vssd1 vssd1 vccd1 vccd1 _6265_/B sky130_fd_sc_hd__or2_1
XANTENNA__5320__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5215_ hold397/X _4864_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6195_ _3652_/Y _3653_/Y _6207_/S vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__mux2_1
X_5146_ _4871_/Y hold465/X _5158_/S vssd1 vssd1 vccd1 vccd1 _7365_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4783__S _4785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5077_ _5159_/C _7193_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5094_/S sky130_fd_sc_hd__and3_4
XFILLER_0_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ _4846_/A _4039_/A _7168_/A _4953_/A vssd1 vssd1 vccd1 vccd1 _4067_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4084__A _4084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit17 _6862_/B vssd1 vssd1 vccd1 vccd1 _6888_/A sky130_fd_sc_hd__buf_1
XFILLER_0_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5387__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5979_ _5979_/A _5979_/B vssd1 vssd1 vccd1 vccd1 _7169_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5119__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6739__A _6875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5643__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5311__A1 _4937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4259__A _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7064__A1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5378__A1 _4111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6413__S _6413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5818__A _6516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4050__A1 hold213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 _5287_/X vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A1 _5022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5000_ _4238_/A _4974_/Y _4999_/X vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__a21bo_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__A2 _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6951_ _6944_/X _6950_/X _7043_/S vssd1 vssd1 vccd1 vccd1 _6952_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6882_ _6882_/A _6882_/B vssd1 vssd1 vccd1 vccd1 _6884_/B sky130_fd_sc_hd__nor2_1
X_5902_ _5927_/B _5902_/B vssd1 vssd1 vccd1 vccd1 _5904_/C sky130_fd_sc_hd__or2_1
XANTENNA__5369__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5833_ _5834_/A _5834_/B _5834_/C vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4632__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7503_ _7541_/CLK hold55/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfxtp_1
X_5764_ _5764_/A _5764_/B vssd1 vssd1 vccd1 vccd1 _5797_/C sky130_fd_sc_hd__nand2_1
X_4715_ _6166_/A _4714_/Y _4986_/S vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5695_ _6273_/A _6637_/A _6338_/A vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7434_ _7434_/CLK _7434_/D vssd1 vssd1 vccd1 vccd1 _7434_/Q sky130_fd_sc_hd__dfxtp_1
X_4646_ _7274_/Q _7614_/Q _7606_/Q _7622_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4646_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4778__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7365_ _4004_/A _7365_/D vssd1 vssd1 vccd1 vccd1 _7365_/Q sky130_fd_sc_hd__dfxtp_1
X_4577_ _4577_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _4625_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7154__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6316_ _6939_/A _6316_/B vssd1 vssd1 vccd1 vccd1 _6934_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5195__C_N _7193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7296_ _7306_/CLK _7296_/D vssd1 vssd1 vccd1 vccd1 _7296_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6278__B _6808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6247_ _6295_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _7019_/A sky130_fd_sc_hd__nand2_1
X_6178_ hold64/X hold46/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ hold568/X _5038_/X _5129_/S vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7046__B2 _6139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5402__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3711__A _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4804__A0 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold161_A _7521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3857__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5638__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4261__B _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4688__S _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5804__C _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4194__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit4 split4/A vssd1 vssd1 vccd1 vccd1 split4/X sky130_fd_sc_hd__clkbuf_2
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold8/X vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__clkbuf_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4559__C1 _4930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4500_ _7375_/Q _7303_/Q _7295_/Q _7287_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4500_/X sky130_fd_sc_hd__mux4_1
X_5480_ _6568_/A _5486_/C vssd1 vssd1 vccd1 vccd1 _5480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4598__S _4692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ _4964_/S _4431_/B _4431_/C vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__and3_1
XANTENNA_1 _4515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7150_ _7211_/B _7150_/B _7193_/C vssd1 vssd1 vccd1 vccd1 _7167_/S sky130_fd_sc_hd__and3_4
X_4362_ _7426_/Q _7358_/Q _7350_/Q _7330_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4362_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4293_ _7401_/Q _7393_/Q _7369_/Q _7385_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4293_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4709__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6101_ _5810_/A _4271_/A _6100_/Y _4122_/C _6027_/Y vssd1 vssd1 vccd1 vccd1 _6101_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7081_ _4031_/B _7079_/X _7080_/X vssd1 vssd1 vccd1 vccd1 _7081_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4185__S1 _4255_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6032_ _6031_/X hold54/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__mux2_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5826__A2 _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer35 _5557_/Y vssd1 vssd1 vccd1 vccd1 _5561_/A3 sky130_fd_sc_hd__clkbuf_1
Xrebuffer13 _6822_/A vssd1 vssd1 vccd1 vccd1 _6803_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6934_ _6949_/A _6934_/B vssd1 vssd1 vccd1 vccd1 _6934_/Y sky130_fd_sc_hd__xnor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout164_A _7551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7200__A1 _4443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5458__A _5854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6865_ _6865_/A _6865_/B vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6796_ _6796_/A _6796_/B vssd1 vssd1 vccd1 vccd1 _6796_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5816_ _6581_/A _6273_/A _5854_/C _6702_/A vssd1 vssd1 vccd1 vccd1 _5816_/X sky130_fd_sc_hd__and4_1
X_5747_ _5747_/A _5764_/A _5747_/C vssd1 vssd1 vccd1 vccd1 _5747_/X sky130_fd_sc_hd__and3_1
XFILLER_0_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4970__C1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7417_ _7441_/CLK _7417_/D vssd1 vssd1 vccd1 vccd1 _7417_/Q sky130_fd_sc_hd__dfxtp_1
X_5678_ _5677_/A _5677_/B _5677_/C vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4629_ _4989_/A _4613_/X _4628_/Y _4591_/Y vssd1 vssd1 vccd1 vccd1 _4629_/X sky130_fd_sc_hd__o31a_4
XANTENNA__6289__A _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 _5235_/X vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _7381_/Q vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _7451_/Q vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
X_7348_ _7423_/CLK _7348_/D vssd1 vssd1 vccd1 vccd1 _7348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold584 _7407_/Q vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _5351_/X vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
X_7279_ _7597_/CLK _7279_/D vssd1 vssd1 vccd1 vccd1 _7279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold595 _5325_/X vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4176__S1 _4686_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_A _6086_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4005__A1 _7542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5202__A0 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput60 _7542_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
Xoutput71 _7520_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_12
XANTENNA__3819__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output58_A _4006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3914__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3989__C _4122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _5024_/S _4980_/B vssd1 vssd1 vccd1 vccd1 _4980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3931_ _3929_/X _3930_/X _3931_/S vssd1 vssd1 vccd1 vccd1 _3931_/X sky130_fd_sc_hd__mux2_1
X_3862_ _7396_/Q _7388_/Q _7364_/Q _7380_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3862_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4182__A _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6650_ _6605_/X _6645_/Y _6646_/Y vssd1 vssd1 vccd1 vccd1 _6658_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5601_ _5605_/B _5601_/B vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__and2_1
X_6581_ _6581_/A _6683_/B vssd1 vssd1 vccd1 vccd1 _6581_/X sky130_fd_sc_hd__and2_1
XFILLER_0_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3793_ _7274_/Q _7614_/Q _7606_/Q _7622_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3793_/X sky130_fd_sc_hd__mux4_1
X_5532_ _5509_/B _5531_/Y _5532_/S vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6941__B1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5725__B _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5217__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5463_ _5457_/S _5460_/Y _5461_/X vssd1 vssd1 vccd1 vccd1 _5465_/B sky130_fd_sc_hd__o21a_1
X_5394_ _7212_/A _7212_/B _7151_/B vssd1 vssd1 vccd1 vccd1 _5409_/S sky130_fd_sc_hd__and3_4
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7202_ hold237/X _4492_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7611_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4704__C1 _4963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4414_ input30/X _5031_/S _4162_/B vssd1 vssd1 vccd1 vccd1 _4414_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4345_ _7316_/Q _7332_/Q _7308_/Q _7444_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4345_/X sky130_fd_sc_hd__mux4_1
X_7133_ _6276_/B _7091_/X _7137_/A vssd1 vssd1 vccd1 vccd1 _7133_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__7249__A1 hold92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4276_ _5024_/S _4262_/X _4270_/X vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__a21bo_1
X_7064_ _6900_/A _7074_/A _7060_/X _7063_/Y _3949_/Y vssd1 vssd1 vccd1 vccd1 _7064_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3905__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6015_ _6015_/A _6015_/B _6015_/C _7232_/B vssd1 vssd1 vccd1 vccd1 _7170_/B sky130_fd_sc_hd__and4_1
XFILLER_0_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4791__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6572__A _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6917_ _6906_/X _6916_/Y _4723_/A vssd1 vssd1 vccd1 vccd1 _6917_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6848_ _6848_/A _6854_/A _6848_/C vssd1 vssd1 vccd1 vccd1 _6848_/X sky130_fd_sc_hd__or3_1
XFILLER_0_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6779_ _6820_/B vssd1 vssd1 vccd1 vccd1 _6779_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5127__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5635__B _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold370 _5220_/X vssd1 vssd1 vccd1 vccd1 _7398_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold381 _7401_/Q vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4966__S _5040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3870__S _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 _7289_/Q vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold660_A _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4226__A1 _4688_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6482__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5726__A1 _6874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5726__B2 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4730__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3832__S0 _3896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer4 _5545_/X vssd1 vssd1 vccd1 vccd1 rebuffer4/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4130_ _7554_/Q _6920_/A _4846_/A vssd1 vssd1 vccd1 vccd1 _4267_/B sky130_fd_sc_hd__and3_1
XANTENNA__4267__A_N _5974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4061_ _6220_/C _4061_/B vssd1 vssd1 vccd1 vccd1 _4061_/X sky130_fd_sc_hd__or2_1
XANTENNA__4905__A _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4312__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4963_ _4960_/X _4962_/X _4963_/S vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3914_ _7375_/Q _7303_/Q _7295_/Q _7287_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3915_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_58_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6702_ _6702_/A _6702_/B vssd1 vssd1 vccd1 vccd1 _6714_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4894_ _4916_/B _4942_/B _4891_/Y _4279_/C _4081_/A vssd1 vssd1 vccd1 vccd1 _4894_/X
+ sky130_fd_sc_hd__a32o_1
X_6633_ _6685_/A _6632_/B _6629_/X vssd1 vssd1 vccd1 vccd1 _6694_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3845_ _3886_/S _3845_/B vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6914__B1 _7020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6390__A1 hold610/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6564_ _6511_/X _6563_/X _7090_/B vssd1 vssd1 vccd1 vccd1 _6568_/B sky130_fd_sc_hd__mux2_1
X_3776_ _6911_/A _7020_/A _6922_/B vssd1 vssd1 vccd1 vccd1 _3777_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5515_ _5526_/A _5514_/B _5498_/A vssd1 vssd1 vccd1 vccd1 _5553_/C sky130_fd_sc_hd__o21bai_4
X_6495_ _6496_/B _6496_/C _6568_/A vssd1 vssd1 vccd1 vccd1 _6529_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5446_ _5460_/A _5445_/B _5442_/X vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4786__S _4786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7162__S _7166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5377_ hold248/X _4385_/X _5391_/S vssd1 vssd1 vccd1 vccd1 _5377_/X sky130_fd_sc_hd__mux2_1
Xfanout113 _3667_/Y vssd1 vssd1 vccd1 vccd1 _4692_/S sky130_fd_sc_hd__buf_4
XANTENNA__5471__A _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 _3685_/Y vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__buf_6
X_4328_ _7422_/Q _7354_/Q _7346_/Q _7326_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4328_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout146 _6702_/A vssd1 vssd1 vccd1 vccd1 _6568_/A sky130_fd_sc_hd__buf_4
Xfanout135 hold662/X vssd1 vssd1 vccd1 vccd1 _6311_/A sky130_fd_sc_hd__buf_6
X_7116_ _7123_/A _6926_/Y _7114_/Y _7115_/X _7245_/C1 vssd1 vssd1 vccd1 vccd1 _7589_/D
+ sky130_fd_sc_hd__o221a_1
Xfanout124 _6628_/A vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__buf_4
Xfanout179 _4686_/S1 vssd1 vssd1 vccd1 vccd1 _4691_/S1 sky130_fd_sc_hd__clkbuf_8
X_4259_ _4999_/B vssd1 vssd1 vccd1 vccd1 _4974_/B sky130_fd_sc_hd__inv_2
Xfanout157 _7573_/Q vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__clkbuf_8
X_7047_ _4030_/B _7045_/X _7046_/X vssd1 vssd1 vccd1 vccd1 _7047_/X sky130_fd_sc_hd__o21ba_1
Xfanout168 _4057_/A vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4179__A1_N _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4456__A1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5410__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3865__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4550__A _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4144__B1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4542__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5556__A _5556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3805__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4907__C1 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6151__S _6160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3630_ _6427_/B vssd1 vssd1 vccd1 vccd1 _6374_/A sky130_fd_sc_hd__inv_6
X_5300_ hold197/X _4996_/X _5302_/S vssd1 vssd1 vccd1 vccd1 _7434_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ _7009_/B vssd1 vssd1 vccd1 vccd1 _6988_/A sky130_fd_sc_hd__inv_2
XANTENNA__4230__S0 _7452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5231_ _5393_/A _5321_/B _7150_/B vssd1 vssd1 vccd1 vccd1 _5248_/S sky130_fd_sc_hd__or3b_4
X_5162_ hold192/X _4111_/X _5176_/S vssd1 vssd1 vccd1 vccd1 _7372_/D sky130_fd_sc_hd__mux2_1
X_5093_ hold198/X _5038_/X _5093_/S vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__mux2_1
X_4113_ _6096_/A _4113_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _4113_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3909__A1_N _3827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4044_ _4044_/A _5804_/D vssd1 vssd1 vccd1 vccd1 _4044_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5230__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6060__A0 _4955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5995_ _6015_/A _5995_/B _6925_/A _5995_/D vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__nand4_2
X_4946_ _4946_/A _4946_/B vssd1 vssd1 vccd1 vccd1 _4946_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4610__A1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7157__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _4873_/A _4953_/B _4900_/B _6096_/A vssd1 vssd1 vccd1 vccd1 _4877_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3828_ _7441_/Q _7433_/Q _7417_/Q _7409_/Q _3896_/S0 _3896_/S1 vssd1 vssd1 vccd1
+ vccd1 _3829_/B sky130_fd_sc_hd__mux4_1
X_7596_ _7596_/CLK _7596_/D vssd1 vssd1 vccd1 vccd1 _7596_/Q sky130_fd_sc_hd__dfxtp_1
X_6616_ _6673_/A _6612_/B _6639_/B _6857_/A vssd1 vssd1 vccd1 vccd1 _6616_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6902__A3 _7098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6547_ _6710_/A _6652_/A vssd1 vssd1 vccd1 vccd1 _6600_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3759_ _3759_/A _7501_/Q vssd1 vssd1 vccd1 vccd1 _6211_/B sky130_fd_sc_hd__nor2_1
X_6478_ _6441_/Y _6475_/X _6477_/X _6435_/Y vssd1 vssd1 vccd1 vccd1 _6521_/D sky130_fd_sc_hd__a31o_4
XFILLER_0_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5405__S _5409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _6871_/A _5428_/B _5428_/C _5422_/Y vssd1 vssd1 vccd1 vccd1 _5438_/B sky130_fd_sc_hd__a31oi_4
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3714__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7076__C1 _3705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__A _4689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4280__A _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6935__A _6935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5093__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5050__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4840__A1 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4800_ _4538_/X _4799_/X _4806_/S vssd1 vssd1 vccd1 vccd1 _7288_/D sky130_fd_sc_hd__mux2_1
X_5780_ _5777_/C _5780_/B vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ hold264/X _4385_/X _4745_/S vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5286__A _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7450_ _7450_/CLK _7450_/D vssd1 vssd1 vccd1 vccd1 _7450_/Q sky130_fd_sc_hd__dfxtp_1
X_4662_ _4113_/Y _4652_/Y _5031_/S vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6401_ input35/X _6400_/X _6413_/S vssd1 vssd1 vccd1 vccd1 _6401_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7381_ _4004_/A _7381_/D vssd1 vssd1 vccd1 vccd1 _7381_/Q sky130_fd_sc_hd__dfxtp_1
X_4593_ _7481_/Q _7469_/Q _7461_/Q _7255_/Q _4686_/S0 _4686_/S1 vssd1 vssd1 vccd1
+ vccd1 _4593_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6332_ _6332_/A _6332_/B _6332_/C vssd1 vssd1 vccd1 vccd1 _6344_/S sky130_fd_sc_hd__or3_1
XFILLER_0_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6263_ _6974_/B _6974_/C _6974_/A vssd1 vssd1 vccd1 vccd1 _6264_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5225__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5214_ _5376_/A _5376_/C _5322_/C vssd1 vssd1 vccd1 vccd1 _5229_/S sky130_fd_sc_hd__and3_4
XANTENNA__4203__S0 _4244_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4659__A1 _6844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6194_ _6204_/A _6194_/B vssd1 vssd1 vccd1 vccd1 _7531_/D sky130_fd_sc_hd__or2_1
XANTENNA_fanout194_A _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5145_ hold464/X _4887_/X _5157_/S vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5084__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5076_ hold177/X _5022_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _7331_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6805__C1 _5788_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4365__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4027_ _7168_/A vssd1 vssd1 vccd1 vccd1 _4027_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4831__A1 _4434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6033__A0 _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit18 _6670_/A vssd1 vssd1 vccd1 vccd1 split18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6580__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _5978_/A _7232_/A vssd1 vssd1 vccd1 vccd1 _6013_/B sky130_fd_sc_hd__nor2_1
X_4929_ _6864_/A _4905_/B _4928_/X _4976_/B vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4690__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3709__A _6328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7579_ _7579_/CLK _7579_/D vssd1 vssd1 vccd1 vccd1 _7579_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5643__B _6311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5847__B1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3858__C1 _7363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4114__A3 _6375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5075__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4822__A1 _4637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6490__A _6754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5818__B _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6327__A1 _4037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4889__A1 _4871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5045__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5066__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6950_ _6989_/A _6978_/C _6948_/Y _6949_/Y _5879_/A vssd1 vssd1 vccd1 vccd1 _6950_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4813__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5901_ _5901_/A _5901_/B vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6881_ _6880_/A _6880_/B _6968_/A _6968_/B _6879_/X vssd1 vssd1 vccd1 vccd1 _7030_/B
+ sky130_fd_sc_hd__o41ai_4
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5832_ _5869_/B _5832_/B vssd1 vssd1 vccd1 vccd1 _5834_/C sky130_fd_sc_hd__nand2_1
X_5763_ _5763_/A _5763_/B _5763_/C vssd1 vssd1 vccd1 vccd1 _5764_/B sky130_fd_sc_hd__or3_1
XFILLER_0_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4632__B _6148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4714_ _6162_/B _4714_/B vssd1 vssd1 vccd1 vccd1 _4714_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4041__A2 _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7502_ _7582_/CLK _7502_/D vssd1 vssd1 vccd1 vccd1 _7502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5694_ _6630_/A _6857_/A vssd1 vssd1 vccd1 vccd1 _6338_/A sky130_fd_sc_hd__nor2_2
X_7433_ _7441_/CLK _7433_/D vssd1 vssd1 vccd1 vccd1 _7433_/Q sky130_fd_sc_hd__dfxtp_1
X_4645_ _7378_/Q _7306_/Q _7298_/Q _7290_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4645_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7364_ _4004_/A _7364_/D vssd1 vssd1 vccd1 vccd1 _7364_/Q sky130_fd_sc_hd__dfxtp_1
X_4576_ _4577_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _4578_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout207_A _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6315_ _7230_/A _6333_/B _6310_/Y _6989_/A _6314_/X vssd1 vssd1 vccd1 vccd1 _6315_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_7295_ _7379_/CLK _7295_/D vssd1 vssd1 vccd1 vccd1 _7295_/Q sky130_fd_sc_hd__dfxtp_1
X_6246_ _6295_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _7040_/B sky130_fd_sc_hd__and2_2
XANTENNA__4794__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6177_ _3751_/Y _6175_/X _6176_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6177_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4620__A_N _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5128_ _5127_/X _4996_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _7358_/D sky130_fd_sc_hd__mux2_1
XANTENNA__7046__A2 _5804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5057__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5059_ _5393_/A _7211_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5076_/S sky130_fd_sc_hd__and3b_4
XFILLER_0_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5638__B _6802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5517__C1 _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5296__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7596_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5048__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__clkbuf_2
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5220__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4879__S _4879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _6111_/A _5034_/B _4428_/Y _4429_/X _4162_/B vssd1 vssd1 vccd1 vccd1 _4431_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA_2 _6076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4361_ _7322_/Q _7338_/Q _7314_/Q _7450_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4361_/X sky130_fd_sc_hd__mux4_1
X_6100_ _6100_/A _6100_/B vssd1 vssd1 vccd1 vccd1 _6100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4292_ _7441_/Q _7433_/Q _7417_/Q _7409_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4292_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5287__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4709__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7080_ _6075_/A _5804_/C _4029_/Y _6148_/A _6326_/C vssd1 vssd1 vccd1 vccd1 _7080_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4908__A _4908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6031_ _4974_/B _6022_/Y _6030_/Y _7472_/Q vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__o22a_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5039__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer36 _5525_/A vssd1 vssd1 vccd1 vccd1 _5577_/B sky130_fd_sc_hd__clkbuf_1
Xrebuffer14 _6803_/A1 vssd1 vssd1 vccd1 vccd1 _6801_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4798__A0 _4492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6933_ _6989_/A _6933_/B _6933_/C vssd1 vssd1 vccd1 vccd1 _6933_/X sky130_fd_sc_hd__and3_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6864_ _6864_/A _6864_/B _6864_/C vssd1 vssd1 vccd1 vccd1 _6880_/A sky130_fd_sc_hd__and3_1
XFILLER_0_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6539__B2 _6481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5815_ _6581_/A _5854_/C _6702_/A _6273_/A vssd1 vssd1 vccd1 vccd1 _5818_/C sky130_fd_sc_hd__a22o_1
XANTENNA__5211__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4645__S0 _4691_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6795_ _6864_/A _6795_/B vssd1 vssd1 vccd1 vccd1 _6813_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5746_ _5747_/A _5764_/A _5747_/C vssd1 vssd1 vccd1 vccd1 _5800_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5677_ _5677_/A _5677_/B _5677_/C vssd1 vssd1 vccd1 vccd1 _5714_/B sky130_fd_sc_hd__or3_1
XANTENNA__7165__S _7167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7416_ _7449_/CLK _7416_/D vssd1 vssd1 vccd1 vccd1 _7416_/Q sky130_fd_sc_hd__dfxtp_1
X_4628_ _6148_/A _5034_/B _4627_/Y _4144_/Y vssd1 vssd1 vccd1 vccd1 _4628_/Y sky130_fd_sc_hd__a211oi_1
Xhold530 _5313_/X vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold563 _5181_/X vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _5337_/X vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _7357_/Q vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
X_7347_ _7423_/CLK _7347_/D vssd1 vssd1 vccd1 vccd1 _7347_/Q sky130_fd_sc_hd__dfxtp_2
X_4559_ _5024_/S _4554_/Y _4558_/Y _4930_/S vssd1 vssd1 vccd1 vccd1 _4559_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold574 _7484_/Q vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
X_7278_ _7483_/CLK _7278_/D vssd1 vssd1 vccd1 vccd1 _7278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold585 _7370_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _7317_/Q vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5278__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6229_ _3733_/A input38/X _6229_/S vssd1 vssd1 vccd1 vccd1 _6230_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4272__B _4879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6950__A1 _6989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4961__B1 _5034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6950__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6163__C1 _3975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput61 hold70/A vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
Xoutput50 _6799_/A vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
XFILLER_0_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5269__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 _7521_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
XANTENNA__5323__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4728__A _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3632__A _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3930_ _7275_/Q _7615_/Q _7607_/Q _7623_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3930_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _3915_/A _3861_/B vssd1 vssd1 vccd1 vccd1 _3861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5729__C1 _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3792_ _7378_/Q _7306_/Q _7298_/Q _7290_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3792_/X sky130_fd_sc_hd__mux4_1
X_5600_ _5660_/B _6840_/A _5561_/X _3659_/Y vssd1 vssd1 vccd1 vccd1 _5605_/C sky130_fd_sc_hd__a31o_1
X_6580_ _6742_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _6618_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4952__B1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5531_ _5536_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5531_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7201_ hold236/X _4529_/X _7209_/S vssd1 vssd1 vccd1 vccd1 _7201_/X sky130_fd_sc_hd__mux2_1
X_5462_ _5457_/S _5460_/Y _5461_/X vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__6154__C1 _3975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5393_ _5393_/A _5393_/B _7150_/B vssd1 vssd1 vccd1 vccd1 _5410_/S sky130_fd_sc_hd__or3b_4
X_4413_ _4930_/S _4413_/B vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4344_ _4343_/X _4360_/B vssd1 vssd1 vccd1 vccd1 _4344_/Y sky130_fd_sc_hd__nand2b_1
X_7132_ _6900_/A _6282_/A _7130_/Y _7131_/X _3949_/Y vssd1 vssd1 vccd1 vccd1 _7132_/X
+ sky130_fd_sc_hd__o221a_1
X_7063_ split4/A _7062_/X _6900_/A vssd1 vssd1 vccd1 vccd1 _7063_/Y sky130_fd_sc_hd__o21ai_1
X_4275_ _6872_/B _4658_/A _4274_/Y _5008_/A vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__a211o_1
X_6014_ _3980_/A _4033_/B _5990_/A vssd1 vssd1 vccd1 vccd1 _7232_/B sky130_fd_sc_hd__o21a_1
XANTENNA__5968__C1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6916_ _6908_/X _6915_/Y _6326_/C vssd1 vssd1 vccd1 vccd1 _6916_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7185__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3994__A1 _5990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6847_ _6848_/A _6854_/A _6848_/C vssd1 vssd1 vccd1 vccd1 _6847_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4618__S0 _4709_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6778_ _6718_/B _6832_/A _6777_/X _6745_/Y vssd1 vssd1 vccd1 vccd1 _6820_/B sky130_fd_sc_hd__o22a_2
X_5729_ _5727_/A _5749_/A _6244_/A _6807_/A vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__o211a_1
XANTENNA__5408__S _5410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3717__A _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold117_A _7524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6145__C1 _3975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold371 _7262_/Q vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _5079_/X vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _5226_/X vssd1 vssd1 vccd1 vccd1 _7401_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _4801_/X vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5143__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold653_A _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4934__A0 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5726__A2 _6869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6923__A1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4730__B _7151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3832__S1 _3896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer5 rebuffer5/A vssd1 vssd1 vccd1 vccd1 _5547_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6136__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7498_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output70_A _7519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5053__S _5057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ hold92/X hold315/X _6023_/S vssd1 vssd1 vccd1 vccd1 _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6673__A _6673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5414__A1 _6683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4962_ _6066_/A _4986_/S _4984_/B _4961_/Y vssd1 vssd1 vccd1 vccd1 _4962_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7167__A1 _4685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3913_ _7479_/Q _7467_/Q _7459_/Q _7253_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3913_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4893_ _4942_/B _4896_/B vssd1 vssd1 vccd1 vccd1 _4893_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6701_ _6702_/B vssd1 vssd1 vccd1 vccd1 _6701_/Y sky130_fd_sc_hd__inv_2
X_3844_ _7439_/Q _7431_/Q _7415_/Q _7407_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3845_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4921__A _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6632_ _6629_/X _6632_/B vssd1 vssd1 vccd1 vccd1 _6676_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5228__S _5230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6563_ _6563_/A _6563_/B vssd1 vssd1 vccd1 vccd1 _6563_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3775_ _6922_/B vssd1 vssd1 vccd1 vccd1 _3775_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6127__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5514_ _5526_/A _5514_/B vssd1 vssd1 vccd1 vccd1 _5520_/C sky130_fd_sc_hd__or2_1
XFILLER_0_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6494_ _6496_/B _6496_/C vssd1 vssd1 vccd1 vccd1 _6494_/Y sky130_fd_sc_hd__nand2_1
X_5445_ _5445_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5460_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5350__A0 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5752__A _6690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5376_ _5376_/A _7212_/B _5376_/C vssd1 vssd1 vccd1 vccd1 _5391_/S sky130_fd_sc_hd__and3_4
XFILLER_0_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7115_ input37/X _4021_/A _6927_/X vssd1 vssd1 vccd1 vccd1 _7115_/X sky130_fd_sc_hd__a21o_1
Xfanout103 _3685_/Y vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__clkbuf_4
Xfanout114 _3665_/Y vssd1 vssd1 vccd1 vccd1 _3827_/S sky130_fd_sc_hd__buf_8
X_4327_ _7318_/Q _7334_/Q _7310_/Q _7446_/Q _4369_/S0 _4369_/S1 vssd1 vssd1 vccd1
+ vccd1 _4327_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6059__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _6793_/A vssd1 vssd1 vccd1 vccd1 _6702_/A sky130_fd_sc_hd__buf_6
Xfanout136 _7583_/Q vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__buf_2
Xfanout125 _7025_/A vssd1 vssd1 vccd1 vccd1 _6628_/A sky130_fd_sc_hd__buf_4
X_4258_ _3668_/Y _4256_/X _4257_/X vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__a21oi_4
X_7046_ _6066_/A _5804_/C _4029_/Y _6139_/A _6329_/A vssd1 vssd1 vccd1 vccd1 _7046_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout158 _6872_/B vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__clkbuf_8
Xfanout169 _5805_/A vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__clkbuf_8
X_4189_ _4873_/A vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__inv_2
XANTENNA__5405__A1 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4307__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4613__C1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7158__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4392__A1 _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold190 _5369_/X vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7149__A1 _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5048__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4460__B _4460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3805__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4887__S _4964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ hold375/X _5022_/X _5230_/S vssd1 vssd1 vccd1 vccd1 _7403_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5332__A0 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4230__S1 _7453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5161_ hold191/X _4385_/X _5175_/S vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5092_ hold185/X _4996_/X _5094_/S vssd1 vssd1 vccd1 vccd1 _7338_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _6096_/A _4113_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__and3_2
XFILLER_0_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4043_ _5979_/A _4065_/C vssd1 vssd1 vccd1 vccd1 _5804_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4916__A _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5994_ _5991_/X _5994_/B _5994_/C _5994_/D vssd1 vssd1 vccd1 vccd1 _5995_/D sky130_fd_sc_hd__and4b_1
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4945_ _6244_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4945_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4651__A _4999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4876_ _4953_/A _4876_/B _4123_/B vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__or3b_4
X_7595_ _7598_/CLK _7595_/D vssd1 vssd1 vccd1 vccd1 _7595_/Q sky130_fd_sc_hd__dfxtp_1
X_3827_ _3823_/X _3826_/X _3827_/S vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5466__B _5660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6615_ _6857_/A _6639_/B vssd1 vssd1 vccd1 vccd1 _6640_/A sky130_fd_sc_hd__and2_1
XFILLER_0_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6546_ _6489_/Y _6545_/Y _7090_/B vssd1 vssd1 vccd1 vccd1 _6652_/A sky130_fd_sc_hd__mux2_1
X_3758_ _3759_/A _6216_/C vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4797__S _4805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3689_ _3983_/A _4044_/A vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__nand2_1
X_6477_ _6485_/B _6485_/C _6485_/D _6480_/B _6485_/A vssd1 vssd1 vccd1 vccd1 _6477_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5428_ _6871_/A _5428_/B _5428_/C vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__and3_1
X_5359_ hold545/X _4385_/X _5373_/S vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4098__A _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3714__B hold97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7029_ _7029_/A split4/A vssd1 vssd1 vccd1 vccd1 _7029_/X sky130_fd_sc_hd__and2_1
XANTENNA__3730__A _6223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5376__B _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7000__B1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3799__S0 _3913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7067__B1 _6900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6935__B _7230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5331__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3640__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _7212_/B _7151_/B _7176_/B vssd1 vssd1 vccd1 vccd1 _4745_/S sky130_fd_sc_hd__and3_4
XFILLER_0_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ _4659_/X _4660_/X _4118_/B vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7380_ _7396_/CLK _7380_/D vssd1 vssd1 vccd1 vccd1 _7380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6400_ _6244_/A _6383_/Y _6399_/X _6383_/A vssd1 vssd1 vccd1 vccd1 _6400_/X sky130_fd_sc_hd__a22o_1
X_4592_ _7281_/Q _7596_/Q _7265_/Q _7489_/Q _4691_/S0 _4691_/S1 vssd1 vssd1 vccd1
+ vccd1 _4592_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6331_ _6331_/A _6331_/B _6919_/B _6331_/D vssd1 vssd1 vccd1 vccd1 _6332_/C sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6262_ _6949_/A _6945_/B vssd1 vssd1 vccd1 vccd1 _6974_/C sky130_fd_sc_hd__or2_2
X_5213_ _5357_/A _5375_/C _5303_/C vssd1 vssd1 vccd1 vccd1 _5230_/S sky130_fd_sc_hd__and3b_4
XANTENNA__4203__S1 _4244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6193_ _5998_/A hold74/X _6207_/S vssd1 vssd1 vccd1 vccd1 _6193_/X sky130_fd_sc_hd__mux2_1
X_5144_ _4849_/X hold481/X _5158_/S vssd1 vssd1 vccd1 vccd1 _7364_/D sky130_fd_sc_hd__mux2_1
X_5075_ hold176/X _5038_/X _5075_/S vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout187_A _7361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4026_ _6374_/A _6223_/A _4030_/B vssd1 vssd1 vccd1 vccd1 _7168_/A sky130_fd_sc_hd__and3_1
XFILLER_0_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5977_ _6417_/B _5977_/B _6920_/A _5977_/D vssd1 vssd1 vccd1 vccd1 _7232_/A sky130_fd_sc_hd__or4_1
X_4928_ _5001_/A _4924_/X _4927_/X vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4690__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4859_ _4854_/X _4858_/X _4982_/A vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7578_ _7587_/CLK _7578_/D vssd1 vssd1 vccd1 vccd1 _7578_/Q sky130_fd_sc_hd__dfxtp_1
X_6529_ _6505_/D _6529_/B vssd1 vssd1 vccd1 vccd1 _6529_/X sky130_fd_sc_hd__and2b_1
XANTENNA__5643__C _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5151__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6024__A1 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4586__A1 _6628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5326__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3635__A _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6011__A _6204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6946__A _7070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5061__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4422__A_N _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5900_ _5901_/A _5901_/B vssd1 vssd1 vccd1 vccd1 _5927_/B sky130_fd_sc_hd__and2_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6681__A _6742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6880_ _6880_/A _6880_/B vssd1 vssd1 vccd1 vccd1 _6998_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _5831_/A _5831_/B vssd1 vssd1 vccd1 vccd1 _5832_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _5766_/A _5766_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5797_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4713_ _4674_/B _4674_/A _4713_/S vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7501_ _7581_/CLK _7501_/D vssd1 vssd1 vccd1 vccd1 _7501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5693_ _5840_/A _5693_/B vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__nand2_1
X_7432_ _7449_/CLK _7432_/D vssd1 vssd1 vccd1 vccd1 _7432_/Q sky130_fd_sc_hd__dfxtp_1
X_4644_ _4689_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4575_ _4479_/A _4478_/B _4526_/A _4574_/X vssd1 vssd1 vccd1 vccd1 _4577_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7363_ _7590_/CLK _7363_/D vssd1 vssd1 vccd1 vccd1 _7363_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5236__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7294_ _7618_/CLK _7294_/D vssd1 vssd1 vccd1 vccd1 _7294_/Q sky130_fd_sc_hd__dfxtp_1
X_6314_ _6314_/A _6333_/C _6313_/X vssd1 vssd1 vccd1 vccd1 _6314_/X sky130_fd_sc_hd__or3b_1
X_6245_ _6630_/A _6793_/A vssd1 vssd1 vccd1 vccd1 _6247_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6856__A _6857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6176_ _6176_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6176_/X sky130_fd_sc_hd__or2_1
X_5127_ hold365/X _5015_/X _5129_/S vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4376__A _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5058_ hold300/X _5022_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _7323_/D sky130_fd_sc_hd__mux2_1
X_4009_ _4009_/A _4039_/A vssd1 vssd1 vccd1 vccd1 _6331_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5638__C _6637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5517__B1 _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4740__A1 _4538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5146__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5670__A _6808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3926__S0 _3930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__buf_1
XFILLER_0_98_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4225__S _4401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5508__B1 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_3 _6085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4731__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _4359_/X _4360_/B vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5056__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4291_ _6098_/B _4672_/B vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__xor2_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5580__A _6445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6030_ _4862_/A _6027_/Y _6029_/X vssd1 vssd1 vccd1 vccd1 _6030_/Y sky130_fd_sc_hd__a21oi_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__B _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4342__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6932_ _6949_/A _6948_/B _6932_/C vssd1 vssd1 vccd1 vccd1 _6933_/C sky130_fd_sc_hd__nand3b_1
X_6863_ _6864_/B _6864_/C vssd1 vssd1 vccd1 vccd1 _6869_/B sky130_fd_sc_hd__nand2_1
X_5814_ _5715_/B _5814_/B vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4645__S1 _4691_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6794_ _6702_/A _6793_/B _6795_/B _6864_/A vssd1 vssd1 vccd1 vccd1 _6794_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4318__A_N _4360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5745_ _5745_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5747_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__4970__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5676_ _5714_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _5677_/C sky130_fd_sc_hd__nand2_1
X_7415_ _7439_/CLK _7415_/D vssd1 vssd1 vccd1 vccd1 _7415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4627_ _4625_/X _4626_/Y _5034_/B vssd1 vssd1 vccd1 vccd1 _4627_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold520 _7385_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold531 _7380_/Q vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _7313_/Q vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _5126_/X vssd1 vssd1 vccd1 vccd1 _7357_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7346_ _7454_/CLK _7346_/D vssd1 vssd1 vccd1 vccd1 _7346_/Q sky130_fd_sc_hd__dfxtp_1
X_4558_ _5024_/S _4601_/B vssd1 vssd1 vccd1 vccd1 _4558_/Y sky130_fd_sc_hd__nor2_1
Xhold575 _5395_/X vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
X_7277_ _7485_/CLK _7277_/D vssd1 vssd1 vccd1 vccd1 _7277_/Q sky130_fd_sc_hd__dfxtp_1
Xhold586 _5155_/X vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _5045_/X vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _7329_/Q vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _6962_/A _4440_/A _4440_/Y _4488_/X vssd1 vssd1 vccd1 vccd1 _4489_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6586__A _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6228_ _7244_/A _6228_/B vssd1 vssd1 vccd1 vccd1 _7554_/D sky130_fd_sc_hd__or2_1
XANTENNA__6475__A1 _6532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6158_/X hold62/X _6168_/S vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__mux2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6227__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4333__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5665__A _6683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5910__B1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput51 _6637_/A vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
XANTENNA__6496__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput62 _7259_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
Xoutput73 _7522_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__4728__B _4728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4324__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3860_ _7436_/Q _7428_/Q _7412_/Q _7404_/Q _3883_/S0 _3883_/S1 vssd1 vssd1 vccd1
+ vccd1 _3861_/B sky130_fd_sc_hd__mux4_1
XANTENNA__5729__B1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3791_ _3886_/S _3791_/B vssd1 vssd1 vccd1 vccd1 _3791_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3794__S _3886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4952__A1 _6793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5530_ _5530_/A _5530_/B vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5575__A _6568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5461_ _5454_/A _5454_/B _5454_/C _5441_/B vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7200_ hold220/X _4443_/X _7210_/S vssd1 vssd1 vccd1 vccd1 _7610_/D sky130_fd_sc_hd__mux2_1
X_4412_ _4407_/B _4406_/X _5024_/S vssd1 vssd1 vccd1 vccd1 _4413_/B sky130_fd_sc_hd__mux2_1
X_5392_ _5391_/X _4685_/X _5392_/S vssd1 vssd1 vccd1 vccd1 _7483_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4704__A1 _3677_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4343_ _4341_/X _4342_/X _4421_/S vssd1 vssd1 vccd1 vccd1 _4343_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7131_ _6840_/B split4/A _7043_/S vssd1 vssd1 vccd1 vccd1 _7131_/X sky130_fd_sc_hd__a21o_1
X_4274_ _4272_/Y _4273_/X _4658_/A vssd1 vssd1 vccd1 vccd1 _4274_/Y sky130_fd_sc_hd__a21oi_1
X_7062_ _7062_/A _7062_/B vssd1 vssd1 vccd1 vccd1 _7062_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_94_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6013_ _7233_/A _6013_/B _4033_/X vssd1 vssd1 vccd1 vccd1 _7171_/A sky130_fd_sc_hd__or3b_1
XANTENNA__4563__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6209__A1 _6922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4315__S0 _4371_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6090__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6915_ _6913_/A _6914_/Y _6910_/X vssd1 vssd1 vccd1 vccd1 _6915_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4640__B1 _4529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4140__A_N _6326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6984__B1_N _6983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6846_ _6887_/A vssd1 vssd1 vccd1 vccd1 _7085_/A sky130_fd_sc_hd__inv_2
XFILLER_0_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4618__S1 _4709_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6777_ _6766_/A _6721_/Y _6782_/A _6775_/Y vssd1 vssd1 vccd1 vccd1 _6777_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6393__A0 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5728_ _7009_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _5749_/A sky130_fd_sc_hd__nor2_1
X_3989_ _6922_/D _4015_/B _4122_/C vssd1 vssd1 vccd1 vccd1 _3989_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3717__B _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5659_ _5659_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5660_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold361 _7392_/Q vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 _7613_/Q vssd1 vssd1 vccd1 vccd1 hold350/X sky130_fd_sc_hd__dlygate4sd3_1
X_7329_ _7424_/CLK _7329_/D vssd1 vssd1 vccd1 vccd1 _7329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold372 _4735_/X vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _7402_/Q vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _7421_/Q vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4459__A0 _6799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5120__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__S0 _4369_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6081__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4631__A0 _4589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5187__A1 _4964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer6 _5547_/A1 vssd1 vssd1 vccd1 vccd1 _5573_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5334__S _5338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7443_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output63_A _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5111__A1 _5038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4474__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4870__B1 _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6072__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5414__A2 _6518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4961_ _4355_/A _4355_/B _5034_/B vssd1 vssd1 vccd1 vccd1 _4961_/Y sky130_fd_sc_hd__a21oi_1
X_3912_ _3931_/S _3912_/B vssd1 vssd1 vccd1 vccd1 _3912_/X sky130_fd_sc_hd__and2_1
X_4892_ _4915_/B _4892_/B vssd1 vssd1 vccd1 vccd1 _4896_/B sky130_fd_sc_hd__nor2_1
X_6700_ _6637_/B _6699_/X _6709_/S vssd1 vssd1 vccd1 vccd1 _6702_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_104_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3843_ _3827_/S _3841_/X _3842_/Y _3838_/Y vssd1 vssd1 vccd1 vccd1 _6066_/A sky130_fd_sc_hd__o2bb2a_2
X_6631_ _6629_/B _6629_/C _6629_/A vssd1 vssd1 vccd1 vccd1 _6632_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4925__A1 _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6562_ _6871_/A _6524_/B _6570_/A vssd1 vssd1 vccd1 vccd1 _6563_/B sky130_fd_sc_hd__a21bo_1
X_3774_ _6911_/B _3962_/C vssd1 vssd1 vccd1 vccd1 _6922_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5513_ _5530_/A _5512_/B _5504_/A _5504_/B vssd1 vssd1 vccd1 vccd1 _5514_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6493_ _6454_/B _6521_/D _6521_/A vssd1 vssd1 vccd1 vccd1 _6496_/C sky130_fd_sc_hd__nand3b_2
X_5444_ _5788_/D _5444_/B _5444_/C vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__and3_1
XFILLER_0_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5752__B _6807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5244__S _5248_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5375_ _5357_/A _7211_/B _5375_/C vssd1 vssd1 vccd1 vccd1 _5392_/S sky130_fd_sc_hd__and3b_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4649__A _4698_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7025__A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7114_ _7107_/X _7113_/X _4723_/A vssd1 vssd1 vccd1 vccd1 _7114_/Y sky130_fd_sc_hd__a21oi_1
Xfanout104 _6413_/S vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__clkbuf_8
Xfanout115 _3664_/Y vssd1 vssd1 vccd1 vccd1 _3886_/S sky130_fd_sc_hd__buf_6
X_4326_ _4325_/X _4360_/B vssd1 vssd1 vccd1 vccd1 _4326_/Y sky130_fd_sc_hd__nand2b_1
Xfanout137 _6710_/A vssd1 vssd1 vccd1 vccd1 _6773_/A sky130_fd_sc_hd__buf_4
Xfanout126 hold635/X vssd1 vssd1 vccd1 vccd1 _7025_/A sky130_fd_sc_hd__buf_4
X_4257_ _4688_/S _4251_/X _4253_/X _4689_/A vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5102__A1 _4897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6864__A _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout148 _7576_/Q vssd1 vssd1 vccd1 vccd1 _6793_/A sky130_fd_sc_hd__buf_8
X_7045_ _6244_/A _6793_/A _4037_/X _7032_/X _7044_/X vssd1 vssd1 vccd1 vccd1 _7045_/X
+ sky130_fd_sc_hd__o32a_1
Xfanout159 _6872_/B vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__clkbuf_4
X_4188_ _4689_/A _4186_/X _4187_/Y _4182_/Y vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__a2bb2o_2
XANTENNA__6063__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5169__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6366__A0 _7527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6829_ _6780_/X _6821_/X _6828_/Y vssd1 vssd1 vccd1 vccd1 _6862_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5341__A1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5154__S _5158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 _7519_/Q vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold191 _7372_/Q vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3910__B _6120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6054__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4080__A1 hold92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5329__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4907__A1 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5064__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5160_ _7212_/B _5376_/C _5322_/B vssd1 vssd1 vccd1 vccd1 _5175_/S sky130_fd_sc_hd__and3_4
X_5091_ hold184/X _5015_/X _5093_/S vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__mux2_1
X_4111_ _5022_/A _4111_/B vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__or2_4
X_4042_ _5977_/B _6220_/B vssd1 vssd1 vccd1 vccd1 _4042_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6045__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5399__A1 _4483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _6922_/D _5987_/X _5992_/X _4013_/Y vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__o211a_1
X_4944_ _4942_/B _4946_/B _4943_/X _4945_/B vssd1 vssd1 vccd1 vccd1 _4944_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4071__A1 hold66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4875_ _4900_/B _4875_/B vssd1 vssd1 vccd1 vccd1 _4875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6348__B1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7594_ _7597_/CLK _7594_/D vssd1 vssd1 vccd1 vccd1 _7594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3826_ _3824_/X _3825_/X _3931_/S vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__mux2_1
X_6614_ _6573_/B _6613_/Y split9/A vssd1 vssd1 vccd1 vccd1 _6639_/B sky130_fd_sc_hd__mux2_2
X_6545_ _6545_/A _6545_/B vssd1 vssd1 vccd1 vccd1 _6545_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3757_ _3757_/A _6207_/S _4267_/D vssd1 vssd1 vccd1 vccd1 _3762_/C sky130_fd_sc_hd__or3_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3688_ _6225_/A _4007_/A vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__nor2_2
X_6476_ _6532_/A _6476_/B vssd1 vssd1 vccd1 vccd1 _6480_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5323__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5427_ _5437_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5428_/C sky130_fd_sc_hd__or2_4
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _5376_/A _7212_/B _7194_/C vssd1 vssd1 vccd1 vccd1 _5373_/S sky130_fd_sc_hd__and3_4
X_4309_ _4474_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__and2_1
XANTENNA__7076__A1 _7043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5289_ hold294/X _4887_/X _5301_/S vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__mux2_1
X_7028_ _7020_/X _7023_/X _7044_/B _7027_/X _6326_/C vssd1 vssd1 vccd1 vccd1 _7028_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6036__C1 _6922_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6587__B1 _6629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5938__A _6235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4929__A1_N _6864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5149__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3799__S1 _3913_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5314__A1 _4947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4752__A _7212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4053__A1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5286__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _5024_/S _4652_/Y _4654_/Y _4930_/S vssd1 vssd1 vccd1 vccd1 _4660_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4591_ hold620/X _4638_/C _4590_/Y vssd1 vssd1 vccd1 vccd1 _4591_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6330_ _4036_/A _6922_/C _4044_/Y _6374_/A vssd1 vssd1 vccd1 vccd1 _6332_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5305__A1 _4864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4199__A _4873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6261_ _6261_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _6939_/A sky130_fd_sc_hd__nand2_2
XANTENNA__6502__B1 _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5212_ _5022_/X hold324/X _5212_/S vssd1 vssd1 vccd1 vccd1 _7395_/D sky130_fd_sc_hd__mux2_1
X_6192_ _3751_/Y _6190_/X _6191_/X _6198_/A vssd1 vssd1 vccd1 vccd1 _6192_/X sky130_fd_sc_hd__o211a_1
X_5143_ hold480/X _4864_/X _5157_/S vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7058__A1 _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5074_ _5073_/X _4996_/X _5076_/S vssd1 vssd1 vccd1 vccd1 _7330_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4025_ _5988_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _5804_/C sky130_fd_sc_hd__nor2_4
XFILLER_0_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5976_ _5976_/A vssd1 vssd1 vccd1 vccd1 _7169_/A sky130_fd_sc_hd__inv_2
X_4927_ _4955_/A _4698_/A _4925_/X _4926_/X _4263_/B vssd1 vssd1 vccd1 vccd1 _4927_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5196__C _5322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4858_ _6872_/B _4976_/B _4857_/X _5008_/A vssd1 vssd1 vccd1 vccd1 _4858_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3809_ _7272_/Q _7612_/Q _7604_/Q _7620_/Q _3930_/S0 _3930_/S1 vssd1 vssd1 vccd1
+ vccd1 _3809_/X sky130_fd_sc_hd__mux4_1
X_4789_ _4964_/S _4789_/B _4789_/C vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__and3_2
X_7577_ _7577_/CLK _7577_/D vssd1 vssd1 vccd1 vccd1 _7577_/Q sky130_fd_sc_hd__dfxtp_2
X_6528_ _6871_/A _6514_/B _6524_/B _6512_/Y vssd1 vssd1 vccd1 vccd1 _6557_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6459_ _6461_/A _6461_/B vssd1 vssd1 vccd1 vccd1 _6522_/A sky130_fd_sc_hd__or2_1
XANTENNA__3858__A1 _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7049__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4048__S _6329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7221__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4374__A_N _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4291__B _4672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__A2 _4440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5342__S _5356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7123__A _7123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6962__A _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _5831_/A _5831_/B vssd1 vssd1 vccd1 vccd1 _5869_/B sky130_fd_sc_hd__nand2_1
X_5761_ _5797_/A _5761_/B vssd1 vssd1 vccd1 vccd1 _5766_/C sky130_fd_sc_hd__and2_1
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4712_ _7343_/Q _4707_/X _4711_/X vssd1 vssd1 vccd1 vccd1 _6162_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7500_ _7581_/CLK _7500_/D vssd1 vssd1 vccd1 vccd1 _7500_/Q sky130_fd_sc_hd__dfxtp_1
X_7431_ _7441_/CLK _7431_/D vssd1 vssd1 vccd1 vccd1 _7431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5692_ _6516_/A _5788_/D _5665_/X _5677_/A vssd1 vssd1 vccd1 vccd1 _5693_/B sky130_fd_sc_hd__a211o_1
XANTENNA_hold70_A hold70/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4643_ _4641_/X _4642_/X _4688_/S vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4421__S _4421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4574_ _4672_/B _6126_/B _4478_/A _4525_/A vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__o211a_1
X_7362_ _7570_/CLK _7362_/D vssd1 vssd1 vccd1 vccd1 _7362_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__6202__A _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7293_ _7372_/CLK _7293_/D vssd1 vssd1 vccd1 vccd1 _7293_/Q sky130_fd_sc_hd__dfxtp_1
X_6313_ _7551_/Q _5805_/A _6421_/B _4037_/A vssd1 vssd1 vccd1 vccd1 _6313_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6244_ _6244_/A _6857_/A vssd1 vssd1 vccd1 vccd1 _7066_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6175_ hold84/X hold48/X _6190_/S vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__mux2_1
X_5126_ _5125_/X _4973_/X _5130_/S vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__mux2_1
X_5057_ hold299/X _5038_/X _5057_/S vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6872__A _6872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4008_ _6417_/B _6329_/A _4030_/B vssd1 vssd1 vccd1 vccd1 _4033_/B sky130_fd_sc_hd__or3_2
XANTENNA__7203__A1 _4580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5488__A _5556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4017__B2 _6374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5638__D _6702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5959_ _5958_/Y _5958_/B _6236_/A vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4973__C1 _5022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5517__A1 _5556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3736__A _6015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3926__S1 _3930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5162__S _5176_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xsplit7 split7/A vssd1 vssd1 vccd1 vccd1 split7/X sky130_fd_sc_hd__clkbuf_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__buf_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5989__D1 _4021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7379_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3862__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5337__S _5337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6022__A _6427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _7542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4290_ _6911_/B _4290_/B _6220_/C _4290_/D vssd1 vssd1 vccd1 vccd1 _4290_/X sky130_fd_sc_hd__or4_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5072__S _5076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6168__S _6168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer16 _6651_/A vssd1 vssd1 vccd1 vccd1 rebuffer16/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4342__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6931_ _6290_/X _6931_/B _7020_/A vssd1 vssd1 vccd1 vccd1 _6931_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6862_ _6799_/B _6862_/B _6874_/C vssd1 vssd1 vccd1 vccd1 _6864_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5813_ hold76/X wire79/X _5812_/X _6198_/A vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__o211a_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6793_ _6793_/A _6793_/B vssd1 vssd1 vccd1 vccd1 _6815_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3853__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ _5763_/A _5763_/B _5763_/C vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5675_ _5675_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__or2_1
X_7414_ _7430_/CLK _7414_/D vssd1 vssd1 vccd1 vccd1 _7414_/Q sky130_fd_sc_hd__dfxtp_1
X_4626_ _4625_/A _4625_/B _4625_/C vssd1 vssd1 vccd1 vccd1 _4626_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4151__S _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 _7459_/Q vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
X_7345_ _7423_/CLK _7345_/D vssd1 vssd1 vccd1 vccd1 _7345_/Q sky130_fd_sc_hd__dfxtp_1
Xhold521 _5190_/X vssd1 vssd1 vccd1 vccd1 _7385_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _7404_/Q vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _5179_/X vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _4992_/X vssd1 vssd1 vccd1 vccd1 _7313_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _5008_/A _4557_/B vssd1 vssd1 vccd1 vccd1 _4557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7276_ _7592_/CLK _7276_/D vssd1 vssd1 vccd1 vccd1 _7276_/Q sky130_fd_sc_hd__dfxtp_1
Xhold587 _5156_/X vssd1 vssd1 vccd1 vccd1 _7370_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _7311_/Q vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _5072_/X vssd1 vssd1 vccd1 vccd1 _7329_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _4488_/A _4533_/B vssd1 vssd1 vccd1 vccd1 _4488_/X sky130_fd_sc_hd__and2_1
Xhold598 _7367_/Q vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6078__S _6142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6227_ _3733_/B input37/X _6229_/S vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__mux2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6427_/B _6156_/X _6157_/Y _4649_/Y _7236_/B1 vssd1 vssd1 vccd1 vccd1 _6158_/X
+ sky130_fd_sc_hd__o32a_1
X_5109_ hold623/X _5015_/X _5111_/S vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__mux2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6153_/A _6089_/B vssd1 vssd1 vccd1 vccd1 _6089_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4333__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6107__A _6162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3844__S0 _3883_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5157__S _5157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5665__B _6962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput52 _6793_/A vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
Xoutput63 _7557_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
Xoutput74 _7523_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
XANTENNA__4324__S1 _4371_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _7482_/Q _7470_/Q _7462_/Q _7256_/Q _3913_/S0 _3913_/S1 vssd1 vssd1 vccd1
+ vccd1 _3791_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_66_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5067__S _5075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5460_ _5460_/A _5460_/B vssd1 vssd1 vccd1 vccd1 _5460_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4411_ _6875_/A _4658_/A _4410_/X _5008_/A vssd1 vssd1 vccd1 vccd1 _4411_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5391_ hold376/X _4719_/Y _5391_/S vssd1 vssd1 vccd1 vccd1 _5391_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4704__A2 _4982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__A _6710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ _7396_/Q _7388_/Q _7364_/Q _7380_/Q _4371_/S0 _4371_/S1 vssd1 vssd1 vccd1
+ vccd1 _4342_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7130_ split4/A _7130_/B vssd1 vssd1 vccd1 vccd1 _7130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4273_ _4262_/X _4266_/Y _4270_/X _4263_/B vssd1 vssd1 vccd1 vccd1 _4273_/X sky130_fd_sc_hd__o2bb2a_1
X_7061_ _7030_/A _7030_/B _6856_/X vssd1 vssd1 vccd1 vccd1 _7062_/B sky130_fd_sc_hd__a21oi_1
X_6012_ _4033_/B _4125_/X _5974_/X vssd1 vssd1 vccd1 vccd1 _7233_/A sky130_fd_sc_hd__o21ai_1
.ends

