magic
tech sky130B
magscale 1 2
timestamp 1717095420
<< obsli1 >>
rect 1104 2159 128892 122417
<< obsm1 >>
rect 658 1368 129246 122448
<< metal2 >>
rect 13082 124200 13138 125000
rect 39026 124200 39082 125000
rect 64970 124200 65026 125000
rect 90914 124200 90970 125000
rect 116858 124200 116914 125000
rect 662 0 718 800
rect 1674 0 1730 800
rect 2686 0 2742 800
rect 3698 0 3754 800
rect 4710 0 4766 800
rect 5722 0 5778 800
rect 6734 0 6790 800
rect 7746 0 7802 800
rect 8758 0 8814 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11794 0 11850 800
rect 12806 0 12862 800
rect 13818 0 13874 800
rect 14830 0 14886 800
rect 15842 0 15898 800
rect 16854 0 16910 800
rect 17866 0 17922 800
rect 18878 0 18934 800
rect 19890 0 19946 800
rect 20902 0 20958 800
rect 21914 0 21970 800
rect 22926 0 22982 800
rect 23938 0 23994 800
rect 24950 0 25006 800
rect 25962 0 26018 800
rect 26974 0 27030 800
rect 27986 0 28042 800
rect 28998 0 29054 800
rect 30010 0 30066 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 33046 0 33102 800
rect 34058 0 34114 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39118 0 39174 800
rect 40130 0 40186 800
rect 41142 0 41198 800
rect 42154 0 42210 800
rect 43166 0 43222 800
rect 44178 0 44234 800
rect 45190 0 45246 800
rect 46202 0 46258 800
rect 47214 0 47270 800
rect 48226 0 48282 800
rect 49238 0 49294 800
rect 50250 0 50306 800
rect 51262 0 51318 800
rect 52274 0 52330 800
rect 53286 0 53342 800
rect 54298 0 54354 800
rect 55310 0 55366 800
rect 56322 0 56378 800
rect 57334 0 57390 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60370 0 60426 800
rect 61382 0 61438 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70490 0 70546 800
rect 71502 0 71558 800
rect 72514 0 72570 800
rect 73526 0 73582 800
rect 74538 0 74594 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77574 0 77630 800
rect 78586 0 78642 800
rect 79598 0 79654 800
rect 80610 0 80666 800
rect 81622 0 81678 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84658 0 84714 800
rect 85670 0 85726 800
rect 86682 0 86738 800
rect 87694 0 87750 800
rect 88706 0 88762 800
rect 89718 0 89774 800
rect 90730 0 90786 800
rect 91742 0 91798 800
rect 92754 0 92810 800
rect 93766 0 93822 800
rect 94778 0 94834 800
rect 95790 0 95846 800
rect 96802 0 96858 800
rect 97814 0 97870 800
rect 98826 0 98882 800
rect 99838 0 99894 800
rect 100850 0 100906 800
rect 101862 0 101918 800
rect 102874 0 102930 800
rect 103886 0 103942 800
rect 104898 0 104954 800
rect 105910 0 105966 800
rect 106922 0 106978 800
rect 107934 0 107990 800
rect 108946 0 109002 800
rect 109958 0 110014 800
rect 110970 0 111026 800
rect 111982 0 112038 800
rect 112994 0 113050 800
rect 114006 0 114062 800
rect 115018 0 115074 800
rect 116030 0 116086 800
rect 117042 0 117098 800
rect 118054 0 118110 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 121090 0 121146 800
rect 122102 0 122158 800
rect 123114 0 123170 800
rect 124126 0 124182 800
rect 125138 0 125194 800
rect 126150 0 126206 800
rect 127162 0 127218 800
rect 128174 0 128230 800
rect 129186 0 129242 800
<< obsm2 >>
rect 664 124144 13026 124200
rect 13194 124144 38970 124200
rect 39138 124144 64914 124200
rect 65082 124144 90858 124200
rect 91026 124144 116802 124200
rect 116970 124144 129240 124200
rect 664 856 129240 124144
rect 774 734 1618 856
rect 1786 734 2630 856
rect 2798 734 3642 856
rect 3810 734 4654 856
rect 4822 734 5666 856
rect 5834 734 6678 856
rect 6846 734 7690 856
rect 7858 734 8702 856
rect 8870 734 9714 856
rect 9882 734 10726 856
rect 10894 734 11738 856
rect 11906 734 12750 856
rect 12918 734 13762 856
rect 13930 734 14774 856
rect 14942 734 15786 856
rect 15954 734 16798 856
rect 16966 734 17810 856
rect 17978 734 18822 856
rect 18990 734 19834 856
rect 20002 734 20846 856
rect 21014 734 21858 856
rect 22026 734 22870 856
rect 23038 734 23882 856
rect 24050 734 24894 856
rect 25062 734 25906 856
rect 26074 734 26918 856
rect 27086 734 27930 856
rect 28098 734 28942 856
rect 29110 734 29954 856
rect 30122 734 30966 856
rect 31134 734 31978 856
rect 32146 734 32990 856
rect 33158 734 34002 856
rect 34170 734 35014 856
rect 35182 734 36026 856
rect 36194 734 37038 856
rect 37206 734 38050 856
rect 38218 734 39062 856
rect 39230 734 40074 856
rect 40242 734 41086 856
rect 41254 734 42098 856
rect 42266 734 43110 856
rect 43278 734 44122 856
rect 44290 734 45134 856
rect 45302 734 46146 856
rect 46314 734 47158 856
rect 47326 734 48170 856
rect 48338 734 49182 856
rect 49350 734 50194 856
rect 50362 734 51206 856
rect 51374 734 52218 856
rect 52386 734 53230 856
rect 53398 734 54242 856
rect 54410 734 55254 856
rect 55422 734 56266 856
rect 56434 734 57278 856
rect 57446 734 58290 856
rect 58458 734 59302 856
rect 59470 734 60314 856
rect 60482 734 61326 856
rect 61494 734 62338 856
rect 62506 734 63350 856
rect 63518 734 64362 856
rect 64530 734 65374 856
rect 65542 734 66386 856
rect 66554 734 67398 856
rect 67566 734 68410 856
rect 68578 734 69422 856
rect 69590 734 70434 856
rect 70602 734 71446 856
rect 71614 734 72458 856
rect 72626 734 73470 856
rect 73638 734 74482 856
rect 74650 734 75494 856
rect 75662 734 76506 856
rect 76674 734 77518 856
rect 77686 734 78530 856
rect 78698 734 79542 856
rect 79710 734 80554 856
rect 80722 734 81566 856
rect 81734 734 82578 856
rect 82746 734 83590 856
rect 83758 734 84602 856
rect 84770 734 85614 856
rect 85782 734 86626 856
rect 86794 734 87638 856
rect 87806 734 88650 856
rect 88818 734 89662 856
rect 89830 734 90674 856
rect 90842 734 91686 856
rect 91854 734 92698 856
rect 92866 734 93710 856
rect 93878 734 94722 856
rect 94890 734 95734 856
rect 95902 734 96746 856
rect 96914 734 97758 856
rect 97926 734 98770 856
rect 98938 734 99782 856
rect 99950 734 100794 856
rect 100962 734 101806 856
rect 101974 734 102818 856
rect 102986 734 103830 856
rect 103998 734 104842 856
rect 105010 734 105854 856
rect 106022 734 106866 856
rect 107034 734 107878 856
rect 108046 734 108890 856
rect 109058 734 109902 856
rect 110070 734 110914 856
rect 111082 734 111926 856
rect 112094 734 112938 856
rect 113106 734 113950 856
rect 114118 734 114962 856
rect 115130 734 115974 856
rect 116142 734 116986 856
rect 117154 734 117998 856
rect 118166 734 119010 856
rect 119178 734 120022 856
rect 120190 734 121034 856
rect 121202 734 122046 856
rect 122214 734 123058 856
rect 123226 734 124070 856
rect 124238 734 125082 856
rect 125250 734 126094 856
rect 126262 734 127106 856
rect 127274 734 128118 856
rect 128286 734 129130 856
<< metal3 >>
rect 129200 121048 130000 121168
rect 129200 116696 130000 116816
rect 0 114248 800 114368
rect 0 113432 800 113552
rect 0 112616 800 112736
rect 129200 112344 130000 112464
rect 0 111800 800 111920
rect 0 110984 800 111104
rect 0 110168 800 110288
rect 0 109352 800 109472
rect 0 108536 800 108656
rect 129200 107992 130000 108112
rect 0 107720 800 107840
rect 0 106904 800 107024
rect 0 106088 800 106208
rect 0 105272 800 105392
rect 0 104456 800 104576
rect 0 103640 800 103760
rect 129200 103640 130000 103760
rect 0 102824 800 102944
rect 0 102008 800 102128
rect 0 101192 800 101312
rect 0 100376 800 100496
rect 0 99560 800 99680
rect 129200 99288 130000 99408
rect 0 98744 800 98864
rect 0 97928 800 98048
rect 0 97112 800 97232
rect 0 96296 800 96416
rect 0 95480 800 95600
rect 129200 94936 130000 95056
rect 0 94664 800 94784
rect 0 93848 800 93968
rect 0 93032 800 93152
rect 0 92216 800 92336
rect 0 91400 800 91520
rect 0 90584 800 90704
rect 129200 90584 130000 90704
rect 0 89768 800 89888
rect 0 88952 800 89072
rect 0 88136 800 88256
rect 0 87320 800 87440
rect 0 86504 800 86624
rect 129200 86232 130000 86352
rect 0 85688 800 85808
rect 0 84872 800 84992
rect 0 84056 800 84176
rect 0 83240 800 83360
rect 0 82424 800 82544
rect 129200 81880 130000 82000
rect 0 81608 800 81728
rect 0 80792 800 80912
rect 0 79976 800 80096
rect 0 79160 800 79280
rect 0 78344 800 78464
rect 0 77528 800 77648
rect 129200 77528 130000 77648
rect 0 76712 800 76832
rect 0 75896 800 76016
rect 0 75080 800 75200
rect 0 74264 800 74384
rect 0 73448 800 73568
rect 129200 73176 130000 73296
rect 0 72632 800 72752
rect 0 71816 800 71936
rect 0 71000 800 71120
rect 0 70184 800 70304
rect 0 69368 800 69488
rect 129200 68824 130000 68944
rect 0 68552 800 68672
rect 0 67736 800 67856
rect 0 66920 800 67040
rect 0 66104 800 66224
rect 0 65288 800 65408
rect 0 64472 800 64592
rect 129200 64472 130000 64592
rect 0 63656 800 63776
rect 0 62840 800 62960
rect 0 62024 800 62144
rect 0 61208 800 61328
rect 0 60392 800 60512
rect 129200 60120 130000 60240
rect 0 59576 800 59696
rect 0 58760 800 58880
rect 0 57944 800 58064
rect 0 57128 800 57248
rect 0 56312 800 56432
rect 129200 55768 130000 55888
rect 0 55496 800 55616
rect 0 54680 800 54800
rect 0 53864 800 53984
rect 0 53048 800 53168
rect 0 52232 800 52352
rect 0 51416 800 51536
rect 129200 51416 130000 51536
rect 0 50600 800 50720
rect 0 49784 800 49904
rect 0 48968 800 49088
rect 0 48152 800 48272
rect 0 47336 800 47456
rect 129200 47064 130000 47184
rect 0 46520 800 46640
rect 0 45704 800 45824
rect 0 44888 800 45008
rect 0 44072 800 44192
rect 0 43256 800 43376
rect 129200 42712 130000 42832
rect 0 42440 800 42560
rect 0 41624 800 41744
rect 0 40808 800 40928
rect 0 39992 800 40112
rect 0 39176 800 39296
rect 0 38360 800 38480
rect 129200 38360 130000 38480
rect 0 37544 800 37664
rect 0 36728 800 36848
rect 0 35912 800 36032
rect 0 35096 800 35216
rect 0 34280 800 34400
rect 129200 34008 130000 34128
rect 0 33464 800 33584
rect 0 32648 800 32768
rect 0 31832 800 31952
rect 0 31016 800 31136
rect 0 30200 800 30320
rect 129200 29656 130000 29776
rect 0 29384 800 29504
rect 0 28568 800 28688
rect 0 27752 800 27872
rect 0 26936 800 27056
rect 0 26120 800 26240
rect 0 25304 800 25424
rect 129200 25304 130000 25424
rect 0 24488 800 24608
rect 0 23672 800 23792
rect 0 22856 800 22976
rect 0 22040 800 22160
rect 0 21224 800 21344
rect 129200 20952 130000 21072
rect 0 20408 800 20528
rect 0 19592 800 19712
rect 0 18776 800 18896
rect 0 17960 800 18080
rect 0 17144 800 17264
rect 129200 16600 130000 16720
rect 0 16328 800 16448
rect 0 15512 800 15632
rect 0 14696 800 14816
rect 0 13880 800 14000
rect 0 13064 800 13184
rect 0 12248 800 12368
rect 129200 12248 130000 12368
rect 0 11432 800 11552
rect 0 10616 800 10736
rect 129200 7896 130000 8016
rect 129200 3544 130000 3664
<< obsm3 >>
rect 798 121248 129200 122433
rect 798 120968 129120 121248
rect 798 116896 129200 120968
rect 798 116616 129120 116896
rect 798 114448 129200 116616
rect 880 114168 129200 114448
rect 798 113632 129200 114168
rect 880 113352 129200 113632
rect 798 112816 129200 113352
rect 880 112544 129200 112816
rect 880 112536 129120 112544
rect 798 112264 129120 112536
rect 798 112000 129200 112264
rect 880 111720 129200 112000
rect 798 111184 129200 111720
rect 880 110904 129200 111184
rect 798 110368 129200 110904
rect 880 110088 129200 110368
rect 798 109552 129200 110088
rect 880 109272 129200 109552
rect 798 108736 129200 109272
rect 880 108456 129200 108736
rect 798 108192 129200 108456
rect 798 107920 129120 108192
rect 880 107912 129120 107920
rect 880 107640 129200 107912
rect 798 107104 129200 107640
rect 880 106824 129200 107104
rect 798 106288 129200 106824
rect 880 106008 129200 106288
rect 798 105472 129200 106008
rect 880 105192 129200 105472
rect 798 104656 129200 105192
rect 880 104376 129200 104656
rect 798 103840 129200 104376
rect 880 103560 129120 103840
rect 798 103024 129200 103560
rect 880 102744 129200 103024
rect 798 102208 129200 102744
rect 880 101928 129200 102208
rect 798 101392 129200 101928
rect 880 101112 129200 101392
rect 798 100576 129200 101112
rect 880 100296 129200 100576
rect 798 99760 129200 100296
rect 880 99488 129200 99760
rect 880 99480 129120 99488
rect 798 99208 129120 99480
rect 798 98944 129200 99208
rect 880 98664 129200 98944
rect 798 98128 129200 98664
rect 880 97848 129200 98128
rect 798 97312 129200 97848
rect 880 97032 129200 97312
rect 798 96496 129200 97032
rect 880 96216 129200 96496
rect 798 95680 129200 96216
rect 880 95400 129200 95680
rect 798 95136 129200 95400
rect 798 94864 129120 95136
rect 880 94856 129120 94864
rect 880 94584 129200 94856
rect 798 94048 129200 94584
rect 880 93768 129200 94048
rect 798 93232 129200 93768
rect 880 92952 129200 93232
rect 798 92416 129200 92952
rect 880 92136 129200 92416
rect 798 91600 129200 92136
rect 880 91320 129200 91600
rect 798 90784 129200 91320
rect 880 90504 129120 90784
rect 798 89968 129200 90504
rect 880 89688 129200 89968
rect 798 89152 129200 89688
rect 880 88872 129200 89152
rect 798 88336 129200 88872
rect 880 88056 129200 88336
rect 798 87520 129200 88056
rect 880 87240 129200 87520
rect 798 86704 129200 87240
rect 880 86432 129200 86704
rect 880 86424 129120 86432
rect 798 86152 129120 86424
rect 798 85888 129200 86152
rect 880 85608 129200 85888
rect 798 85072 129200 85608
rect 880 84792 129200 85072
rect 798 84256 129200 84792
rect 880 83976 129200 84256
rect 798 83440 129200 83976
rect 880 83160 129200 83440
rect 798 82624 129200 83160
rect 880 82344 129200 82624
rect 798 82080 129200 82344
rect 798 81808 129120 82080
rect 880 81800 129120 81808
rect 880 81528 129200 81800
rect 798 80992 129200 81528
rect 880 80712 129200 80992
rect 798 80176 129200 80712
rect 880 79896 129200 80176
rect 798 79360 129200 79896
rect 880 79080 129200 79360
rect 798 78544 129200 79080
rect 880 78264 129200 78544
rect 798 77728 129200 78264
rect 880 77448 129120 77728
rect 798 76912 129200 77448
rect 880 76632 129200 76912
rect 798 76096 129200 76632
rect 880 75816 129200 76096
rect 798 75280 129200 75816
rect 880 75000 129200 75280
rect 798 74464 129200 75000
rect 880 74184 129200 74464
rect 798 73648 129200 74184
rect 880 73376 129200 73648
rect 880 73368 129120 73376
rect 798 73096 129120 73368
rect 798 72832 129200 73096
rect 880 72552 129200 72832
rect 798 72016 129200 72552
rect 880 71736 129200 72016
rect 798 71200 129200 71736
rect 880 70920 129200 71200
rect 798 70384 129200 70920
rect 880 70104 129200 70384
rect 798 69568 129200 70104
rect 880 69288 129200 69568
rect 798 69024 129200 69288
rect 798 68752 129120 69024
rect 880 68744 129120 68752
rect 880 68472 129200 68744
rect 798 67936 129200 68472
rect 880 67656 129200 67936
rect 798 67120 129200 67656
rect 880 66840 129200 67120
rect 798 66304 129200 66840
rect 880 66024 129200 66304
rect 798 65488 129200 66024
rect 880 65208 129200 65488
rect 798 64672 129200 65208
rect 880 64392 129120 64672
rect 798 63856 129200 64392
rect 880 63576 129200 63856
rect 798 63040 129200 63576
rect 880 62760 129200 63040
rect 798 62224 129200 62760
rect 880 61944 129200 62224
rect 798 61408 129200 61944
rect 880 61128 129200 61408
rect 798 60592 129200 61128
rect 880 60320 129200 60592
rect 880 60312 129120 60320
rect 798 60040 129120 60312
rect 798 59776 129200 60040
rect 880 59496 129200 59776
rect 798 58960 129200 59496
rect 880 58680 129200 58960
rect 798 58144 129200 58680
rect 880 57864 129200 58144
rect 798 57328 129200 57864
rect 880 57048 129200 57328
rect 798 56512 129200 57048
rect 880 56232 129200 56512
rect 798 55968 129200 56232
rect 798 55696 129120 55968
rect 880 55688 129120 55696
rect 880 55416 129200 55688
rect 798 54880 129200 55416
rect 880 54600 129200 54880
rect 798 54064 129200 54600
rect 880 53784 129200 54064
rect 798 53248 129200 53784
rect 880 52968 129200 53248
rect 798 52432 129200 52968
rect 880 52152 129200 52432
rect 798 51616 129200 52152
rect 880 51336 129120 51616
rect 798 50800 129200 51336
rect 880 50520 129200 50800
rect 798 49984 129200 50520
rect 880 49704 129200 49984
rect 798 49168 129200 49704
rect 880 48888 129200 49168
rect 798 48352 129200 48888
rect 880 48072 129200 48352
rect 798 47536 129200 48072
rect 880 47264 129200 47536
rect 880 47256 129120 47264
rect 798 46984 129120 47256
rect 798 46720 129200 46984
rect 880 46440 129200 46720
rect 798 45904 129200 46440
rect 880 45624 129200 45904
rect 798 45088 129200 45624
rect 880 44808 129200 45088
rect 798 44272 129200 44808
rect 880 43992 129200 44272
rect 798 43456 129200 43992
rect 880 43176 129200 43456
rect 798 42912 129200 43176
rect 798 42640 129120 42912
rect 880 42632 129120 42640
rect 880 42360 129200 42632
rect 798 41824 129200 42360
rect 880 41544 129200 41824
rect 798 41008 129200 41544
rect 880 40728 129200 41008
rect 798 40192 129200 40728
rect 880 39912 129200 40192
rect 798 39376 129200 39912
rect 880 39096 129200 39376
rect 798 38560 129200 39096
rect 880 38280 129120 38560
rect 798 37744 129200 38280
rect 880 37464 129200 37744
rect 798 36928 129200 37464
rect 880 36648 129200 36928
rect 798 36112 129200 36648
rect 880 35832 129200 36112
rect 798 35296 129200 35832
rect 880 35016 129200 35296
rect 798 34480 129200 35016
rect 880 34208 129200 34480
rect 880 34200 129120 34208
rect 798 33928 129120 34200
rect 798 33664 129200 33928
rect 880 33384 129200 33664
rect 798 32848 129200 33384
rect 880 32568 129200 32848
rect 798 32032 129200 32568
rect 880 31752 129200 32032
rect 798 31216 129200 31752
rect 880 30936 129200 31216
rect 798 30400 129200 30936
rect 880 30120 129200 30400
rect 798 29856 129200 30120
rect 798 29584 129120 29856
rect 880 29576 129120 29584
rect 880 29304 129200 29576
rect 798 28768 129200 29304
rect 880 28488 129200 28768
rect 798 27952 129200 28488
rect 880 27672 129200 27952
rect 798 27136 129200 27672
rect 880 26856 129200 27136
rect 798 26320 129200 26856
rect 880 26040 129200 26320
rect 798 25504 129200 26040
rect 880 25224 129120 25504
rect 798 24688 129200 25224
rect 880 24408 129200 24688
rect 798 23872 129200 24408
rect 880 23592 129200 23872
rect 798 23056 129200 23592
rect 880 22776 129200 23056
rect 798 22240 129200 22776
rect 880 21960 129200 22240
rect 798 21424 129200 21960
rect 880 21152 129200 21424
rect 880 21144 129120 21152
rect 798 20872 129120 21144
rect 798 20608 129200 20872
rect 880 20328 129200 20608
rect 798 19792 129200 20328
rect 880 19512 129200 19792
rect 798 18976 129200 19512
rect 880 18696 129200 18976
rect 798 18160 129200 18696
rect 880 17880 129200 18160
rect 798 17344 129200 17880
rect 880 17064 129200 17344
rect 798 16800 129200 17064
rect 798 16528 129120 16800
rect 880 16520 129120 16528
rect 880 16248 129200 16520
rect 798 15712 129200 16248
rect 880 15432 129200 15712
rect 798 14896 129200 15432
rect 880 14616 129200 14896
rect 798 14080 129200 14616
rect 880 13800 129200 14080
rect 798 13264 129200 13800
rect 880 12984 129200 13264
rect 798 12448 129200 12984
rect 880 12168 129120 12448
rect 798 11632 129200 12168
rect 880 11352 129200 11632
rect 798 10816 129200 11352
rect 880 10536 129200 10816
rect 798 8096 129200 10536
rect 798 7816 129120 8096
rect 798 3744 129200 7816
rect 798 3464 129120 3744
rect 798 2143 129200 3464
<< metal4 >>
rect 4208 2128 4528 122448
rect 19568 2128 19888 122448
rect 34928 2128 35248 122448
rect 50288 2128 50608 122448
rect 65648 2128 65968 122448
rect 81008 2128 81328 122448
rect 96368 2128 96688 122448
rect 111728 2128 112048 122448
rect 127088 2128 127408 122448
<< obsm4 >>
rect 1715 2347 4128 122093
rect 4608 2347 19488 122093
rect 19968 2347 34848 122093
rect 35328 2347 50208 122093
rect 50688 2347 65568 122093
rect 66048 2347 80928 122093
rect 81408 2347 96288 122093
rect 96768 2347 111648 122093
rect 112128 2347 127008 122093
rect 127488 2347 128005 122093
<< labels >>
rlabel metal2 s 662 0 718 800 6 cache_entry[0]
port 1 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 cache_entry[100]
port 2 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 cache_entry[101]
port 3 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 cache_entry[102]
port 4 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 cache_entry[103]
port 5 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 cache_entry[104]
port 6 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 cache_entry[105]
port 7 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 cache_entry[106]
port 8 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 cache_entry[107]
port 9 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 cache_entry[108]
port 10 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 cache_entry[109]
port 11 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 cache_entry[10]
port 12 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 cache_entry[110]
port 13 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 cache_entry[111]
port 14 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 cache_entry[112]
port 15 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 cache_entry[113]
port 16 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 cache_entry[114]
port 17 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 cache_entry[115]
port 18 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 cache_entry[116]
port 19 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 cache_entry[117]
port 20 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 cache_entry[118]
port 21 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 cache_entry[119]
port 22 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 cache_entry[11]
port 23 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 cache_entry[120]
port 24 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 cache_entry[121]
port 25 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 cache_entry[122]
port 26 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 cache_entry[123]
port 27 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 cache_entry[124]
port 28 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 cache_entry[125]
port 29 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 cache_entry[126]
port 30 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 cache_entry[127]
port 31 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 cache_entry[12]
port 32 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 cache_entry[13]
port 33 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 cache_entry[14]
port 34 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 cache_entry[15]
port 35 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 cache_entry[16]
port 36 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 cache_entry[17]
port 37 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 cache_entry[18]
port 38 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 cache_entry[19]
port 39 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 cache_entry[1]
port 40 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 cache_entry[20]
port 41 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 cache_entry[21]
port 42 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 cache_entry[22]
port 43 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 cache_entry[23]
port 44 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 cache_entry[24]
port 45 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 cache_entry[25]
port 46 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 cache_entry[26]
port 47 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 cache_entry[27]
port 48 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 cache_entry[28]
port 49 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 cache_entry[29]
port 50 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 cache_entry[2]
port 51 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 cache_entry[30]
port 52 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 cache_entry[31]
port 53 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 cache_entry[32]
port 54 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 cache_entry[33]
port 55 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 cache_entry[34]
port 56 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 cache_entry[35]
port 57 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 cache_entry[36]
port 58 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 cache_entry[37]
port 59 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 cache_entry[38]
port 60 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 cache_entry[39]
port 61 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 cache_entry[3]
port 62 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 cache_entry[40]
port 63 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 cache_entry[41]
port 64 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 cache_entry[42]
port 65 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 cache_entry[43]
port 66 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 cache_entry[44]
port 67 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 cache_entry[45]
port 68 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 cache_entry[46]
port 69 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 cache_entry[47]
port 70 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 cache_entry[48]
port 71 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 cache_entry[49]
port 72 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 cache_entry[4]
port 73 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 cache_entry[50]
port 74 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 cache_entry[51]
port 75 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 cache_entry[52]
port 76 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 cache_entry[53]
port 77 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 cache_entry[54]
port 78 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 cache_entry[55]
port 79 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 cache_entry[56]
port 80 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 cache_entry[57]
port 81 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 cache_entry[58]
port 82 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 cache_entry[59]
port 83 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 cache_entry[5]
port 84 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 cache_entry[60]
port 85 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 cache_entry[61]
port 86 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 cache_entry[62]
port 87 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 cache_entry[63]
port 88 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 cache_entry[64]
port 89 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 cache_entry[65]
port 90 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 cache_entry[66]
port 91 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 cache_entry[67]
port 92 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 cache_entry[68]
port 93 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 cache_entry[69]
port 94 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 cache_entry[6]
port 95 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 cache_entry[70]
port 96 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 cache_entry[71]
port 97 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 cache_entry[72]
port 98 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 cache_entry[73]
port 99 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 cache_entry[74]
port 100 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 cache_entry[75]
port 101 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 cache_entry[76]
port 102 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 cache_entry[77]
port 103 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 cache_entry[78]
port 104 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 cache_entry[79]
port 105 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 cache_entry[7]
port 106 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 cache_entry[80]
port 107 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 cache_entry[81]
port 108 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 cache_entry[82]
port 109 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 cache_entry[83]
port 110 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 cache_entry[84]
port 111 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 cache_entry[85]
port 112 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 cache_entry[86]
port 113 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 cache_entry[87]
port 114 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 cache_entry[88]
port 115 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 cache_entry[89]
port 116 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 cache_entry[8]
port 117 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 cache_entry[90]
port 118 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 cache_entry[91]
port 119 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 cache_entry[92]
port 120 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 cache_entry[93]
port 121 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 cache_entry[94]
port 122 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 cache_entry[95]
port 123 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 cache_entry[96]
port 124 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 cache_entry[97]
port 125 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 cache_entry[98]
port 126 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 cache_entry[99]
port 127 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 cache_entry[9]
port 128 nsew signal output
rlabel metal2 s 90914 124200 90970 125000 6 cache_hit
port 129 nsew signal output
rlabel metal2 s 13082 124200 13138 125000 6 clk
port 130 nsew signal input
rlabel metal3 s 129200 3544 130000 3664 6 curr_PC[0]
port 131 nsew signal input
rlabel metal3 s 129200 47064 130000 47184 6 curr_PC[10]
port 132 nsew signal input
rlabel metal3 s 129200 51416 130000 51536 6 curr_PC[11]
port 133 nsew signal input
rlabel metal3 s 129200 55768 130000 55888 6 curr_PC[12]
port 134 nsew signal input
rlabel metal3 s 129200 60120 130000 60240 6 curr_PC[13]
port 135 nsew signal input
rlabel metal3 s 129200 64472 130000 64592 6 curr_PC[14]
port 136 nsew signal input
rlabel metal3 s 129200 68824 130000 68944 6 curr_PC[15]
port 137 nsew signal input
rlabel metal3 s 129200 73176 130000 73296 6 curr_PC[16]
port 138 nsew signal input
rlabel metal3 s 129200 77528 130000 77648 6 curr_PC[17]
port 139 nsew signal input
rlabel metal3 s 129200 81880 130000 82000 6 curr_PC[18]
port 140 nsew signal input
rlabel metal3 s 129200 86232 130000 86352 6 curr_PC[19]
port 141 nsew signal input
rlabel metal3 s 129200 7896 130000 8016 6 curr_PC[1]
port 142 nsew signal input
rlabel metal3 s 129200 90584 130000 90704 6 curr_PC[20]
port 143 nsew signal input
rlabel metal3 s 129200 94936 130000 95056 6 curr_PC[21]
port 144 nsew signal input
rlabel metal3 s 129200 99288 130000 99408 6 curr_PC[22]
port 145 nsew signal input
rlabel metal3 s 129200 103640 130000 103760 6 curr_PC[23]
port 146 nsew signal input
rlabel metal3 s 129200 107992 130000 108112 6 curr_PC[24]
port 147 nsew signal input
rlabel metal3 s 129200 112344 130000 112464 6 curr_PC[25]
port 148 nsew signal input
rlabel metal3 s 129200 116696 130000 116816 6 curr_PC[26]
port 149 nsew signal input
rlabel metal3 s 129200 121048 130000 121168 6 curr_PC[27]
port 150 nsew signal input
rlabel metal3 s 129200 12248 130000 12368 6 curr_PC[2]
port 151 nsew signal input
rlabel metal3 s 129200 16600 130000 16720 6 curr_PC[3]
port 152 nsew signal input
rlabel metal3 s 129200 20952 130000 21072 6 curr_PC[4]
port 153 nsew signal input
rlabel metal3 s 129200 25304 130000 25424 6 curr_PC[5]
port 154 nsew signal input
rlabel metal3 s 129200 29656 130000 29776 6 curr_PC[6]
port 155 nsew signal input
rlabel metal3 s 129200 34008 130000 34128 6 curr_PC[7]
port 156 nsew signal input
rlabel metal3 s 129200 38360 130000 38480 6 curr_PC[8]
port 157 nsew signal input
rlabel metal3 s 129200 42712 130000 42832 6 curr_PC[9]
port 158 nsew signal input
rlabel metal2 s 116858 124200 116914 125000 6 entry_valid
port 159 nsew signal input
rlabel metal2 s 64970 124200 65026 125000 6 invalidate
port 160 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 new_entry[0]
port 161 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 new_entry[100]
port 162 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 new_entry[101]
port 163 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 new_entry[102]
port 164 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 new_entry[103]
port 165 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 new_entry[104]
port 166 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 new_entry[105]
port 167 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 new_entry[106]
port 168 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 new_entry[107]
port 169 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 new_entry[108]
port 170 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 new_entry[109]
port 171 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 new_entry[10]
port 172 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 new_entry[110]
port 173 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 new_entry[111]
port 174 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 new_entry[112]
port 175 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 new_entry[113]
port 176 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 new_entry[114]
port 177 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 new_entry[115]
port 178 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 new_entry[116]
port 179 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 new_entry[117]
port 180 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 new_entry[118]
port 181 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 new_entry[119]
port 182 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 new_entry[11]
port 183 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 new_entry[120]
port 184 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 new_entry[121]
port 185 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 new_entry[122]
port 186 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 new_entry[123]
port 187 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 new_entry[124]
port 188 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 new_entry[125]
port 189 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 new_entry[126]
port 190 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 new_entry[127]
port 191 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 new_entry[12]
port 192 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 new_entry[13]
port 193 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 new_entry[14]
port 194 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 new_entry[15]
port 195 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 new_entry[16]
port 196 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 new_entry[17]
port 197 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 new_entry[18]
port 198 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 new_entry[19]
port 199 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 new_entry[1]
port 200 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 new_entry[20]
port 201 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 new_entry[21]
port 202 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 new_entry[22]
port 203 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 new_entry[23]
port 204 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 new_entry[24]
port 205 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 new_entry[25]
port 206 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 new_entry[26]
port 207 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 new_entry[27]
port 208 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 new_entry[28]
port 209 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 new_entry[29]
port 210 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 new_entry[2]
port 211 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 new_entry[30]
port 212 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 new_entry[31]
port 213 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 new_entry[32]
port 214 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 new_entry[33]
port 215 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 new_entry[34]
port 216 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 new_entry[35]
port 217 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 new_entry[36]
port 218 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 new_entry[37]
port 219 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 new_entry[38]
port 220 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 new_entry[39]
port 221 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 new_entry[3]
port 222 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 new_entry[40]
port 223 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 new_entry[41]
port 224 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 new_entry[42]
port 225 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 new_entry[43]
port 226 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 new_entry[44]
port 227 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 new_entry[45]
port 228 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 new_entry[46]
port 229 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 new_entry[47]
port 230 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 new_entry[48]
port 231 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 new_entry[49]
port 232 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 new_entry[4]
port 233 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 new_entry[50]
port 234 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 new_entry[51]
port 235 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 new_entry[52]
port 236 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 new_entry[53]
port 237 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 new_entry[54]
port 238 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 new_entry[55]
port 239 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 new_entry[56]
port 240 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 new_entry[57]
port 241 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 new_entry[58]
port 242 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 new_entry[59]
port 243 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 new_entry[5]
port 244 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 new_entry[60]
port 245 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 new_entry[61]
port 246 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 new_entry[62]
port 247 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 new_entry[63]
port 248 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 new_entry[64]
port 249 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 new_entry[65]
port 250 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 new_entry[66]
port 251 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 new_entry[67]
port 252 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 new_entry[68]
port 253 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 new_entry[69]
port 254 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 new_entry[6]
port 255 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 new_entry[70]
port 256 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 new_entry[71]
port 257 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 new_entry[72]
port 258 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 new_entry[73]
port 259 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 new_entry[74]
port 260 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 new_entry[75]
port 261 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 new_entry[76]
port 262 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 new_entry[77]
port 263 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 new_entry[78]
port 264 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 new_entry[79]
port 265 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 new_entry[7]
port 266 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 new_entry[80]
port 267 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 new_entry[81]
port 268 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 new_entry[82]
port 269 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 new_entry[83]
port 270 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 new_entry[84]
port 271 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 new_entry[85]
port 272 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 new_entry[86]
port 273 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 new_entry[87]
port 274 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 new_entry[88]
port 275 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 new_entry[89]
port 276 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 new_entry[8]
port 277 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 new_entry[90]
port 278 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 new_entry[91]
port 279 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 new_entry[92]
port 280 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 new_entry[93]
port 281 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 new_entry[94]
port 282 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 new_entry[95]
port 283 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 new_entry[96]
port 284 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 new_entry[97]
port 285 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 new_entry[98]
port 286 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 new_entry[99]
port 287 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 new_entry[9]
port 288 nsew signal input
rlabel metal2 s 39026 124200 39082 125000 6 rst
port 289 nsew signal input
rlabel metal4 s 4208 2128 4528 122448 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 122448 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 122448 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 122448 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 122448 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 122448 6 vssd1
port 291 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 122448 6 vssd1
port 291 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 122448 6 vssd1
port 291 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 122448 6 vssd1
port 291 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 130000 125000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 62040570
string GDS_FILE /run/media/tholin/8a6b8802-051e-45a8-8492-771202e4c08a/ci2406-rej-pommedeterrible-tholin/openlane/icache/runs/24_05_30_20_24/results/signoff/icache.magic.gds
string GDS_START 656218
<< end >>

