// This is the unpowered netlist.
module execution_unit (busy,
    dest_pred_val,
    int_return,
    is_load,
    is_store,
    pred_val,
    rst,
    sign_extend,
    take_branch,
    wb_clk_i,
    curr_PC,
    dest_idx,
    dest_mask,
    dest_pred,
    dest_val,
    instruction,
    loadstore_address,
    loadstore_dest,
    loadstore_size,
    new_PC,
    pred_idx,
    reg1_idx,
    reg1_val,
    reg2_idx,
    reg2_val);
 output busy;
 output dest_pred_val;
 output int_return;
 output is_load;
 output is_store;
 input pred_val;
 input rst;
 output sign_extend;
 output take_branch;
 input wb_clk_i;
 input [27:0] curr_PC;
 output [5:0] dest_idx;
 output [1:0] dest_mask;
 output [2:0] dest_pred;
 output [31:0] dest_val;
 input [41:0] instruction;
 output [31:0] loadstore_address;
 output [5:0] loadstore_dest;
 output [1:0] loadstore_size;
 output [27:0] new_PC;
 output [2:0] pred_idx;
 output [5:0] reg1_idx;
 input [31:0] reg1_val;
 output [5:0] reg2_idx;
 input [31:0] reg2_val;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire busy_l;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire div_complete;
 wire \div_counter[0] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_res[0] ;
 wire \div_res[10] ;
 wire \div_res[11] ;
 wire \div_res[12] ;
 wire \div_res[13] ;
 wire \div_res[14] ;
 wire \div_res[15] ;
 wire \div_res[16] ;
 wire \div_res[17] ;
 wire \div_res[18] ;
 wire \div_res[19] ;
 wire \div_res[1] ;
 wire \div_res[20] ;
 wire \div_res[21] ;
 wire \div_res[22] ;
 wire \div_res[23] ;
 wire \div_res[24] ;
 wire \div_res[25] ;
 wire \div_res[26] ;
 wire \div_res[27] ;
 wire \div_res[28] ;
 wire \div_res[29] ;
 wire \div_res[2] ;
 wire \div_res[30] ;
 wire \div_res[31] ;
 wire \div_res[3] ;
 wire \div_res[4] ;
 wire \div_res[5] ;
 wire \div_res[6] ;
 wire \div_res[7] ;
 wire \div_res[8] ;
 wire \div_res[9] ;
 wire \div_shifter[0] ;
 wire \div_shifter[10] ;
 wire \div_shifter[11] ;
 wire \div_shifter[12] ;
 wire \div_shifter[13] ;
 wire \div_shifter[14] ;
 wire \div_shifter[15] ;
 wire \div_shifter[16] ;
 wire \div_shifter[17] ;
 wire \div_shifter[18] ;
 wire \div_shifter[19] ;
 wire \div_shifter[1] ;
 wire \div_shifter[20] ;
 wire \div_shifter[21] ;
 wire \div_shifter[22] ;
 wire \div_shifter[23] ;
 wire \div_shifter[24] ;
 wire \div_shifter[25] ;
 wire \div_shifter[26] ;
 wire \div_shifter[27] ;
 wire \div_shifter[28] ;
 wire \div_shifter[29] ;
 wire \div_shifter[2] ;
 wire \div_shifter[30] ;
 wire \div_shifter[31] ;
 wire \div_shifter[32] ;
 wire \div_shifter[33] ;
 wire \div_shifter[34] ;
 wire \div_shifter[35] ;
 wire \div_shifter[36] ;
 wire \div_shifter[37] ;
 wire \div_shifter[38] ;
 wire \div_shifter[39] ;
 wire \div_shifter[3] ;
 wire \div_shifter[40] ;
 wire \div_shifter[41] ;
 wire \div_shifter[42] ;
 wire \div_shifter[43] ;
 wire \div_shifter[44] ;
 wire \div_shifter[45] ;
 wire \div_shifter[46] ;
 wire \div_shifter[47] ;
 wire \div_shifter[48] ;
 wire \div_shifter[49] ;
 wire \div_shifter[4] ;
 wire \div_shifter[50] ;
 wire \div_shifter[51] ;
 wire \div_shifter[52] ;
 wire \div_shifter[53] ;
 wire \div_shifter[54] ;
 wire \div_shifter[55] ;
 wire \div_shifter[56] ;
 wire \div_shifter[57] ;
 wire \div_shifter[58] ;
 wire \div_shifter[59] ;
 wire \div_shifter[5] ;
 wire \div_shifter[60] ;
 wire \div_shifter[61] ;
 wire \div_shifter[62] ;
 wire \div_shifter[63] ;
 wire \div_shifter[6] ;
 wire \div_shifter[7] ;
 wire \div_shifter[8] ;
 wire \div_shifter[9] ;
 wire divi1_sign;
 wire \divi2_l[0] ;
 wire \divi2_l[10] ;
 wire \divi2_l[11] ;
 wire \divi2_l[12] ;
 wire \divi2_l[13] ;
 wire \divi2_l[14] ;
 wire \divi2_l[15] ;
 wire \divi2_l[16] ;
 wire \divi2_l[17] ;
 wire \divi2_l[18] ;
 wire \divi2_l[19] ;
 wire \divi2_l[1] ;
 wire \divi2_l[20] ;
 wire \divi2_l[21] ;
 wire \divi2_l[22] ;
 wire \divi2_l[23] ;
 wire \divi2_l[24] ;
 wire \divi2_l[25] ;
 wire \divi2_l[26] ;
 wire \divi2_l[27] ;
 wire \divi2_l[28] ;
 wire \divi2_l[29] ;
 wire \divi2_l[2] ;
 wire \divi2_l[30] ;
 wire \divi2_l[31] ;
 wire \divi2_l[3] ;
 wire \divi2_l[4] ;
 wire \divi2_l[5] ;
 wire \divi2_l[6] ;
 wire \divi2_l[7] ;
 wire \divi2_l[8] ;
 wire \divi2_l[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(reg1_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(reg1_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(reg1_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(reg1_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(reg1_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(reg1_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(reg1_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(reg1_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(reg1_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(reg1_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(reg1_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(reg1_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(reg1_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(reg1_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(reg2_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(reg2_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(reg2_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(reg2_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(reg2_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(reg2_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(reg2_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(reg2_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(reg2_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(reg2_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(reg2_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04209_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(reg2_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(reg2_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(reg2_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(reg2_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(reg2_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(reg2_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(reg2_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(reg2_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(reg2_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(reg2_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(reg2_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(reg2_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(reg2_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(reg2_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(reg2_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(reg2_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(instruction[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(instruction[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(reg1_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(reg1_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(reg1_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(reg1_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(reg1_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(reg1_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(reg1_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(reg1_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(reg1_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(reg1_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(reg1_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06553__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06555__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06557__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__C1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__B (.DIODE(_04764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__B (.DIODE(_04764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06573__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__A2 (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__B (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A_N (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__B (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__A_N (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__B (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__B (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__A_N (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__B (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__B (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__B (.DIODE(_05132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A_N (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__B (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__B (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06606__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__A2_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__B (.DIODE(_05284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06615__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__B (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__B (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__A (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__B (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__B (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A2_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__B (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__B (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__B (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06650__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06652__B (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06653__B (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__B (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06657__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__A_N (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__B (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__B (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__B (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A2_N (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__B1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__B (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06688__A2_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A2_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__A2 (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__B (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__B (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A3 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__B (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__B (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__B (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06707__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06707__A3 (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__A3 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__B (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__A3 (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06724__A3 (.DIODE(_05284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__A3 (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A3 (.DIODE(_05132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__A3 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__A3 (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__C1 (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__D1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__C_N (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__B1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__B1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A3 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A3 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__A3 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A3 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06773__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06773__A3 (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A3 (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__B (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__B (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A3 (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__A3 (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__B (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__B (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__B (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__A_N (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__A_N (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A_N (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A_N (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__B (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__B (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__B (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__B (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__B (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__B (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06840__B (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A1 (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A2 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__D (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A1 (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__B (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__B (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__B (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__C (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__B (.DIODE(_04618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A2 (.DIODE(_04764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__C1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A2 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A3 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A3 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A4 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__B (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__A (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__B (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__C (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__D (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__B (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__C (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__D (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A2 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A3 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__B (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__C1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__B1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__C1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__A (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__C (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__D (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__B (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__B (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A3 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__B (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__C_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__C_N (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__B (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__B (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__B (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__C (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__C (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__D (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A1 (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B1 (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__B (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__B (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A1 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__C1 (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__C1 (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A2 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__B1 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__B (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__B (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__C (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__C (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__C (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__D (.DIODE(_00218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__B (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__A2 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__A3 (.DIODE(_00218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__B (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__B (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__B (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__B (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__B (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__C_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B2 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__B (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__B (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__A_N (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__A (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__B (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__A (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__A1 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__B (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__B (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__A (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A1 (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A1 (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A2 (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A2 (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A3 (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A_N (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A2 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__A (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__B (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__B (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A1 (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A1 (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__B (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__B (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__B (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A1 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B (.DIODE(_00432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B1 (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B (.DIODE(_00432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__C_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__B (.DIODE(_00432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__C (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A (.DIODE(_00438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__B (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A2 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A2 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__B (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__B1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__B1 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B1 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07436__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07436__B1 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__A2 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__B2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__B2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B (.DIODE(_00657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__B1 (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__B1 (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__D1 (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__A3 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__A4 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A1 (.DIODE(_00438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__B (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__A1 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__A2 (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A1 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__B1 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__B2 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__B1 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B2 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A1 (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B2 (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A1 (.DIODE(_00438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A1 (.DIODE(_00205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A1 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A2 (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__C (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B2 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A1 (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A (.DIODE(_00173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B1 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A2 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B1 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B2 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(_00241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A2 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__B (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07853__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__A_N (.DIODE(_00985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__B (.DIODE(_00985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A1 (.DIODE(_00241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A2 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__B1 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07867__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__B1 (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__A1 (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A2 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B1 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B2 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A2 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A1 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A2 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B1 (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A1 (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A2_N (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A1 (.DIODE(_00438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B2 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__B1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__B1 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A2 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B1 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A1 (.DIODE(_01150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A2 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B2 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A2 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__A2 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__B1 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A2 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B1 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__B1 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__B2 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A2 (.DIODE(_00241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__B2 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A2 (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08311__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A1 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A2 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B1 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__B (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__B1 (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A2 (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B2 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__B2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__B2 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08518__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__B1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__C (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__B2 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__B (.DIODE(_00241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B (.DIODE(_00241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A2 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B1 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__B2 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__A1 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__A2 (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__B1 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__C (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A2 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__B (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__A2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A2 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__B (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__A2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__B1 (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__B2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A1 (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B2 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08836__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08838__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A2 (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08842__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__A1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__B1 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__B2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__B1 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__A (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09002__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__A1 (.DIODE(_01150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__B (.DIODE(_02179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__B1 (.DIODE(_02179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__B (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__B (.DIODE(_02192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__C (.DIODE(_02193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__B (.DIODE(_02195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__C (.DIODE(_02196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__B (.DIODE(_02198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09069__B (.DIODE(_02200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__B (.DIODE(_02198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__C (.DIODE(_02200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__D (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__B (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__B (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__C_N (.DIODE(_02208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__D_N (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__B (.DIODE(_02210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A1 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__B1 (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__C1 (.DIODE(_02210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B1_N (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A1_N (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__B (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__B (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__A (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__B (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__B (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__A1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__C1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__A0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__S (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__B (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__B (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A1_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A2_N (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__B1 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__A1 (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A2 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__A1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A3 (.DIODE(_00657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__B (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__B (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A3 (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A3 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A4 (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__C1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__S (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__S (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__S (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__B (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__A1 (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__A3 (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A1 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A2 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A1 (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A3 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__B (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__B (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A (.DIODE(_02636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__B (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__S (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__S (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B2 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A1 (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__B1 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__S (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__A (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A2 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__A (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__A (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__D (.DIODE(_02636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__C1 (.DIODE(_02636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__A1 (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__S (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__S (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__A2 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__B1 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__A2 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09728__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09742__A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A1 (.DIODE(_00438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__A2 (.DIODE(_00349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__B2 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A (.DIODE(_02636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A1 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__S (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__A (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09852__A2 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A2 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__B2 (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__S (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A2 (.DIODE(_03123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__A1_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__A2_N (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__B2 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10056__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10056__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A3 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10058__B (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A1 (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__A1 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__S (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A2 (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__B1 (.DIODE(_03263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__A2 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__B (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__A (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__S (.DIODE(_06321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__A2_N (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__A2 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__D (.DIODE(_03393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A2 (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A1 (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B2 (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__A (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A3 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A1 (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A2 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__B1 (.DIODE(_02179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__C (.DIODE(_02179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__C1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A2 (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__S (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__S (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__C1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10535__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A1_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A2_N (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A1 (.DIODE(_00438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__B2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__B1 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__B2 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__C1 (.DIODE(_03766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A1 (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A2 (.DIODE(_00452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A3 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__A (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__B2 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A2 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A1 (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__A2 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A3 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__B (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10876__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A1_N (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A2_N (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__B1 (.DIODE(_04006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A1 (.DIODE(_00349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A2 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__B (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__B1 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A3 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__A1_N (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__A2_N (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__A2 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__B (.DIODE(_04130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__B (.DIODE(_04130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__B2 (.DIODE(_00349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A3 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__B (.DIODE(_04157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B (.DIODE(_04157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__11075__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__11075__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A2 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11097__B1 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A2 (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__11105__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__B1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__B1 (.DIODE(_04224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__B (.DIODE(_04264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__B1 (.DIODE(_02192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__C (.DIODE(_02192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__A (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A1_N (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A2_N (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A1_N (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__A1 (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__B1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__B1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__B2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__B (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__B (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A2 (.DIODE(_04264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A2 (.DIODE(_02192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__B1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A (.DIODE(_02193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A1 (.DIODE(_02193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__B2 (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A1_N (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__B2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A2 (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11334__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11346__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__C (.DIODE(_02195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__B1 (.DIODE(_02195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A2 (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__B2 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A2 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A3 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11418__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__B2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__B (.DIODE(_00432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__A1_N (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__A2_N (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__A (.DIODE(_04559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A2 (.DIODE(_02195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A (.DIODE(_02196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__C1 (.DIODE(_04599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A (.DIODE(_04559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A (.DIODE(_04559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A3 (.DIODE(_04559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__B1 (.DIODE(_02198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__C (.DIODE(_02198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__C1 (.DIODE(_04695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__B1 (.DIODE(_02200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__A3 (.DIODE(_02200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__S (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__A2 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__C1 (.DIODE(_04784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A1 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11697__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__B1 (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__A3 (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__11761__A1 (.DIODE(_04881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A1 (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__A2 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__A (.DIODE(_04935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__B (.DIODE(_04938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__B1 (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__C (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__A (.DIODE(_04935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__A (.DIODE(_04935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A2 (.DIODE(_04938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__B1 (.DIODE(_02208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A3 (.DIODE(_02208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__C1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__C1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__B1 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__B2 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A2_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__A2 (.DIODE(_02208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__C1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(_05154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12001__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__A2 (.DIODE(_02210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__B1 (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A2 (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A3 (.DIODE(_02210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A1 (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__C1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__A (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__B1 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__A2_N (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__B1 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__B2 (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A1 (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__B1 (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__A2 (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__A (.DIODE(_02220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__B2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__B (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__B1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A4 (.DIODE(_05441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__A (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__B1_N (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__C1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__A (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A1 (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__B2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A2 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__A2 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__C1 (.DIODE(_02318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A2 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A2_N (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__B2 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__B1 (.DIODE(_05526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__B1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A2 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__B (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A2 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A1 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__A0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__A (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__S (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__A (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__A (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__A (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__A (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__A (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__A (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__A (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__A (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A (.DIODE(_05132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__A (.DIODE(_05132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__A (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__A (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A (.DIODE(_05284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A (.DIODE(_05284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__S (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__A (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__A (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__A (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__A (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__A (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__S (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__B (.DIODE(_05736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__B (.DIODE(_05736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A2_N (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__B (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__B (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__S (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__B (.DIODE(_05749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__B (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__B (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__B (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__B (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__B (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__B (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__B (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__B (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__B (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__B (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__B (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__B (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__B (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__B (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__B (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__B (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B (.DIODE(_05132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__B (.DIODE(_05132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__B (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__B (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__B (.DIODE(_05284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__B (.DIODE(_05284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__B (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__B (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__B (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__B (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A2 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__B2 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__A2 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__B (.DIODE(_00218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A (.DIODE(_04552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A1 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__A1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__C1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__A1 (.DIODE(_00450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__A1 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A1 (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A1 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A1 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__A1 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__C1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__A1 (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__A (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A1 (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A1 (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A (.DIODE(_00349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A1 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__A1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__A2 (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A2 (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A1 (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__A2 (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__A1 (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A1 (.DIODE(_00146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__A1 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A1 (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A1 (.DIODE(_00432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A1 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A1 (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A1 (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__C1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__A1 (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__A1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13110__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13110__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout11_A (.DIODE(_00454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(_00451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(_00451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(_00454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(_00205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_A (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(_00349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_00173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(_00173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(_00173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(_00349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(_00256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_00285_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(_00285_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap10_A (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap110_A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap119_A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap128_A (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap250_A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap97_A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap99_A (.DIODE(_00300_));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06531_ (.A(net548),
    .Y(_04400_));
 sky130_fd_sc_hd__inv_2 _06532_ (.A(net550),
    .Y(_04411_));
 sky130_fd_sc_hd__inv_2 _06533_ (.A(net602),
    .Y(_04422_));
 sky130_fd_sc_hd__inv_2 _06534_ (.A(net353),
    .Y(_04432_));
 sky130_fd_sc_hd__inv_2 _06535_ (.A(net357),
    .Y(_04443_));
 sky130_fd_sc_hd__inv_2 _06536_ (.A(net346),
    .Y(_04454_));
 sky130_fd_sc_hd__inv_2 _06537_ (.A(net272),
    .Y(_04465_));
 sky130_fd_sc_hd__inv_2 _06538_ (.A(instruction[3]),
    .Y(_04476_));
 sky130_fd_sc_hd__inv_6 _06539_ (.A(instruction[5]),
    .Y(_04487_));
 sky130_fd_sc_hd__inv_2 _06540_ (.A(net302),
    .Y(_04498_));
 sky130_fd_sc_hd__inv_2 _06541_ (.A(instruction[41]),
    .Y(_04509_));
 sky130_fd_sc_hd__inv_2 _06542_ (.A(reg1_val[8]),
    .Y(_04520_));
 sky130_fd_sc_hd__inv_2 _06543_ (.A(reg1_val[16]),
    .Y(_04531_));
 sky130_fd_sc_hd__inv_2 _06544_ (.A(reg1_val[26]),
    .Y(_04541_));
 sky130_fd_sc_hd__inv_6 _06545_ (.A(reg1_val[31]),
    .Y(_04552_));
 sky130_fd_sc_hd__inv_2 _06546_ (.A(net304),
    .Y(_04563_));
 sky130_fd_sc_hd__inv_2 _06547_ (.A(rst),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2_1 _06548_ (.A(instruction[0]),
    .B(pred_val),
    .Y(_04585_));
 sky130_fd_sc_hd__and2_1 _06549_ (.A(pred_val),
    .B(instruction[1]),
    .X(_04596_));
 sky130_fd_sc_hd__o31a_1 _06550_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(pred_val),
    .X(_04607_));
 sky130_fd_sc_hd__and4b_4 _06551_ (.A_N(instruction[1]),
    .B(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04618_));
 sky130_fd_sc_hd__or3b_4 _06552_ (.A(_04596_),
    .B(_04585_),
    .C_N(instruction[2]),
    .X(_04629_));
 sky130_fd_sc_hd__or2_1 _06553_ (.A(instruction[23]),
    .B(_04618_),
    .X(_04639_));
 sky130_fd_sc_hd__o211a_4 _06554_ (.A1(instruction[16]),
    .A2(_04629_),
    .B1(_04639_),
    .C1(net285),
    .X(reg1_idx[5]));
 sky130_fd_sc_hd__or2_1 _06555_ (.A(instruction[20]),
    .B(_04618_),
    .X(_04660_));
 sky130_fd_sc_hd__o211a_4 _06556_ (.A1(instruction[13]),
    .A2(_04629_),
    .B1(_04660_),
    .C1(net285),
    .X(reg1_idx[2]));
 sky130_fd_sc_hd__or2_1 _06557_ (.A(instruction[21]),
    .B(_04618_),
    .X(_04681_));
 sky130_fd_sc_hd__o211a_4 _06558_ (.A1(instruction[14]),
    .A2(_04629_),
    .B1(_04681_),
    .C1(net285),
    .X(reg1_idx[3]));
 sky130_fd_sc_hd__or2_1 _06559_ (.A(instruction[18]),
    .B(_04618_),
    .X(_04702_));
 sky130_fd_sc_hd__o211a_4 _06560_ (.A1(instruction[11]),
    .A2(_04629_),
    .B1(_04702_),
    .C1(net285),
    .X(reg1_idx[0]));
 sky130_fd_sc_hd__or2_1 _06561_ (.A(instruction[19]),
    .B(_04618_),
    .X(_04723_));
 sky130_fd_sc_hd__o211a_4 _06562_ (.A1(instruction[12]),
    .A2(_04629_),
    .B1(_04723_),
    .C1(net285),
    .X(reg1_idx[1]));
 sky130_fd_sc_hd__or2_1 _06563_ (.A(instruction[22]),
    .B(_04618_),
    .X(_04743_));
 sky130_fd_sc_hd__o211a_4 _06564_ (.A1(instruction[15]),
    .A2(_04629_),
    .B1(_04743_),
    .C1(net286),
    .X(reg1_idx[4]));
 sky130_fd_sc_hd__or4bb_4 _06565_ (.A(instruction[0]),
    .B(instruction[1]),
    .C_N(instruction[2]),
    .D_N(pred_val),
    .X(_04764_));
 sky130_fd_sc_hd__nor2_8 _06566_ (.A(instruction[3]),
    .B(_04764_),
    .Y(is_load));
 sky130_fd_sc_hd__nor2_8 _06567_ (.A(_04476_),
    .B(_04764_),
    .Y(is_store));
 sky130_fd_sc_hd__and4bb_1 _06568_ (.A_N(instruction[0]),
    .B_N(instruction[2]),
    .C(instruction[1]),
    .D(pred_val),
    .X(_04795_));
 sky130_fd_sc_hd__or4bb_4 _06569_ (.A(instruction[0]),
    .B(instruction[2]),
    .C_N(instruction[1]),
    .D_N(pred_val),
    .X(_04806_));
 sky130_fd_sc_hd__o311a_4 _06570_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[41]),
    .C1(pred_val),
    .X(_04817_));
 sky130_fd_sc_hd__and4bb_1 _06571_ (.A_N(instruction[1]),
    .B_N(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04827_));
 sky130_fd_sc_hd__or4bb_2 _06572_ (.A(instruction[1]),
    .B(instruction[2]),
    .C_N(instruction[0]),
    .D_N(pred_val),
    .X(_04838_));
 sky130_fd_sc_hd__and2_4 _06573_ (.A(instruction[25]),
    .B(net286),
    .X(_04849_));
 sky130_fd_sc_hd__o211a_1 _06574_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .X(_04860_));
 sky130_fd_sc_hd__o211ai_1 _06575_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .Y(_04871_));
 sky130_fd_sc_hd__a21o_1 _06576_ (.A1(instruction[41]),
    .A2(_04827_),
    .B1(_04860_),
    .X(_04882_));
 sky130_fd_sc_hd__a21oi_1 _06577_ (.A1(instruction[41]),
    .A2(_04827_),
    .B1(_04860_),
    .Y(_04893_));
 sky130_fd_sc_hd__a221o_1 _06578_ (.A1(instruction[24]),
    .A2(_04817_),
    .B1(_04827_),
    .B2(instruction[41]),
    .C1(_04860_),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _06579_ (.A(net284),
    .B(_04904_),
    .Y(_04915_));
 sky130_fd_sc_hd__and2_4 _06580_ (.A(instruction[39]),
    .B(net286),
    .X(_04925_));
 sky130_fd_sc_hd__nor2_1 _06581_ (.A(net264),
    .B(_04925_),
    .Y(_04936_));
 sky130_fd_sc_hd__o2bb2a_4 _06582_ (.A1_N(reg2_val[29]),
    .A2_N(net282),
    .B1(net231),
    .B2(_04936_),
    .X(_04947_));
 sky130_fd_sc_hd__and2b_1 _06583_ (.A_N(_04947_),
    .B(reg1_val[29]),
    .X(_04958_));
 sky130_fd_sc_hd__nand2b_1 _06584_ (.A_N(reg1_val[29]),
    .B(_04947_),
    .Y(_04969_));
 sky130_fd_sc_hd__and2b_1 _06585_ (.A_N(_04958_),
    .B(_04969_),
    .X(_04980_));
 sky130_fd_sc_hd__and2_4 _06586_ (.A(instruction[38]),
    .B(net286),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _06587_ (.A(net264),
    .B(_04991_),
    .Y(_05002_));
 sky130_fd_sc_hd__o2bb2a_4 _06588_ (.A1_N(reg2_val[28]),
    .A2_N(net282),
    .B1(net231),
    .B2(_05002_),
    .X(_05012_));
 sky130_fd_sc_hd__nand2b_1 _06589_ (.A_N(_05012_),
    .B(reg1_val[28]),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2b_1 _06590_ (.A_N(reg1_val[28]),
    .B(_05012_),
    .Y(_05034_));
 sky130_fd_sc_hd__and2_1 _06591_ (.A(_05023_),
    .B(_05034_),
    .X(_05045_));
 sky130_fd_sc_hd__inv_2 _06592_ (.A(_05045_),
    .Y(_05056_));
 sky130_fd_sc_hd__and2_4 _06593_ (.A(instruction[35]),
    .B(net286),
    .X(_05067_));
 sky130_fd_sc_hd__nor2_1 _06594_ (.A(net264),
    .B(_05067_),
    .Y(_05078_));
 sky130_fd_sc_hd__o2bb2a_4 _06595_ (.A1_N(reg2_val[25]),
    .A2_N(net282),
    .B1(net231),
    .B2(_05078_),
    .X(_05089_));
 sky130_fd_sc_hd__nand2b_1 _06596_ (.A_N(_05089_),
    .B(reg1_val[25]),
    .Y(_05099_));
 sky130_fd_sc_hd__and2b_1 _06597_ (.A_N(reg1_val[25]),
    .B(_05089_),
    .X(_05110_));
 sky130_fd_sc_hd__xor2_2 _06598_ (.A(reg1_val[25]),
    .B(_05089_),
    .X(_05121_));
 sky130_fd_sc_hd__and2_4 _06599_ (.A(instruction[34]),
    .B(net286),
    .X(_05132_));
 sky130_fd_sc_hd__nor2_1 _06600_ (.A(net264),
    .B(_05132_),
    .Y(_05143_));
 sky130_fd_sc_hd__o2bb2a_4 _06601_ (.A1_N(reg2_val[24]),
    .A2_N(net282),
    .B1(net231),
    .B2(_05143_),
    .X(_05154_));
 sky130_fd_sc_hd__nand2b_2 _06602_ (.A_N(_05154_),
    .B(reg1_val[24]),
    .Y(_05165_));
 sky130_fd_sc_hd__and2b_1 _06603_ (.A_N(reg1_val[24]),
    .B(_05154_),
    .X(_05176_));
 sky130_fd_sc_hd__xor2_2 _06604_ (.A(reg1_val[24]),
    .B(_05154_),
    .X(_05186_));
 sky130_fd_sc_hd__or4bb_1 _06605_ (.A(_04980_),
    .B(_05045_),
    .C_N(_05121_),
    .D_N(_05186_),
    .X(_05197_));
 sky130_fd_sc_hd__and2_4 _06606_ (.A(instruction[37]),
    .B(net286),
    .X(_05208_));
 sky130_fd_sc_hd__nor2_1 _06607_ (.A(net262),
    .B(_05208_),
    .Y(_05219_));
 sky130_fd_sc_hd__o2bb2a_1 _06608_ (.A1_N(reg2_val[27]),
    .A2_N(net280),
    .B1(net230),
    .B2(_05219_),
    .X(_05230_));
 sky130_fd_sc_hd__a2bb2o_2 _06609_ (.A1_N(_05219_),
    .A2_N(net230),
    .B1(net280),
    .B2(reg2_val[27]),
    .X(_05241_));
 sky130_fd_sc_hd__nor2_1 _06610_ (.A(reg1_val[27]),
    .B(_05241_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_2 _06611_ (.A(reg1_val[27]),
    .B(_05241_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2b_2 _06612_ (.A_N(_05251_),
    .B(_05262_),
    .Y(_05273_));
 sky130_fd_sc_hd__and2_4 _06613_ (.A(instruction[36]),
    .B(net286),
    .X(_05284_));
 sky130_fd_sc_hd__nor2_1 _06614_ (.A(net264),
    .B(_05284_),
    .Y(_05295_));
 sky130_fd_sc_hd__a2bb2o_4 _06615_ (.A1_N(_05295_),
    .A2_N(net231),
    .B1(net282),
    .B2(reg2_val[26]),
    .X(_05306_));
 sky130_fd_sc_hd__nand2_2 _06616_ (.A(reg1_val[26]),
    .B(_05306_),
    .Y(_05317_));
 sky130_fd_sc_hd__inv_2 _06617_ (.A(_05317_),
    .Y(_05327_));
 sky130_fd_sc_hd__or2_1 _06618_ (.A(reg1_val[26]),
    .B(_05306_),
    .X(_05338_));
 sky130_fd_sc_hd__nand2_2 _06619_ (.A(_05317_),
    .B(_05338_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _06620_ (.A(_05273_),
    .B(_05349_),
    .Y(_05360_));
 sky130_fd_sc_hd__and2_1 _06621_ (.A(reg2_val[31]),
    .B(net282),
    .X(_05371_));
 sky130_fd_sc_hd__o21ba_2 _06622_ (.A1(_04509_),
    .A2(net231),
    .B1_N(_05371_),
    .X(_05382_));
 sky130_fd_sc_hd__a31o_4 _06623_ (.A1(instruction[41]),
    .A2(net284),
    .A3(_04904_),
    .B1(_05371_),
    .X(_05392_));
 sky130_fd_sc_hd__xnor2_4 _06624_ (.A(_04552_),
    .B(_05392_),
    .Y(_05403_));
 sky130_fd_sc_hd__and2_4 _06625_ (.A(instruction[40]),
    .B(net286),
    .X(_05414_));
 sky130_fd_sc_hd__nor2_1 _06626_ (.A(net262),
    .B(_05414_),
    .Y(_05425_));
 sky130_fd_sc_hd__o2bb2a_1 _06627_ (.A1_N(reg2_val[30]),
    .A2_N(net280),
    .B1(net230),
    .B2(_05425_),
    .X(_05436_));
 sky130_fd_sc_hd__a2bb2o_2 _06628_ (.A1_N(_05425_),
    .A2_N(net230),
    .B1(net280),
    .B2(reg2_val[30]),
    .X(_05446_));
 sky130_fd_sc_hd__and2_1 _06629_ (.A(reg1_val[30]),
    .B(_05446_),
    .X(_05457_));
 sky130_fd_sc_hd__nor2_1 _06630_ (.A(reg1_val[30]),
    .B(_05446_),
    .Y(_05468_));
 sky130_fd_sc_hd__nor2_2 _06631_ (.A(_05457_),
    .B(_05468_),
    .Y(_05479_));
 sky130_fd_sc_hd__or4_1 _06632_ (.A(_05197_),
    .B(_05360_),
    .C(_05403_),
    .D(_05479_),
    .X(_05490_));
 sky130_fd_sc_hd__and2_4 _06633_ (.A(instruction[33]),
    .B(net286),
    .X(_05500_));
 sky130_fd_sc_hd__nor2_1 _06634_ (.A(net263),
    .B(_05500_),
    .Y(_05511_));
 sky130_fd_sc_hd__o2bb2a_2 _06635_ (.A1_N(reg2_val[23]),
    .A2_N(net281),
    .B1(net230),
    .B2(_05511_),
    .X(_05522_));
 sky130_fd_sc_hd__a2bb2o_1 _06636_ (.A1_N(_05511_),
    .A2_N(net230),
    .B1(net281),
    .B2(reg2_val[23]),
    .X(_05533_));
 sky130_fd_sc_hd__and2_1 _06637_ (.A(reg1_val[23]),
    .B(_05533_),
    .X(_05544_));
 sky130_fd_sc_hd__nor2_1 _06638_ (.A(reg1_val[23]),
    .B(_05533_),
    .Y(_05554_));
 sky130_fd_sc_hd__nor2_1 _06639_ (.A(_05544_),
    .B(_05554_),
    .Y(_05565_));
 sky130_fd_sc_hd__and2_4 _06640_ (.A(instruction[32]),
    .B(net285),
    .X(_05576_));
 sky130_fd_sc_hd__nor2_1 _06641_ (.A(net263),
    .B(_05576_),
    .Y(_05585_));
 sky130_fd_sc_hd__o2bb2a_4 _06642_ (.A1_N(reg2_val[22]),
    .A2_N(net281),
    .B1(net230),
    .B2(_05585_),
    .X(_05595_));
 sky130_fd_sc_hd__a2bb2o_2 _06643_ (.A1_N(_05585_),
    .A2_N(net230),
    .B1(net281),
    .B2(reg2_val[22]),
    .X(_05604_));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(reg1_val[22]),
    .B(_05604_),
    .Y(_05614_));
 sky130_fd_sc_hd__inv_2 _06645_ (.A(_05614_),
    .Y(_05623_));
 sky130_fd_sc_hd__nor2_1 _06646_ (.A(reg1_val[22]),
    .B(_05604_),
    .Y(_05633_));
 sky130_fd_sc_hd__nor2_2 _06647_ (.A(_05623_),
    .B(_05633_),
    .Y(_05643_));
 sky130_fd_sc_hd__and2_4 _06648_ (.A(instruction[30]),
    .B(net285),
    .X(_05652_));
 sky130_fd_sc_hd__nor2_1 _06649_ (.A(net262),
    .B(_05652_),
    .Y(_05662_));
 sky130_fd_sc_hd__o2bb2a_2 _06650_ (.A1_N(reg2_val[20]),
    .A2_N(net281),
    .B1(net230),
    .B2(_05662_),
    .X(_05671_));
 sky130_fd_sc_hd__a2bb2o_2 _06651_ (.A1_N(_05662_),
    .A2_N(net230),
    .B1(net280),
    .B2(reg2_val[20]),
    .X(_05681_));
 sky130_fd_sc_hd__nand2_1 _06652_ (.A(reg1_val[20]),
    .B(_05681_),
    .Y(_05690_));
 sky130_fd_sc_hd__or2_1 _06653_ (.A(reg1_val[20]),
    .B(_05681_),
    .X(_05700_));
 sky130_fd_sc_hd__and2_1 _06654_ (.A(_05690_),
    .B(_05700_),
    .X(_05709_));
 sky130_fd_sc_hd__o311a_4 _06655_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[31]),
    .C1(pred_val),
    .X(_05718_));
 sky130_fd_sc_hd__nor2_1 _06656_ (.A(net264),
    .B(_05718_),
    .Y(_05728_));
 sky130_fd_sc_hd__o2bb2a_2 _06657_ (.A1_N(reg2_val[21]),
    .A2_N(net282),
    .B1(net231),
    .B2(_05728_),
    .X(_05737_));
 sky130_fd_sc_hd__and2b_1 _06658_ (.A_N(_05737_),
    .B(reg1_val[21]),
    .X(_05747_));
 sky130_fd_sc_hd__and2b_1 _06659_ (.A_N(reg1_val[21]),
    .B(_05737_),
    .X(_05755_));
 sky130_fd_sc_hd__nor2_2 _06660_ (.A(_05747_),
    .B(_05755_),
    .Y(_05764_));
 sky130_fd_sc_hd__nor4_1 _06661_ (.A(_05565_),
    .B(_05643_),
    .C(_05709_),
    .D(_05764_),
    .Y(_05773_));
 sky130_fd_sc_hd__and2_4 _06662_ (.A(instruction[29]),
    .B(net285),
    .X(_05782_));
 sky130_fd_sc_hd__nor2_1 _06663_ (.A(net264),
    .B(_05782_),
    .Y(_05791_));
 sky130_fd_sc_hd__o2bb2a_2 _06664_ (.A1_N(reg2_val[19]),
    .A2_N(net282),
    .B1(net230),
    .B2(_05791_),
    .X(_05800_));
 sky130_fd_sc_hd__and2b_1 _06665_ (.A_N(_05800_),
    .B(reg1_val[19]),
    .X(_05810_));
 sky130_fd_sc_hd__inv_2 _06666_ (.A(_05810_),
    .Y(_05819_));
 sky130_fd_sc_hd__and2b_1 _06667_ (.A_N(reg1_val[19]),
    .B(_05800_),
    .X(_05828_));
 sky130_fd_sc_hd__nor2_2 _06668_ (.A(_05810_),
    .B(_05828_),
    .Y(_05836_));
 sky130_fd_sc_hd__and2_4 _06669_ (.A(instruction[28]),
    .B(net285),
    .X(_05845_));
 sky130_fd_sc_hd__nor2_1 _06670_ (.A(net264),
    .B(_05845_),
    .Y(_05854_));
 sky130_fd_sc_hd__o2bb2a_1 _06671_ (.A1_N(reg2_val[18]),
    .A2_N(net282),
    .B1(net230),
    .B2(_05854_),
    .X(_05863_));
 sky130_fd_sc_hd__a2bb2o_2 _06672_ (.A1_N(_05854_),
    .A2_N(net230),
    .B1(net282),
    .B2(reg2_val[18]),
    .X(_05871_));
 sky130_fd_sc_hd__and2_1 _06673_ (.A(reg1_val[18]),
    .B(_05871_),
    .X(_05881_));
 sky130_fd_sc_hd__nand2_1 _06674_ (.A(reg1_val[18]),
    .B(_05871_),
    .Y(_05890_));
 sky130_fd_sc_hd__nor2_1 _06675_ (.A(reg1_val[18]),
    .B(_05871_),
    .Y(_05899_));
 sky130_fd_sc_hd__nor2_2 _06676_ (.A(_05881_),
    .B(_05899_),
    .Y(_05905_));
 sky130_fd_sc_hd__inv_2 _06677_ (.A(_05905_),
    .Y(_05911_));
 sky130_fd_sc_hd__and2_4 _06678_ (.A(instruction[27]),
    .B(net285),
    .X(_05917_));
 sky130_fd_sc_hd__nor2_1 _06679_ (.A(net264),
    .B(_05917_),
    .Y(_05923_));
 sky130_fd_sc_hd__o2bb2a_2 _06680_ (.A1_N(reg2_val[17]),
    .A2_N(_04806_),
    .B1(net230),
    .B2(_05923_),
    .X(_05929_));
 sky130_fd_sc_hd__a2bb2o_2 _06681_ (.A1_N(_05923_),
    .A2_N(net230),
    .B1(_04806_),
    .B2(reg2_val[17]),
    .X(_05935_));
 sky130_fd_sc_hd__nor2_1 _06682_ (.A(reg1_val[17]),
    .B(_05935_),
    .Y(_05943_));
 sky130_fd_sc_hd__or2_1 _06683_ (.A(reg1_val[17]),
    .B(_05935_),
    .X(_05954_));
 sky130_fd_sc_hd__and2_1 _06684_ (.A(reg1_val[17]),
    .B(_05935_),
    .X(_05965_));
 sky130_fd_sc_hd__nor2_1 _06685_ (.A(_05943_),
    .B(_05965_),
    .Y(_05976_));
 sky130_fd_sc_hd__o311a_4 _06686_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[26]),
    .C1(pred_val),
    .X(_05987_));
 sky130_fd_sc_hd__nor2_1 _06687_ (.A(net264),
    .B(_05987_),
    .Y(_05998_));
 sky130_fd_sc_hd__o2bb2a_2 _06688_ (.A1_N(reg2_val[16]),
    .A2_N(net282),
    .B1(net231),
    .B2(_05998_),
    .X(_06009_));
 sky130_fd_sc_hd__a2bb2o_2 _06689_ (.A1_N(_05998_),
    .A2_N(net230),
    .B1(net282),
    .B2(reg2_val[16]),
    .X(_06020_));
 sky130_fd_sc_hd__nor2_1 _06690_ (.A(reg1_val[16]),
    .B(_06020_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(_04531_),
    .B(_06009_),
    .Y(_06042_));
 sky130_fd_sc_hd__nor2_1 _06692_ (.A(_04531_),
    .B(_06009_),
    .Y(_06053_));
 sky130_fd_sc_hd__nor2_2 _06693_ (.A(_06031_),
    .B(_06053_),
    .Y(_06059_));
 sky130_fd_sc_hd__and2_1 _06694_ (.A(reg2_val[15]),
    .B(net281),
    .X(_06065_));
 sky130_fd_sc_hd__a31o_4 _06695_ (.A1(net283),
    .A2(_04817_),
    .A3(net263),
    .B1(_06065_),
    .X(_06071_));
 sky130_fd_sc_hd__nor2_1 _06696_ (.A(reg1_val[15]),
    .B(_06071_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_1 _06697_ (.A(reg1_val[15]),
    .B(_06071_),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2b_2 _06698_ (.A_N(_06077_),
    .B(_06083_),
    .Y(_06089_));
 sky130_fd_sc_hd__and2_1 _06699_ (.A(reg2_val[14]),
    .B(net281),
    .X(_06095_));
 sky130_fd_sc_hd__a31o_4 _06700_ (.A1(net284),
    .A2(net263),
    .A3(_05414_),
    .B1(_06095_),
    .X(_06101_));
 sky130_fd_sc_hd__nor2_1 _06701_ (.A(reg1_val[14]),
    .B(_06101_),
    .Y(_06107_));
 sky130_fd_sc_hd__or2_1 _06702_ (.A(reg1_val[14]),
    .B(_06101_),
    .X(_06113_));
 sky130_fd_sc_hd__and2_1 _06703_ (.A(reg1_val[14]),
    .B(_06101_),
    .X(_06119_));
 sky130_fd_sc_hd__nor2_2 _06704_ (.A(_06107_),
    .B(_06119_),
    .Y(_06125_));
 sky130_fd_sc_hd__inv_2 _06705_ (.A(_06125_),
    .Y(_06132_));
 sky130_fd_sc_hd__and2_1 _06706_ (.A(reg2_val[13]),
    .B(net281),
    .X(_06140_));
 sky130_fd_sc_hd__a31o_4 _06707_ (.A1(net284),
    .A2(net263),
    .A3(_04925_),
    .B1(_06140_),
    .X(_06149_));
 sky130_fd_sc_hd__nor2_1 _06708_ (.A(reg1_val[13]),
    .B(_06149_),
    .Y(_06158_));
 sky130_fd_sc_hd__nand2_1 _06709_ (.A(reg1_val[13]),
    .B(_06149_),
    .Y(_06167_));
 sky130_fd_sc_hd__nand2b_2 _06710_ (.A_N(_06158_),
    .B(_06167_),
    .Y(_06176_));
 sky130_fd_sc_hd__and2_1 _06711_ (.A(reg2_val[12]),
    .B(net281),
    .X(_06185_));
 sky130_fd_sc_hd__a31o_4 _06712_ (.A1(net284),
    .A2(net263),
    .A3(_04991_),
    .B1(_06185_),
    .X(_06194_));
 sky130_fd_sc_hd__nor2_1 _06713_ (.A(reg1_val[12]),
    .B(_06194_),
    .Y(_06203_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(reg1_val[12]),
    .B(_06194_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2b_2 _06715_ (.A_N(_06203_),
    .B(_06212_),
    .Y(_06221_));
 sky130_fd_sc_hd__and2_1 _06716_ (.A(reg2_val[11]),
    .B(net281),
    .X(_06230_));
 sky130_fd_sc_hd__a31o_2 _06717_ (.A1(net283),
    .A2(net263),
    .A3(_05208_),
    .B1(_06230_),
    .X(_06238_));
 sky130_fd_sc_hd__inv_2 _06718_ (.A(_06238_),
    .Y(_06247_));
 sky130_fd_sc_hd__nor2_1 _06719_ (.A(reg1_val[11]),
    .B(_06238_),
    .Y(_06256_));
 sky130_fd_sc_hd__and2_1 _06720_ (.A(reg1_val[11]),
    .B(_06238_),
    .X(_06263_));
 sky130_fd_sc_hd__nor2_1 _06721_ (.A(_06256_),
    .B(_06263_),
    .Y(_06269_));
 sky130_fd_sc_hd__or2_1 _06722_ (.A(_06256_),
    .B(_06263_),
    .X(_06270_));
 sky130_fd_sc_hd__and2_1 _06723_ (.A(reg2_val[10]),
    .B(net281),
    .X(_06271_));
 sky130_fd_sc_hd__a31o_4 _06724_ (.A1(net283),
    .A2(net263),
    .A3(_05284_),
    .B1(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__inv_2 _06725_ (.A(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__or2_1 _06726_ (.A(reg1_val[10]),
    .B(_06272_),
    .X(_06274_));
 sky130_fd_sc_hd__nand2_1 _06727_ (.A(reg1_val[10]),
    .B(_06272_),
    .Y(_06275_));
 sky130_fd_sc_hd__nand2_2 _06728_ (.A(_06274_),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__and2_1 _06729_ (.A(reg2_val[9]),
    .B(net281),
    .X(_06277_));
 sky130_fd_sc_hd__a31o_4 _06730_ (.A1(net283),
    .A2(net263),
    .A3(_05067_),
    .B1(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__inv_2 _06731_ (.A(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_1 _06732_ (.A(reg1_val[9]),
    .B(_06278_),
    .Y(_06280_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(reg1_val[9]),
    .B(_06278_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2b_2 _06734_ (.A_N(_06280_),
    .B(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__and2_1 _06735_ (.A(reg2_val[8]),
    .B(net280),
    .X(_06283_));
 sky130_fd_sc_hd__a31o_4 _06736_ (.A1(net283),
    .A2(net262),
    .A3(_05132_),
    .B1(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__or2_1 _06737_ (.A(reg1_val[8]),
    .B(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__nand2_1 _06738_ (.A(reg1_val[8]),
    .B(_06284_),
    .Y(_06286_));
 sky130_fd_sc_hd__and2_1 _06739_ (.A(_06285_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__and2_1 _06740_ (.A(reg2_val[7]),
    .B(net280),
    .X(_06288_));
 sky130_fd_sc_hd__a31o_4 _06741_ (.A1(net283),
    .A2(net262),
    .A3(_05500_),
    .B1(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__nor2_1 _06742_ (.A(reg1_val[7]),
    .B(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2_1 _06743_ (.A(reg1_val[7]),
    .B(_06289_),
    .Y(_06291_));
 sky130_fd_sc_hd__nand2b_2 _06744_ (.A_N(_06290_),
    .B(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__and2_1 _06745_ (.A(reg2_val[6]),
    .B(net280),
    .X(_06293_));
 sky130_fd_sc_hd__a31o_4 _06746_ (.A1(net283),
    .A2(net262),
    .A3(_05576_),
    .B1(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__or2_1 _06747_ (.A(reg1_val[6]),
    .B(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__and2_1 _06748_ (.A(reg1_val[6]),
    .B(_06294_),
    .X(_06296_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(reg1_val[6]),
    .B(_06294_),
    .Y(_06297_));
 sky130_fd_sc_hd__and2_1 _06750_ (.A(_06295_),
    .B(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__o2111a_4 _06751_ (.A1(_04509_),
    .A2(_04838_),
    .B1(_04871_),
    .C1(_05718_),
    .D1(net284),
    .X(_06299_));
 sky130_fd_sc_hd__or3b_4 _06752_ (.A(net282),
    .B(_04882_),
    .C_N(_05718_),
    .X(_06300_));
 sky130_fd_sc_hd__a21oi_2 _06753_ (.A1(reg2_val[5]),
    .A2(net280),
    .B1(_06299_),
    .Y(_06301_));
 sky130_fd_sc_hd__a21o_2 _06754_ (.A1(reg2_val[5]),
    .A2(net280),
    .B1(_06299_),
    .X(_06302_));
 sky130_fd_sc_hd__nor2_1 _06755_ (.A(reg1_val[5]),
    .B(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__or2_1 _06756_ (.A(reg1_val[5]),
    .B(_06302_),
    .X(_06304_));
 sky130_fd_sc_hd__nand2_1 _06757_ (.A(reg1_val[5]),
    .B(_06302_),
    .Y(_06305_));
 sky130_fd_sc_hd__and2_1 _06758_ (.A(_06304_),
    .B(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__and2_1 _06759_ (.A(reg2_val[4]),
    .B(net280),
    .X(_06307_));
 sky130_fd_sc_hd__a31o_1 _06760_ (.A1(net283),
    .A2(net262),
    .A3(_05652_),
    .B1(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__a31oi_2 _06761_ (.A1(net283),
    .A2(net262),
    .A3(_05652_),
    .B1(_06307_),
    .Y(_06309_));
 sky130_fd_sc_hd__nor2_1 _06762_ (.A(reg1_val[4]),
    .B(net228),
    .Y(_06310_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(reg1_val[4]),
    .B(net228),
    .Y(_06311_));
 sky130_fd_sc_hd__nand2b_2 _06764_ (.A_N(_06310_),
    .B(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__and2_1 _06765_ (.A(reg2_val[3]),
    .B(net280),
    .X(_06313_));
 sky130_fd_sc_hd__a31oi_4 _06766_ (.A1(net283),
    .A2(net262),
    .A3(_05782_),
    .B1(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__a31o_1 _06767_ (.A1(net283),
    .A2(net262),
    .A3(_05782_),
    .B1(_06313_),
    .X(_06315_));
 sky130_fd_sc_hd__nor2_1 _06768_ (.A(reg1_val[3]),
    .B(net223),
    .Y(_06316_));
 sky130_fd_sc_hd__nand2_1 _06769_ (.A(reg1_val[3]),
    .B(net223),
    .Y(_06317_));
 sky130_fd_sc_hd__and2b_1 _06770_ (.A_N(_06316_),
    .B(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__nand2b_1 _06771_ (.A_N(_06316_),
    .B(_06317_),
    .Y(_06319_));
 sky130_fd_sc_hd__and2_1 _06772_ (.A(reg2_val[2]),
    .B(net280),
    .X(_06320_));
 sky130_fd_sc_hd__a31oi_4 _06773_ (.A1(net283),
    .A2(net262),
    .A3(_05845_),
    .B1(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a31o_4 _06774_ (.A1(net283),
    .A2(net262),
    .A3(_05845_),
    .B1(_06320_),
    .X(_06322_));
 sky130_fd_sc_hd__nor2_1 _06775_ (.A(reg1_val[2]),
    .B(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2_1 _06776_ (.A(reg1_val[2]),
    .B(_06322_),
    .Y(_06324_));
 sky130_fd_sc_hd__nand2b_2 _06777_ (.A_N(_06323_),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__and2_1 _06778_ (.A(reg2_val[1]),
    .B(net280),
    .X(_06326_));
 sky130_fd_sc_hd__a31oi_4 _06779_ (.A1(net283),
    .A2(net262),
    .A3(_05917_),
    .B1(_06326_),
    .Y(_06327_));
 sky130_fd_sc_hd__a31o_1 _06780_ (.A1(net283),
    .A2(net262),
    .A3(_05917_),
    .B1(_06326_),
    .X(_06328_));
 sky130_fd_sc_hd__or2_1 _06781_ (.A(net301),
    .B(net219),
    .X(_06329_));
 sky130_fd_sc_hd__xnor2_2 _06782_ (.A(net301),
    .B(net219),
    .Y(_06330_));
 sky130_fd_sc_hd__and2_1 _06783_ (.A(net283),
    .B(_05987_),
    .X(_06331_));
 sky130_fd_sc_hd__a22oi_1 _06784_ (.A1(reg2_val[0]),
    .A2(net280),
    .B1(net262),
    .B2(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__a22o_1 _06785_ (.A1(reg2_val[0]),
    .A2(net280),
    .B1(net262),
    .B2(_06331_),
    .X(_06333_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(net299),
    .B(net213),
    .Y(_06334_));
 sky130_fd_sc_hd__and2_1 _06787_ (.A(net301),
    .B(_06327_),
    .X(_06335_));
 sky130_fd_sc_hd__a21o_1 _06788_ (.A1(_06330_),
    .A2(_06334_),
    .B1(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__and2_1 _06789_ (.A(reg1_val[2]),
    .B(_06321_),
    .X(_06337_));
 sky130_fd_sc_hd__a21oi_1 _06790_ (.A1(_06325_),
    .A2(_06336_),
    .B1(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(reg1_val[3]),
    .B(_06314_),
    .Y(_06339_));
 sky130_fd_sc_hd__o21ai_1 _06792_ (.A1(_06318_),
    .A2(_06338_),
    .B1(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__and2_1 _06793_ (.A(reg1_val[4]),
    .B(net225),
    .X(_06341_));
 sky130_fd_sc_hd__a21oi_1 _06794_ (.A1(_06312_),
    .A2(_06340_),
    .B1(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(reg1_val[5]),
    .B(_06301_),
    .Y(_06343_));
 sky130_fd_sc_hd__o21a_1 _06796_ (.A1(_06306_),
    .A2(_06342_),
    .B1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__nand2b_1 _06797_ (.A_N(_06294_),
    .B(reg1_val[6]),
    .Y(_06345_));
 sky130_fd_sc_hd__o21ai_1 _06798_ (.A1(_06298_),
    .A2(_06344_),
    .B1(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__and2b_1 _06799_ (.A_N(_06289_),
    .B(reg1_val[7]),
    .X(_06347_));
 sky130_fd_sc_hd__a21oi_1 _06800_ (.A1(_06292_),
    .A2(_06346_),
    .B1(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__or2_1 _06801_ (.A(_06287_),
    .B(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__o21ai_1 _06802_ (.A1(_04520_),
    .A2(_06284_),
    .B1(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__and2_1 _06803_ (.A(reg1_val[9]),
    .B(_06279_),
    .X(_06351_));
 sky130_fd_sc_hd__a21o_1 _06804_ (.A1(_06282_),
    .A2(_06350_),
    .B1(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__and2_1 _06805_ (.A(reg1_val[10]),
    .B(_06273_),
    .X(_06353_));
 sky130_fd_sc_hd__a21oi_1 _06806_ (.A1(_06276_),
    .A2(_06352_),
    .B1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(reg1_val[11]),
    .B(_06247_),
    .Y(_06355_));
 sky130_fd_sc_hd__o21ai_1 _06808_ (.A1(_06269_),
    .A2(_06354_),
    .B1(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__and2b_1 _06809_ (.A_N(_06194_),
    .B(reg1_val[12]),
    .X(_06357_));
 sky130_fd_sc_hd__a21o_1 _06810_ (.A1(_06221_),
    .A2(_06356_),
    .B1(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__and2b_1 _06811_ (.A_N(_06149_),
    .B(reg1_val[13]),
    .X(_06359_));
 sky130_fd_sc_hd__a21oi_1 _06812_ (.A1(_06176_),
    .A2(_06358_),
    .B1(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2b_1 _06813_ (.A_N(_06101_),
    .B(reg1_val[14]),
    .Y(_06361_));
 sky130_fd_sc_hd__o21ai_1 _06814_ (.A1(_06125_),
    .A2(_06360_),
    .B1(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__and2b_1 _06815_ (.A_N(_06071_),
    .B(reg1_val[15]),
    .X(_06363_));
 sky130_fd_sc_hd__a21oi_1 _06816_ (.A1(_06089_),
    .A2(_06362_),
    .B1(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__nand2_1 _06817_ (.A(reg1_val[16]),
    .B(_06009_),
    .Y(_06365_));
 sky130_fd_sc_hd__o21a_1 _06818_ (.A1(_06059_),
    .A2(_06364_),
    .B1(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__nand2_1 _06819_ (.A(reg1_val[17]),
    .B(_05929_),
    .Y(_06367_));
 sky130_fd_sc_hd__o21ai_1 _06820_ (.A1(_05976_),
    .A2(_06366_),
    .B1(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__and2_1 _06821_ (.A(reg1_val[18]),
    .B(_05863_),
    .X(_06369_));
 sky130_fd_sc_hd__a21oi_2 _06822_ (.A1(_05911_),
    .A2(_06368_),
    .B1(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nand2_1 _06823_ (.A(reg1_val[19]),
    .B(_05800_),
    .Y(_06371_));
 sky130_fd_sc_hd__o21a_1 _06824_ (.A1(_05836_),
    .A2(_06370_),
    .B1(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__o21ai_1 _06825_ (.A1(_05836_),
    .A2(_06370_),
    .B1(_06371_),
    .Y(_06373_));
 sky130_fd_sc_hd__nand2_1 _06826_ (.A(reg1_val[21]),
    .B(_05737_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_1 _06827_ (.A(reg1_val[20]),
    .B(_05671_),
    .Y(_06375_));
 sky130_fd_sc_hd__o21a_1 _06828_ (.A1(_05764_),
    .A2(_06375_),
    .B1(_06374_),
    .X(_06376_));
 sky130_fd_sc_hd__or2_1 _06829_ (.A(_05643_),
    .B(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__nand2_1 _06830_ (.A(reg1_val[22]),
    .B(_05595_),
    .Y(_06378_));
 sky130_fd_sc_hd__a21oi_1 _06831_ (.A1(_06377_),
    .A2(_06378_),
    .B1(_05565_),
    .Y(_06379_));
 sky130_fd_sc_hd__a221o_1 _06832_ (.A1(reg1_val[23]),
    .A2(_05522_),
    .B1(_05773_),
    .B2(_06373_),
    .C1(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__nand2b_1 _06833_ (.A_N(_05490_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(reg1_val[30]),
    .B(_05436_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(reg1_val[29]),
    .B(_04947_),
    .Y(_06383_));
 sky130_fd_sc_hd__and2_1 _06836_ (.A(reg1_val[28]),
    .B(_05012_),
    .X(_06384_));
 sky130_fd_sc_hd__nand2_1 _06837_ (.A(reg1_val[27]),
    .B(_05230_),
    .Y(_06385_));
 sky130_fd_sc_hd__nor2_1 _06838_ (.A(_04541_),
    .B(_05306_),
    .Y(_06386_));
 sky130_fd_sc_hd__and2_1 _06839_ (.A(reg1_val[25]),
    .B(_05089_),
    .X(_06387_));
 sky130_fd_sc_hd__and2_1 _06840_ (.A(reg1_val[24]),
    .B(_05154_),
    .X(_06388_));
 sky130_fd_sc_hd__a21o_1 _06841_ (.A1(_05121_),
    .A2(_06388_),
    .B1(_06387_),
    .X(_06389_));
 sky130_fd_sc_hd__a21o_1 _06842_ (.A1(_05349_),
    .A2(_06389_),
    .B1(_06386_),
    .X(_06390_));
 sky130_fd_sc_hd__nand2_1 _06843_ (.A(_05273_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__a21oi_1 _06844_ (.A1(_06385_),
    .A2(_06391_),
    .B1(_05045_),
    .Y(_06392_));
 sky130_fd_sc_hd__nor2_1 _06845_ (.A(_06384_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__o21a_1 _06846_ (.A1(_04980_),
    .A2(_06393_),
    .B1(_06383_),
    .X(_06394_));
 sky130_fd_sc_hd__o21a_1 _06847_ (.A1(_05479_),
    .A2(_06394_),
    .B1(_06382_),
    .X(_06395_));
 sky130_fd_sc_hd__a21oi_1 _06848_ (.A1(reg1_val[31]),
    .A2(_05382_),
    .B1(net305),
    .Y(_06396_));
 sky130_fd_sc_hd__o211a_1 _06849_ (.A1(_05403_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06381_),
    .X(_06397_));
 sky130_fd_sc_hd__a21o_1 _06850_ (.A1(_05186_),
    .A2(_06380_),
    .B1(_06388_),
    .X(_06398_));
 sky130_fd_sc_hd__a21o_1 _06851_ (.A1(_05121_),
    .A2(_06398_),
    .B1(_06387_),
    .X(_06399_));
 sky130_fd_sc_hd__a21o_1 _06852_ (.A1(_05349_),
    .A2(_06399_),
    .B1(_06386_),
    .X(_06400_));
 sky130_fd_sc_hd__a21bo_1 _06853_ (.A1(_05273_),
    .A2(_06400_),
    .B1_N(_06385_),
    .X(_06401_));
 sky130_fd_sc_hd__a21oi_1 _06854_ (.A1(_05056_),
    .A2(_06401_),
    .B1(_06384_),
    .Y(_06402_));
 sky130_fd_sc_hd__o21a_1 _06855_ (.A1(_04980_),
    .A2(_06402_),
    .B1(_06383_),
    .X(_06403_));
 sky130_fd_sc_hd__nor2_1 _06856_ (.A(_05479_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__o21a_1 _06857_ (.A1(_05479_),
    .A2(_06403_),
    .B1(_06382_),
    .X(_06405_));
 sky130_fd_sc_hd__or3b_1 _06858_ (.A(_06404_),
    .B(_05403_),
    .C_N(_06382_),
    .X(_06406_));
 sky130_fd_sc_hd__o21ai_1 _06859_ (.A1(_04552_),
    .A2(_05392_),
    .B1(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__a21o_1 _06860_ (.A1(net305),
    .A2(_06407_),
    .B1(_06397_),
    .X(_06408_));
 sky130_fd_sc_hd__or2_4 _06861_ (.A(instruction[4]),
    .B(instruction[3]),
    .X(_06409_));
 sky130_fd_sc_hd__inv_2 _06862_ (.A(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__nand2_2 _06863_ (.A(net302),
    .B(net213),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(net299),
    .B(net216),
    .Y(_06412_));
 sky130_fd_sc_hd__nor4_1 _06865_ (.A(_05836_),
    .B(_05905_),
    .C(_05976_),
    .D(_06059_),
    .Y(_06413_));
 sky130_fd_sc_hd__and4_1 _06866_ (.A(_06270_),
    .B(_06276_),
    .C(_06282_),
    .D(_06292_),
    .X(_06414_));
 sky130_fd_sc_hd__and4_1 _06867_ (.A(_06089_),
    .B(_06132_),
    .C(_06176_),
    .D(_06221_),
    .X(_06415_));
 sky130_fd_sc_hd__and4bb_1 _06868_ (.A_N(_06298_),
    .B_N(_06306_),
    .C(_06312_),
    .D(_06319_),
    .X(_06416_));
 sky130_fd_sc_hd__a21oi_1 _06869_ (.A1(_06411_),
    .A2(_06412_),
    .B1(_06287_),
    .Y(_06417_));
 sky130_fd_sc_hd__and4_1 _06870_ (.A(_06325_),
    .B(_06330_),
    .C(_06416_),
    .D(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__and3_1 _06871_ (.A(_06414_),
    .B(_06415_),
    .C(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__and4b_1 _06872_ (.A_N(_05490_),
    .B(_05773_),
    .C(_06413_),
    .D(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__nand2_1 _06873_ (.A(net306),
    .B(_05403_),
    .Y(_06421_));
 sky130_fd_sc_hd__o211a_1 _06874_ (.A1(net305),
    .A2(_06420_),
    .B1(_06421_),
    .C1(_06410_),
    .X(_06422_));
 sky130_fd_sc_hd__nand2_2 _06875_ (.A(instruction[4]),
    .B(instruction[3]),
    .Y(_06423_));
 sky130_fd_sc_hd__inv_2 _06876_ (.A(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__or2_2 _06877_ (.A(instruction[4]),
    .B(_04476_),
    .X(_06425_));
 sky130_fd_sc_hd__a221o_2 _06878_ (.A1(instruction[3]),
    .A2(_06408_),
    .B1(_06420_),
    .B2(_06424_),
    .C1(_06422_),
    .X(_06426_));
 sky130_fd_sc_hd__xnor2_4 _06879_ (.A(_04487_),
    .B(_06426_),
    .Y(dest_pred_val));
 sky130_fd_sc_hd__and3_4 _06880_ (.A(instruction[2]),
    .B(_04585_),
    .C(_04596_),
    .X(_06427_));
 sky130_fd_sc_hd__nand3_1 _06881_ (.A(instruction[2]),
    .B(_04585_),
    .C(_04596_),
    .Y(_06428_));
 sky130_fd_sc_hd__a21o_4 _06882_ (.A1(_04618_),
    .A2(dest_pred_val),
    .B1(net259),
    .X(take_branch));
 sky130_fd_sc_hd__and3_1 _06883_ (.A(reg1_idx[0]),
    .B(reg1_idx[1]),
    .C(reg1_idx[4]),
    .X(_06429_));
 sky130_fd_sc_hd__and2_1 _06884_ (.A(reg1_idx[5]),
    .B(_06427_),
    .X(_06430_));
 sky130_fd_sc_hd__and4_4 _06885_ (.A(reg1_idx[2]),
    .B(reg1_idx[3]),
    .C(_06429_),
    .D(_06430_),
    .X(int_return));
 sky130_fd_sc_hd__nand2_8 _06886_ (.A(net305),
    .B(_04487_),
    .Y(_06431_));
 sky130_fd_sc_hd__nand2_2 _06887_ (.A(net305),
    .B(instruction[5]),
    .Y(_06432_));
 sky130_fd_sc_hd__a21oi_1 _06888_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(instruction[4]),
    .Y(_06433_));
 sky130_fd_sc_hd__a221oi_2 _06889_ (.A1(net282),
    .A2(_04838_),
    .B1(_06431_),
    .B2(instruction[4]),
    .C1(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__a221o_1 _06890_ (.A1(net282),
    .A2(_04838_),
    .B1(_06431_),
    .B2(instruction[4]),
    .C1(_06433_),
    .X(_06435_));
 sky130_fd_sc_hd__nor2_1 _06891_ (.A(net271),
    .B(_06434_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _06892_ (.A(net266),
    .B(_06435_),
    .Y(_06437_));
 sky130_fd_sc_hd__nor2_8 _06893_ (.A(div_complete),
    .B(net196),
    .Y(busy));
 sky130_fd_sc_hd__and4b_4 _06894_ (.A_N(instruction[2]),
    .B(instruction[1]),
    .C(pred_val),
    .D(instruction[0]),
    .X(_06438_));
 sky130_fd_sc_hd__and2_4 _06895_ (.A(instruction[11]),
    .B(_06438_),
    .X(dest_pred[0]));
 sky130_fd_sc_hd__and2_4 _06896_ (.A(instruction[12]),
    .B(_06438_),
    .X(dest_pred[1]));
 sky130_fd_sc_hd__and2_4 _06897_ (.A(instruction[13]),
    .B(_06438_),
    .X(dest_pred[2]));
 sky130_fd_sc_hd__or3_2 _06898_ (.A(net284),
    .B(_04827_),
    .C(_06427_),
    .X(_06439_));
 sky130_fd_sc_hd__and2_4 _06899_ (.A(instruction[11]),
    .B(_06439_),
    .X(dest_idx[0]));
 sky130_fd_sc_hd__and2_4 _06900_ (.A(instruction[12]),
    .B(_06439_),
    .X(dest_idx[1]));
 sky130_fd_sc_hd__and2_4 _06901_ (.A(instruction[13]),
    .B(_06439_),
    .X(dest_idx[2]));
 sky130_fd_sc_hd__and2_4 _06902_ (.A(instruction[14]),
    .B(_06439_),
    .X(dest_idx[3]));
 sky130_fd_sc_hd__and2_4 _06903_ (.A(instruction[15]),
    .B(_06439_),
    .X(dest_idx[4]));
 sky130_fd_sc_hd__and2_4 _06904_ (.A(instruction[16]),
    .B(_06439_),
    .X(dest_idx[5]));
 sky130_fd_sc_hd__or2_1 _06905_ (.A(instruction[25]),
    .B(_04618_),
    .X(_06440_));
 sky130_fd_sc_hd__o211a_4 _06906_ (.A1(instruction[18]),
    .A2(_04629_),
    .B1(_06440_),
    .C1(net285),
    .X(reg2_idx[0]));
 sky130_fd_sc_hd__or2_1 _06907_ (.A(instruction[26]),
    .B(_04618_),
    .X(_06441_));
 sky130_fd_sc_hd__o211a_4 _06908_ (.A1(instruction[19]),
    .A2(_04629_),
    .B1(_06441_),
    .C1(net285),
    .X(reg2_idx[1]));
 sky130_fd_sc_hd__or2_1 _06909_ (.A(instruction[27]),
    .B(_04618_),
    .X(_06442_));
 sky130_fd_sc_hd__o211a_4 _06910_ (.A1(instruction[20]),
    .A2(_04629_),
    .B1(_06442_),
    .C1(net285),
    .X(reg2_idx[2]));
 sky130_fd_sc_hd__or2_1 _06911_ (.A(instruction[28]),
    .B(_04618_),
    .X(_06443_));
 sky130_fd_sc_hd__o211a_4 _06912_ (.A1(instruction[21]),
    .A2(_04629_),
    .B1(_06443_),
    .C1(net285),
    .X(reg2_idx[3]));
 sky130_fd_sc_hd__or2_1 _06913_ (.A(instruction[29]),
    .B(_04618_),
    .X(_06444_));
 sky130_fd_sc_hd__o211a_4 _06914_ (.A1(instruction[22]),
    .A2(_04629_),
    .B1(_06444_),
    .C1(net285),
    .X(reg2_idx[4]));
 sky130_fd_sc_hd__or2_1 _06915_ (.A(instruction[30]),
    .B(_04618_),
    .X(_06445_));
 sky130_fd_sc_hd__o211a_4 _06916_ (.A1(instruction[23]),
    .A2(_04629_),
    .B1(_06445_),
    .C1(net285),
    .X(reg2_idx[5]));
 sky130_fd_sc_hd__nor3_2 _06917_ (.A(net306),
    .B(instruction[5]),
    .C(_06425_),
    .Y(_06446_));
 sky130_fd_sc_hd__or3_2 _06918_ (.A(net306),
    .B(instruction[5]),
    .C(_06425_),
    .X(_06447_));
 sky130_fd_sc_hd__and4b_1 _06919_ (.A_N(net306),
    .B(instruction[4]),
    .C(_04476_),
    .D(_04487_),
    .X(_06448_));
 sky130_fd_sc_hd__or4b_4 _06920_ (.A(instruction[3]),
    .B(instruction[6]),
    .C(instruction[5]),
    .D_N(instruction[4]),
    .X(_06449_));
 sky130_fd_sc_hd__a31o_1 _06921_ (.A1(instruction[17]),
    .A2(net209),
    .A3(_06449_),
    .B1(net282),
    .X(_06450_));
 sky130_fd_sc_hd__o221a_1 _06922_ (.A1(instruction[3]),
    .A2(_04764_),
    .B1(_04838_),
    .B2(instruction[40]),
    .C1(_06431_),
    .X(_06451_));
 sky130_fd_sc_hd__and3_1 _06923_ (.A(_04882_),
    .B(_06450_),
    .C(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__a31o_2 _06924_ (.A1(instruction[24]),
    .A2(net304),
    .A3(is_load),
    .B1(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__nand2_8 _06925_ (.A(net257),
    .B(_06453_),
    .Y(dest_mask[0]));
 sky130_fd_sc_hd__a32o_2 _06926_ (.A1(net264),
    .A2(_06450_),
    .A3(_06451_),
    .B1(is_load),
    .B2(net304),
    .X(_06454_));
 sky130_fd_sc_hd__nand2_8 _06927_ (.A(net257),
    .B(_06454_),
    .Y(dest_mask[1]));
 sky130_fd_sc_hd__and4b_4 _06928_ (.A_N(net306),
    .B(instruction[5]),
    .C(net303),
    .D(_06410_),
    .X(_06455_));
 sky130_fd_sc_hd__or4_2 _06929_ (.A(net305),
    .B(_04487_),
    .C(net298),
    .D(_06409_),
    .X(_06456_));
 sky130_fd_sc_hd__o21ai_4 _06930_ (.A1(_06410_),
    .A2(_06432_),
    .B1(net251),
    .Y(_06457_));
 sky130_fd_sc_hd__and2_1 _06931_ (.A(reg1_val[31]),
    .B(net303),
    .X(_06458_));
 sky130_fd_sc_hd__or4_2 _06932_ (.A(net302),
    .B(net301),
    .C(reg1_val[2]),
    .D(reg1_val[3]),
    .X(_06459_));
 sky130_fd_sc_hd__or4_2 _06933_ (.A(reg1_val[4]),
    .B(reg1_val[5]),
    .C(reg1_val[6]),
    .D(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__or4_2 _06934_ (.A(reg1_val[7]),
    .B(reg1_val[8]),
    .C(reg1_val[9]),
    .D(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__or4_4 _06935_ (.A(reg1_val[10]),
    .B(reg1_val[11]),
    .C(reg1_val[12]),
    .D(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__or4_4 _06936_ (.A(reg1_val[13]),
    .B(reg1_val[14]),
    .C(reg1_val[15]),
    .D(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__or3_1 _06937_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .C(reg1_val[22]),
    .X(_06464_));
 sky130_fd_sc_hd__or2_2 _06938_ (.A(reg1_val[16]),
    .B(reg1_val[17]),
    .X(_06465_));
 sky130_fd_sc_hd__or3_4 _06939_ (.A(reg1_val[18]),
    .B(reg1_val[19]),
    .C(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__or3_4 _06940_ (.A(reg1_val[23]),
    .B(_06464_),
    .C(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__or2_2 _06941_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .X(_06468_));
 sky130_fd_sc_hd__o31a_2 _06942_ (.A1(_06463_),
    .A2(_06467_),
    .A3(_06468_),
    .B1(net274),
    .X(_06469_));
 sky130_fd_sc_hd__o41a_4 _06943_ (.A1(reg1_val[26]),
    .A2(_06463_),
    .A3(_06467_),
    .A4(_06468_),
    .B1(net274),
    .X(_06470_));
 sky130_fd_sc_hd__xor2_2 _06944_ (.A(reg1_val[27]),
    .B(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__xnor2_4 _06945_ (.A(reg1_val[27]),
    .B(_06470_),
    .Y(_06472_));
 sky130_fd_sc_hd__and2_1 _06946_ (.A(net304),
    .B(_05392_),
    .X(_06473_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(net304),
    .B(_05392_),
    .Y(_06474_));
 sky130_fd_sc_hd__and4_1 _06948_ (.A(_06314_),
    .B(_06321_),
    .C(_06327_),
    .D(net214),
    .X(_06475_));
 sky130_fd_sc_hd__or4_4 _06949_ (.A(net223),
    .B(_06322_),
    .C(net219),
    .D(net213),
    .X(_06476_));
 sky130_fd_sc_hd__a21o_1 _06950_ (.A1(net190),
    .A2(_06476_),
    .B1(net228),
    .X(_06477_));
 sky130_fd_sc_hd__or3_2 _06951_ (.A(net225),
    .B(net189),
    .C(_06475_),
    .X(_06478_));
 sky130_fd_sc_hd__nand2_2 _06952_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__o21ai_2 _06953_ (.A1(_06463_),
    .A2(_06467_),
    .B1(net274),
    .Y(_06480_));
 sky130_fd_sc_hd__o31a_2 _06954_ (.A1(reg1_val[24]),
    .A2(_06463_),
    .A3(_06467_),
    .B1(net274),
    .X(_06481_));
 sky130_fd_sc_hd__xor2_4 _06955_ (.A(reg1_val[25]),
    .B(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__xnor2_4 _06956_ (.A(_04541_),
    .B(_06469_),
    .Y(_06483_));
 sky130_fd_sc_hd__and2_1 _06957_ (.A(net117),
    .B(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__nor2_1 _06958_ (.A(net117),
    .B(_06483_),
    .Y(_06485_));
 sky130_fd_sc_hd__nor2_1 _06959_ (.A(_06484_),
    .B(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__or2_1 _06960_ (.A(_06484_),
    .B(_06485_),
    .X(_06487_));
 sky130_fd_sc_hd__o211a_1 _06961_ (.A1(net219),
    .A2(net213),
    .B1(net304),
    .C1(_05392_),
    .X(_06488_));
 sky130_fd_sc_hd__o311a_2 _06962_ (.A1(_06322_),
    .A2(net219),
    .A3(net213),
    .B1(_05392_),
    .C1(net303),
    .X(_06489_));
 sky130_fd_sc_hd__xnor2_2 _06963_ (.A(net223),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__xnor2_4 _06964_ (.A(_06314_),
    .B(_06489_),
    .Y(_06491_));
 sky130_fd_sc_hd__and3_1 _06965_ (.A(_06472_),
    .B(net117),
    .C(_06483_),
    .X(_06492_));
 sky130_fd_sc_hd__a21oi_1 _06966_ (.A1(net120),
    .A2(_06485_),
    .B1(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__o22a_1 _06967_ (.A1(net147),
    .A2(net38),
    .B1(net174),
    .B2(net36),
    .X(_06494_));
 sky130_fd_sc_hd__xnor2_1 _06968_ (.A(net121),
    .B(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__o21ai_2 _06969_ (.A1(_06463_),
    .A2(_06466_),
    .B1(net275),
    .Y(_06496_));
 sky130_fd_sc_hd__o31a_2 _06970_ (.A1(_06463_),
    .A2(_06464_),
    .A3(_06466_),
    .B1(net274),
    .X(_06497_));
 sky130_fd_sc_hd__xor2_4 _06971_ (.A(reg1_val[23]),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__or4_4 _06972_ (.A(_06289_),
    .B(_06294_),
    .C(_06302_),
    .D(net228),
    .X(_06499_));
 sky130_fd_sc_hd__o21ai_4 _06973_ (.A1(_06476_),
    .A2(_06499_),
    .B1(net190),
    .Y(_06500_));
 sky130_fd_sc_hd__xor2_1 _06974_ (.A(_06284_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__xnor2_4 _06975_ (.A(_06284_),
    .B(_06500_),
    .Y(_06502_));
 sky130_fd_sc_hd__o31a_4 _06976_ (.A1(reg1_val[20]),
    .A2(_06463_),
    .A3(_06466_),
    .B1(net275),
    .X(_06503_));
 sky130_fd_sc_hd__xor2_4 _06977_ (.A(reg1_val[21]),
    .B(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__xnor2_4 _06978_ (.A(reg1_val[21]),
    .B(_06503_),
    .Y(_06505_));
 sky130_fd_sc_hd__o41a_2 _06979_ (.A1(reg1_val[20]),
    .A2(reg1_val[21]),
    .A3(_06463_),
    .A4(_06466_),
    .B1(net274),
    .X(_06506_));
 sky130_fd_sc_hd__xor2_4 _06980_ (.A(reg1_val[22]),
    .B(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__xnor2_2 _06981_ (.A(_06505_),
    .B(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__xnor2_2 _06982_ (.A(net112),
    .B(_06507_),
    .Y(_06509_));
 sky130_fd_sc_hd__a31o_2 _06983_ (.A1(_06301_),
    .A2(net225),
    .A3(_06475_),
    .B1(net189),
    .X(_06510_));
 sky130_fd_sc_hd__o41ai_4 _06984_ (.A1(_06294_),
    .A2(_06302_),
    .A3(net228),
    .A4(_06476_),
    .B1(net190),
    .Y(_06511_));
 sky130_fd_sc_hd__xor2_1 _06985_ (.A(_06289_),
    .B(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__xnor2_4 _06986_ (.A(_06289_),
    .B(_06511_),
    .Y(_06513_));
 sky130_fd_sc_hd__or3b_4 _06987_ (.A(net111),
    .B(_06507_),
    .C_N(net114),
    .X(_06514_));
 sky130_fd_sc_hd__or3b_4 _06988_ (.A(net114),
    .B(net110),
    .C_N(_06507_),
    .X(_06515_));
 sky130_fd_sc_hd__and2_1 _06989_ (.A(_06514_),
    .B(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__o22a_1 _06990_ (.A1(net145),
    .A2(net80),
    .B1(net143),
    .B2(net33),
    .X(_06517_));
 sky130_fd_sc_hd__xnor2_1 _06991_ (.A(net114),
    .B(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__and2_1 _06992_ (.A(_06495_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__nor2_1 _06993_ (.A(_06495_),
    .B(_06518_),
    .Y(_06520_));
 sky130_fd_sc_hd__or2_1 _06994_ (.A(_06519_),
    .B(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__xnor2_4 _06995_ (.A(_06294_),
    .B(_06510_),
    .Y(_06522_));
 sky130_fd_sc_hd__xor2_2 _06996_ (.A(_06294_),
    .B(_06510_),
    .X(_06523_));
 sky130_fd_sc_hd__xnor2_4 _06997_ (.A(reg1_val[24]),
    .B(_06480_),
    .Y(_06524_));
 sky130_fd_sc_hd__and2_1 _06998_ (.A(_06498_),
    .B(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__nor2_1 _06999_ (.A(_06498_),
    .B(_06524_),
    .Y(_06526_));
 sky130_fd_sc_hd__or2_4 _07000_ (.A(_06525_),
    .B(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__and3_1 _07001_ (.A(net303),
    .B(_05392_),
    .C(net228),
    .X(_06528_));
 sky130_fd_sc_hd__a211o_1 _07002_ (.A1(_06309_),
    .A2(_06475_),
    .B1(net189),
    .C1(_06302_),
    .X(_06529_));
 sky130_fd_sc_hd__a211o_1 _07003_ (.A1(net190),
    .A2(_06476_),
    .B1(_06528_),
    .C1(_06301_),
    .X(_06530_));
 sky130_fd_sc_hd__and2_2 _07004_ (.A(_06529_),
    .B(_06530_),
    .X(_00136_));
 sky130_fd_sc_hd__nand3b_1 _07005_ (.A_N(net116),
    .B(net113),
    .C(_06524_),
    .Y(_00137_));
 sky130_fd_sc_hd__a21boi_4 _07006_ (.A1(net116),
    .A2(_06526_),
    .B1_N(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__o22a_1 _07007_ (.A1(net141),
    .A2(net31),
    .B1(net139),
    .B2(net30),
    .X(_00139_));
 sky130_fd_sc_hd__xor2_1 _07008_ (.A(net118),
    .B(_00139_),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _07009_ (.A(_06521_),
    .B(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__and2_1 _07010_ (.A(_06521_),
    .B(_00140_),
    .X(_00142_));
 sky130_fd_sc_hd__nor2_1 _07011_ (.A(_00141_),
    .B(_00142_),
    .Y(_00143_));
 sky130_fd_sc_hd__o21a_1 _07012_ (.A1(reg1_val[10]),
    .A2(_06461_),
    .B1(net275),
    .X(_00144_));
 sky130_fd_sc_hd__xnor2_4 _07013_ (.A(reg1_val[11]),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_4 _07014_ (.A(net173),
    .Y(_00146_));
 sky130_fd_sc_hd__or2_1 _07015_ (.A(_06278_),
    .B(_06284_),
    .X(_00147_));
 sky130_fd_sc_hd__nor3_1 _07016_ (.A(_06476_),
    .B(_06499_),
    .C(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__or3_1 _07017_ (.A(_06476_),
    .B(_06499_),
    .C(_00147_),
    .X(_00149_));
 sky130_fd_sc_hd__or2_1 _07018_ (.A(_06238_),
    .B(_06272_),
    .X(_00150_));
 sky130_fd_sc_hd__or4_1 _07019_ (.A(_06071_),
    .B(_06101_),
    .C(_06149_),
    .D(_06194_),
    .X(_00151_));
 sky130_fd_sc_hd__nor2_1 _07020_ (.A(_00150_),
    .B(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__or2_1 _07021_ (.A(_00150_),
    .B(_00151_),
    .X(_00153_));
 sky130_fd_sc_hd__o41a_4 _07022_ (.A1(_05935_),
    .A2(_06020_),
    .A3(_00149_),
    .A4(_00153_),
    .B1(net190),
    .X(_00154_));
 sky130_fd_sc_hd__xnor2_4 _07023_ (.A(_05871_),
    .B(_00154_),
    .Y(_00155_));
 sky130_fd_sc_hd__o21a_1 _07024_ (.A1(reg1_val[7]),
    .A2(_06460_),
    .B1(net275),
    .X(_00156_));
 sky130_fd_sc_hd__o31a_1 _07025_ (.A1(reg1_val[7]),
    .A2(reg1_val[8]),
    .A3(_06460_),
    .B1(net275),
    .X(_00157_));
 sky130_fd_sc_hd__xnor2_2 _07026_ (.A(reg1_val[9]),
    .B(_00157_),
    .Y(_00158_));
 sky130_fd_sc_hd__nand2_1 _07027_ (.A(net275),
    .B(_06461_),
    .Y(_00159_));
 sky130_fd_sc_hd__xor2_2 _07028_ (.A(reg1_val[10]),
    .B(_00159_),
    .X(_00160_));
 sky130_fd_sc_hd__nand2_1 _07029_ (.A(net187),
    .B(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__or2_1 _07030_ (.A(net187),
    .B(_00160_),
    .X(_00162_));
 sky130_fd_sc_hd__nand2_2 _07031_ (.A(_00161_),
    .B(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__a21o_2 _07032_ (.A1(_00148_),
    .A2(_00152_),
    .B1(net189),
    .X(_00164_));
 sky130_fd_sc_hd__a31o_1 _07033_ (.A1(_06009_),
    .A2(_00148_),
    .A3(_00152_),
    .B1(net189),
    .X(_00165_));
 sky130_fd_sc_hd__xnor2_4 _07034_ (.A(_05929_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__mux2_2 _07035_ (.A0(_00161_),
    .A1(_00162_),
    .S(net172),
    .X(_00167_));
 sky130_fd_sc_hd__o22a_1 _07036_ (.A1(_00155_),
    .A2(net107),
    .B1(_00166_),
    .B2(net103),
    .X(_00168_));
 sky130_fd_sc_hd__xnor2_1 _07037_ (.A(net173),
    .B(_00168_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_2 _07038_ (.A(net275),
    .B(_06460_),
    .Y(_00170_));
 sky130_fd_sc_hd__xor2_4 _07039_ (.A(reg1_val[7]),
    .B(_00170_),
    .X(_00171_));
 sky130_fd_sc_hd__o21a_1 _07040_ (.A1(reg1_val[4]),
    .A2(_06459_),
    .B1(net275),
    .X(_00172_));
 sky130_fd_sc_hd__xnor2_4 _07041_ (.A(reg1_val[5]),
    .B(_00172_),
    .Y(_00173_));
 sky130_fd_sc_hd__o31a_2 _07042_ (.A1(reg1_val[4]),
    .A2(reg1_val[5]),
    .A3(_06459_),
    .B1(net275),
    .X(_00174_));
 sky130_fd_sc_hd__xnor2_4 _07043_ (.A(reg1_val[6]),
    .B(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__and2_1 _07044_ (.A(net206),
    .B(_00175_),
    .X(_00176_));
 sky130_fd_sc_hd__nand2_1 _07045_ (.A(net206),
    .B(_00175_),
    .Y(_00177_));
 sky130_fd_sc_hd__nor2_1 _07046_ (.A(net206),
    .B(_00175_),
    .Y(_00178_));
 sky130_fd_sc_hd__or2_2 _07047_ (.A(_00176_),
    .B(_00178_),
    .X(_00179_));
 sky130_fd_sc_hd__inv_2 _07048_ (.A(net170),
    .Y(_00180_));
 sky130_fd_sc_hd__and4_1 _07049_ (.A(_05800_),
    .B(_05863_),
    .C(_05929_),
    .D(_06009_),
    .X(_00181_));
 sky130_fd_sc_hd__and3_2 _07050_ (.A(_00148_),
    .B(_00152_),
    .C(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__or3b_2 _07051_ (.A(_00149_),
    .B(_00153_),
    .C_N(_00181_),
    .X(_00183_));
 sky130_fd_sc_hd__and2_1 _07052_ (.A(_05671_),
    .B(_05737_),
    .X(_00184_));
 sky130_fd_sc_hd__a21o_2 _07053_ (.A1(_00182_),
    .A2(_00184_),
    .B1(net189),
    .X(_00185_));
 sky130_fd_sc_hd__xnor2_4 _07054_ (.A(_05604_),
    .B(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__xnor2_4 _07055_ (.A(_05595_),
    .B(_00185_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _07056_ (.A(net183),
    .B(_00178_),
    .Y(_00188_));
 sky130_fd_sc_hd__o21a_2 _07057_ (.A1(net183),
    .A2(_00177_),
    .B1(_00188_),
    .X(_00189_));
 sky130_fd_sc_hd__inv_2 _07058_ (.A(net136),
    .Y(_00190_));
 sky130_fd_sc_hd__nor2_1 _07059_ (.A(_05671_),
    .B(net189),
    .Y(_00191_));
 sky130_fd_sc_hd__o211ai_1 _07060_ (.A1(_05681_),
    .A2(_00183_),
    .B1(net190),
    .C1(_05737_),
    .Y(_00192_));
 sky130_fd_sc_hd__a211o_1 _07061_ (.A1(net190),
    .A2(_00183_),
    .B1(_00191_),
    .C1(_05737_),
    .X(_00193_));
 sky130_fd_sc_hd__and2_1 _07062_ (.A(_00192_),
    .B(_00193_),
    .X(_00194_));
 sky130_fd_sc_hd__o22a_1 _07063_ (.A1(net170),
    .A2(_00187_),
    .B1(net136),
    .B2(net76),
    .X(_00195_));
 sky130_fd_sc_hd__xnor2_1 _07064_ (.A(net184),
    .B(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__nor2_1 _07065_ (.A(_00169_),
    .B(_00196_),
    .Y(_00197_));
 sky130_fd_sc_hd__xor2_1 _07066_ (.A(_00169_),
    .B(_00196_),
    .X(_00198_));
 sky130_fd_sc_hd__a21o_1 _07067_ (.A1(net190),
    .A2(_00183_),
    .B1(_05681_),
    .X(_00199_));
 sky130_fd_sc_hd__or3_1 _07068_ (.A(_05671_),
    .B(net189),
    .C(_00182_),
    .X(_00200_));
 sky130_fd_sc_hd__nand2_1 _07069_ (.A(_00199_),
    .B(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__xnor2_4 _07070_ (.A(reg1_val[8]),
    .B(_00156_),
    .Y(_00202_));
 sky130_fd_sc_hd__nor2_1 _07071_ (.A(net183),
    .B(_00202_),
    .Y(_00203_));
 sky130_fd_sc_hd__and2_1 _07072_ (.A(net183),
    .B(_00202_),
    .X(_00204_));
 sky130_fd_sc_hd__or2_2 _07073_ (.A(_00203_),
    .B(_00204_),
    .X(_00205_));
 sky130_fd_sc_hd__inv_2 _07074_ (.A(net134),
    .Y(_00206_));
 sky130_fd_sc_hd__nor2_1 _07075_ (.A(_05863_),
    .B(_06474_),
    .Y(_00207_));
 sky130_fd_sc_hd__o21ai_4 _07076_ (.A1(_00154_),
    .A2(_00207_),
    .B1(_05800_),
    .Y(_00208_));
 sky130_fd_sc_hd__or3_2 _07077_ (.A(_05800_),
    .B(_00154_),
    .C(_00207_),
    .X(_00209_));
 sky130_fd_sc_hd__and2_1 _07078_ (.A(_00208_),
    .B(_00209_),
    .X(_00210_));
 sky130_fd_sc_hd__nand2_4 _07079_ (.A(_00208_),
    .B(_00209_),
    .Y(_00211_));
 sky130_fd_sc_hd__and3b_1 _07080_ (.A_N(net186),
    .B(net183),
    .C(_00202_),
    .X(_00212_));
 sky130_fd_sc_hd__a21oi_2 _07081_ (.A1(net186),
    .A2(_00203_),
    .B1(_00212_),
    .Y(_00213_));
 sky130_fd_sc_hd__o22a_1 _07082_ (.A1(net71),
    .A2(net135),
    .B1(net69),
    .B2(net133),
    .X(_00214_));
 sky130_fd_sc_hd__xnor2_1 _07083_ (.A(net186),
    .B(_00214_),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _07084_ (.A(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__a21oi_1 _07085_ (.A1(_00198_),
    .A2(_00216_),
    .B1(_00197_),
    .Y(_00217_));
 sky130_fd_sc_hd__or3_2 _07086_ (.A(reg1_val[26]),
    .B(reg1_val[27]),
    .C(_06468_),
    .X(_00218_));
 sky130_fd_sc_hd__or4_2 _07087_ (.A(reg1_val[28]),
    .B(_06463_),
    .C(_06467_),
    .D(_00218_),
    .X(_00219_));
 sky130_fd_sc_hd__a21oi_1 _07088_ (.A1(net274),
    .A2(_00219_),
    .B1(reg1_val[29]),
    .Y(_00220_));
 sky130_fd_sc_hd__and3_1 _07089_ (.A(reg1_val[29]),
    .B(net274),
    .C(_00219_),
    .X(_00221_));
 sky130_fd_sc_hd__or2_2 _07090_ (.A(_00220_),
    .B(_00221_),
    .X(_00222_));
 sky130_fd_sc_hd__and3_2 _07091_ (.A(net303),
    .B(_05392_),
    .C(net213),
    .X(_00223_));
 sky130_fd_sc_hd__xnor2_4 _07092_ (.A(_06327_),
    .B(_00223_),
    .Y(_00224_));
 sky130_fd_sc_hd__xnor2_1 _07093_ (.A(net219),
    .B(_00223_),
    .Y(_00225_));
 sky130_fd_sc_hd__o31a_2 _07094_ (.A1(_06463_),
    .A2(_06467_),
    .A3(_00218_),
    .B1(net274),
    .X(_00226_));
 sky130_fd_sc_hd__xor2_4 _07095_ (.A(reg1_val[28]),
    .B(_00226_),
    .X(_00227_));
 sky130_fd_sc_hd__or2_1 _07096_ (.A(net121),
    .B(_00227_),
    .X(_00228_));
 sky130_fd_sc_hd__nand2_1 _07097_ (.A(net121),
    .B(_00227_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_4 _07098_ (.A(_00228_),
    .B(_00229_),
    .Y(_00230_));
 sky130_fd_sc_hd__mux2_2 _07099_ (.A0(_00228_),
    .A1(_00229_),
    .S(net68),
    .X(_00231_));
 sky130_fd_sc_hd__o22a_1 _07100_ (.A1(net168),
    .A2(net28),
    .B1(net26),
    .B2(net214),
    .X(_00232_));
 sky130_fd_sc_hd__xor2_1 _07101_ (.A(net68),
    .B(_00232_),
    .X(_00233_));
 sky130_fd_sc_hd__and2b_1 _07102_ (.A_N(_00217_),
    .B(_00233_),
    .X(_00234_));
 sky130_fd_sc_hd__o31a_2 _07103_ (.A1(reg1_val[0]),
    .A2(net301),
    .A3(reg1_val[2]),
    .B1(net274),
    .X(_00235_));
 sky130_fd_sc_hd__xnor2_4 _07104_ (.A(reg1_val[3]),
    .B(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_2 _07105_ (.A(net275),
    .B(_06459_),
    .Y(_00237_));
 sky130_fd_sc_hd__xor2_4 _07106_ (.A(reg1_val[4]),
    .B(_00237_),
    .X(_00238_));
 sky130_fd_sc_hd__nand2_2 _07107_ (.A(net203),
    .B(_00238_),
    .Y(_00239_));
 sky130_fd_sc_hd__or2_1 _07108_ (.A(net203),
    .B(_00238_),
    .X(_00240_));
 sky130_fd_sc_hd__and2_2 _07109_ (.A(_00239_),
    .B(_00240_),
    .X(_00241_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(_00239_),
    .B(_00240_),
    .Y(_00242_));
 sky130_fd_sc_hd__and3_1 _07111_ (.A(_05522_),
    .B(_05595_),
    .C(_00184_),
    .X(_00243_));
 sky130_fd_sc_hd__or3b_1 _07112_ (.A(_05533_),
    .B(_05604_),
    .C_N(_00184_),
    .X(_00244_));
 sky130_fd_sc_hd__a21o_1 _07113_ (.A1(_00182_),
    .A2(_00243_),
    .B1(net189),
    .X(_00245_));
 sky130_fd_sc_hd__xnor2_4 _07114_ (.A(_05154_),
    .B(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__or3b_2 _07115_ (.A(net203),
    .B(_00238_),
    .C_N(net206),
    .X(_00247_));
 sky130_fd_sc_hd__o21a_1 _07116_ (.A1(net206),
    .A2(_00239_),
    .B1(_00247_),
    .X(_00248_));
 sky130_fd_sc_hd__o21ai_2 _07117_ (.A1(net206),
    .A2(_00239_),
    .B1(_00247_),
    .Y(_00249_));
 sky130_fd_sc_hd__a31o_1 _07118_ (.A1(_05595_),
    .A2(_00182_),
    .A3(_00184_),
    .B1(net189),
    .X(_00250_));
 sky130_fd_sc_hd__xnor2_4 _07119_ (.A(_05522_),
    .B(_00250_),
    .Y(_00251_));
 sky130_fd_sc_hd__o22a_1 _07120_ (.A1(net166),
    .A2(net65),
    .B1(net164),
    .B2(_00251_),
    .X(_00252_));
 sky130_fd_sc_hd__xnor2_1 _07121_ (.A(net207),
    .B(_00252_),
    .Y(_00253_));
 sky130_fd_sc_hd__and3_4 _07122_ (.A(reg1_val[0]),
    .B(reg1_val[31]),
    .C(net303),
    .X(_00254_));
 sky130_fd_sc_hd__xor2_4 _07123_ (.A(net301),
    .B(_00254_),
    .X(_00255_));
 sky130_fd_sc_hd__xnor2_4 _07124_ (.A(net301),
    .B(_00254_),
    .Y(_00256_));
 sky130_fd_sc_hd__and2_1 _07125_ (.A(_05089_),
    .B(_05154_),
    .X(_00257_));
 sky130_fd_sc_hd__nand2_1 _07126_ (.A(_05089_),
    .B(_05154_),
    .Y(_00258_));
 sky130_fd_sc_hd__and3_1 _07127_ (.A(_00182_),
    .B(_00243_),
    .C(_00257_),
    .X(_00259_));
 sky130_fd_sc_hd__and4b_1 _07128_ (.A_N(_05306_),
    .B(_00182_),
    .C(_00243_),
    .D(_00257_),
    .X(_00260_));
 sky130_fd_sc_hd__or4_1 _07129_ (.A(_05306_),
    .B(_00183_),
    .C(_00244_),
    .D(_00258_),
    .X(_00261_));
 sky130_fd_sc_hd__nor2_1 _07130_ (.A(_05241_),
    .B(_05306_),
    .Y(_00262_));
 sky130_fd_sc_hd__a21o_1 _07131_ (.A1(_05230_),
    .A2(_00260_),
    .B1(net189),
    .X(_00263_));
 sky130_fd_sc_hd__xnor2_4 _07132_ (.A(_05012_),
    .B(_00263_),
    .Y(_00264_));
 sky130_fd_sc_hd__and2_4 _07133_ (.A(net300),
    .B(net301),
    .X(_00265_));
 sky130_fd_sc_hd__nand2_4 _07134_ (.A(net300),
    .B(reg1_val[1]),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_2 _07135_ (.A(_05241_),
    .B(net189),
    .Y(_00267_));
 sky130_fd_sc_hd__o41a_1 _07136_ (.A1(_05306_),
    .A2(_00183_),
    .A3(_00244_),
    .A4(_00258_),
    .B1(_05241_),
    .X(_00268_));
 sky130_fd_sc_hd__a211o_2 _07137_ (.A1(_00259_),
    .A2(_00262_),
    .B1(_00268_),
    .C1(net189),
    .X(_00269_));
 sky130_fd_sc_hd__and2_2 _07138_ (.A(_00267_),
    .B(_00269_),
    .X(_00270_));
 sky130_fd_sc_hd__nand2_4 _07139_ (.A(_00267_),
    .B(_00269_),
    .Y(_00271_));
 sky130_fd_sc_hd__o22a_1 _07140_ (.A1(net299),
    .A2(net24),
    .B1(net247),
    .B2(net22),
    .X(_00272_));
 sky130_fd_sc_hd__xnor2_1 _07141_ (.A(net248),
    .B(_00272_),
    .Y(_00273_));
 sky130_fd_sc_hd__nor2_1 _07142_ (.A(_00253_),
    .B(_00273_),
    .Y(_00274_));
 sky130_fd_sc_hd__o21a_1 _07143_ (.A1(net302),
    .A2(reg1_val[1]),
    .B1(net275),
    .X(_00275_));
 sky130_fd_sc_hd__xnor2_4 _07144_ (.A(reg1_val[2]),
    .B(_00275_),
    .Y(_00276_));
 sky130_fd_sc_hd__and2_1 _07145_ (.A(net249),
    .B(_00276_),
    .X(_00277_));
 sky130_fd_sc_hd__nand2_1 _07146_ (.A(_00256_),
    .B(_00276_),
    .Y(_00278_));
 sky130_fd_sc_hd__nor2_1 _07147_ (.A(net249),
    .B(_00276_),
    .Y(_00279_));
 sky130_fd_sc_hd__or2_1 _07148_ (.A(_00256_),
    .B(_00276_),
    .X(_00280_));
 sky130_fd_sc_hd__nor2_2 _07149_ (.A(_00277_),
    .B(_00279_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _07150_ (.A(_00278_),
    .B(_00280_),
    .Y(_00282_));
 sky130_fd_sc_hd__a31o_4 _07151_ (.A1(_00182_),
    .A2(_00243_),
    .A3(_00257_),
    .B1(net189),
    .X(_00283_));
 sky130_fd_sc_hd__xnor2_4 _07152_ (.A(_05306_),
    .B(_00283_),
    .Y(_00284_));
 sky130_fd_sc_hd__xor2_4 _07153_ (.A(_05306_),
    .B(_00283_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_2 _07154_ (.A0(_00278_),
    .A1(_00280_),
    .S(net205),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_2 _07155_ (.A0(_00277_),
    .A1(_00279_),
    .S(net205),
    .X(_00287_));
 sky130_fd_sc_hd__a31o_1 _07156_ (.A1(_05154_),
    .A2(_00182_),
    .A3(_00243_),
    .B1(net189),
    .X(_00288_));
 sky130_fd_sc_hd__xnor2_4 _07157_ (.A(_05089_),
    .B(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__o22a_1 _07158_ (.A1(net162),
    .A2(net61),
    .B1(net160),
    .B2(net58),
    .X(_00290_));
 sky130_fd_sc_hd__xnor2_1 _07159_ (.A(net203),
    .B(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__xnor2_1 _07160_ (.A(_00253_),
    .B(_00273_),
    .Y(_00292_));
 sky130_fd_sc_hd__nor2_1 _07161_ (.A(_00291_),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__xnor2_1 _07162_ (.A(_00217_),
    .B(_00233_),
    .Y(_00294_));
 sky130_fd_sc_hd__o21a_1 _07163_ (.A1(_00274_),
    .A2(_00293_),
    .B1(_00294_),
    .X(_00295_));
 sky130_fd_sc_hd__or2_1 _07164_ (.A(_00234_),
    .B(_00295_),
    .X(_00296_));
 sky130_fd_sc_hd__nand2_2 _07165_ (.A(net274),
    .B(_06462_),
    .Y(_00297_));
 sky130_fd_sc_hd__xor2_4 _07166_ (.A(reg1_val[13]),
    .B(_00297_),
    .X(_00298_));
 sky130_fd_sc_hd__xnor2_1 _07167_ (.A(_06009_),
    .B(_00164_),
    .Y(_00299_));
 sky130_fd_sc_hd__xnor2_4 _07168_ (.A(_06020_),
    .B(_00164_),
    .Y(_00300_));
 sky130_fd_sc_hd__o31a_2 _07169_ (.A1(reg1_val[10]),
    .A2(reg1_val[11]),
    .A3(_06461_),
    .B1(net275),
    .X(_00301_));
 sky130_fd_sc_hd__xnor2_4 _07170_ (.A(reg1_val[12]),
    .B(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__and2_1 _07171_ (.A(net172),
    .B(_00302_),
    .X(_00303_));
 sky130_fd_sc_hd__nor2_4 _07172_ (.A(net172),
    .B(_00302_),
    .Y(_00304_));
 sky130_fd_sc_hd__nor2_4 _07173_ (.A(_00303_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__or2_4 _07174_ (.A(_00303_),
    .B(_00304_),
    .X(_00306_));
 sky130_fd_sc_hd__or4_4 _07175_ (.A(_06476_),
    .B(_06499_),
    .C(_00147_),
    .D(_00150_),
    .X(_00307_));
 sky130_fd_sc_hd__o31a_2 _07176_ (.A1(_06149_),
    .A2(_06194_),
    .A3(_00307_),
    .B1(net190),
    .X(_00308_));
 sky130_fd_sc_hd__o41a_2 _07177_ (.A1(_06101_),
    .A2(_06149_),
    .A3(_06194_),
    .A4(_00307_),
    .B1(net190),
    .X(_00309_));
 sky130_fd_sc_hd__xor2_4 _07178_ (.A(_06071_),
    .B(_00309_),
    .X(_00310_));
 sky130_fd_sc_hd__clkinv_4 _07179_ (.A(net97),
    .Y(_00311_));
 sky130_fd_sc_hd__and2b_1 _07180_ (.A_N(net130),
    .B(_00303_),
    .X(_00312_));
 sky130_fd_sc_hd__a21oi_4 _07181_ (.A1(net130),
    .A2(_00304_),
    .B1(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__a21o_4 _07182_ (.A1(net130),
    .A2(_00304_),
    .B1(_00312_),
    .X(_00314_));
 sky130_fd_sc_hd__a22o_1 _07183_ (.A1(net99),
    .A2(_00305_),
    .B1(net97),
    .B2(_00314_),
    .X(_00315_));
 sky130_fd_sc_hd__xor2_1 _07184_ (.A(net130),
    .B(_00315_),
    .X(_00316_));
 sky130_fd_sc_hd__o21a_1 _07185_ (.A1(reg1_val[13]),
    .A2(_06462_),
    .B1(net275),
    .X(_00317_));
 sky130_fd_sc_hd__o31a_4 _07186_ (.A1(reg1_val[13]),
    .A2(reg1_val[14]),
    .A3(_06462_),
    .B1(net275),
    .X(_00318_));
 sky130_fd_sc_hd__xor2_4 _07187_ (.A(reg1_val[15]),
    .B(_00318_),
    .X(_00319_));
 sky130_fd_sc_hd__xnor2_4 _07188_ (.A(reg1_val[15]),
    .B(_00318_),
    .Y(_00320_));
 sky130_fd_sc_hd__xnor2_4 _07189_ (.A(reg1_val[14]),
    .B(_00317_),
    .Y(_00321_));
 sky130_fd_sc_hd__xnor2_4 _07190_ (.A(net130),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__xor2_4 _07191_ (.A(_06101_),
    .B(_00308_),
    .X(_00323_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(_06101_),
    .B(_00308_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand3_1 _07193_ (.A(net130),
    .B(_00319_),
    .C(_00321_),
    .Y(_00325_));
 sky130_fd_sc_hd__or3_2 _07194_ (.A(net130),
    .B(_00319_),
    .C(_00321_),
    .X(_00326_));
 sky130_fd_sc_hd__and2_2 _07195_ (.A(_00325_),
    .B(_00326_),
    .X(_00327_));
 sky130_fd_sc_hd__o21a_1 _07196_ (.A1(_06194_),
    .A2(_00307_),
    .B1(net190),
    .X(_00328_));
 sky130_fd_sc_hd__xnor2_4 _07197_ (.A(_06149_),
    .B(_00328_),
    .Y(_00329_));
 sky130_fd_sc_hd__o22a_1 _07198_ (.A1(net96),
    .A2(net94),
    .B1(net55),
    .B2(net92),
    .X(_00330_));
 sky130_fd_sc_hd__xnor2_1 _07199_ (.A(net127),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__or2_2 _07200_ (.A(_00316_),
    .B(_00331_),
    .X(_00332_));
 sky130_fd_sc_hd__o22a_1 _07201_ (.A1(net108),
    .A2(net103),
    .B1(net69),
    .B2(net107),
    .X(_00333_));
 sky130_fd_sc_hd__xnor2_1 _07202_ (.A(net173),
    .B(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__o22a_1 _07203_ (.A1(net77),
    .A2(net136),
    .B1(net62),
    .B2(net170),
    .X(_00335_));
 sky130_fd_sc_hd__xnor2_1 _07204_ (.A(net184),
    .B(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__xor2_1 _07205_ (.A(_00334_),
    .B(_00336_),
    .X(_00337_));
 sky130_fd_sc_hd__o22a_1 _07206_ (.A1(net74),
    .A2(net135),
    .B1(net133),
    .B2(net71),
    .X(_00338_));
 sky130_fd_sc_hd__xnor2_1 _07207_ (.A(net188),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2b_1 _07208_ (.A_N(_00339_),
    .B(_00337_),
    .Y(_00340_));
 sky130_fd_sc_hd__xnor2_1 _07209_ (.A(_00337_),
    .B(_00339_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2b_1 _07210_ (.A_N(_00332_),
    .B(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__o22a_1 _07211_ (.A1(net22),
    .A2(net162),
    .B1(net61),
    .B2(net160),
    .X(_00343_));
 sky130_fd_sc_hd__xnor2_1 _07212_ (.A(net203),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__inv_2 _07213_ (.A(_00344_),
    .Y(_00345_));
 sky130_fd_sc_hd__o22a_1 _07214_ (.A1(_00246_),
    .A2(net164),
    .B1(net58),
    .B2(net166),
    .X(_00346_));
 sky130_fd_sc_hd__xnor2_1 _07215_ (.A(net207),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__a31o_1 _07216_ (.A1(_05012_),
    .A2(_05230_),
    .A3(_00260_),
    .B1(net189),
    .X(_00348_));
 sky130_fd_sc_hd__xnor2_4 _07217_ (.A(_04947_),
    .B(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__o22a_1 _07218_ (.A1(net24),
    .A2(net247),
    .B1(net20),
    .B2(net299),
    .X(_00350_));
 sky130_fd_sc_hd__xnor2_1 _07219_ (.A(net248),
    .B(_00350_),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_1 _07220_ (.A(_00347_),
    .B(_00351_),
    .Y(_00352_));
 sky130_fd_sc_hd__xor2_1 _07221_ (.A(_00347_),
    .B(_00351_),
    .X(_00353_));
 sky130_fd_sc_hd__xnor2_1 _07222_ (.A(_00344_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__xnor2_1 _07223_ (.A(_00332_),
    .B(_00341_),
    .Y(_00355_));
 sky130_fd_sc_hd__a21bo_1 _07224_ (.A1(_00354_),
    .A2(_00355_),
    .B1_N(_00342_),
    .X(_00356_));
 sky130_fd_sc_hd__xnor2_1 _07225_ (.A(_00143_),
    .B(_00296_),
    .Y(_00357_));
 sky130_fd_sc_hd__and2b_1 _07226_ (.A_N(_00357_),
    .B(_00356_),
    .X(_00358_));
 sky130_fd_sc_hd__a21o_2 _07227_ (.A1(_00143_),
    .A2(_00296_),
    .B1(_00358_),
    .X(_00359_));
 sky130_fd_sc_hd__o22a_1 _07228_ (.A1(net170),
    .A2(net65),
    .B1(net62),
    .B2(net136),
    .X(_00360_));
 sky130_fd_sc_hd__xnor2_1 _07229_ (.A(net184),
    .B(_00360_),
    .Y(_00361_));
 sky130_fd_sc_hd__o22a_1 _07230_ (.A1(net107),
    .A2(net72),
    .B1(net69),
    .B2(net103),
    .X(_00362_));
 sky130_fd_sc_hd__xnor2_1 _07231_ (.A(net173),
    .B(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__nor2_1 _07232_ (.A(_00361_),
    .B(_00363_),
    .Y(_00364_));
 sky130_fd_sc_hd__and2_1 _07233_ (.A(_00361_),
    .B(_00363_),
    .X(_00365_));
 sky130_fd_sc_hd__nor2_1 _07234_ (.A(_00364_),
    .B(_00365_),
    .Y(_00366_));
 sky130_fd_sc_hd__o22a_1 _07235_ (.A1(net77),
    .A2(net135),
    .B1(net133),
    .B2(net75),
    .X(_00367_));
 sky130_fd_sc_hd__xnor2_2 _07236_ (.A(net188),
    .B(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__xnor2_2 _07237_ (.A(_00366_),
    .B(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__o22a_1 _07238_ (.A1(net24),
    .A2(net162),
    .B1(net160),
    .B2(net22),
    .X(_00370_));
 sky130_fd_sc_hd__xnor2_1 _07239_ (.A(net203),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _07240_ (.A(_00371_),
    .Y(_00372_));
 sky130_fd_sc_hd__o22a_2 _07241_ (.A1(net166),
    .A2(net61),
    .B1(net58),
    .B2(net164),
    .X(_00373_));
 sky130_fd_sc_hd__xnor2_4 _07242_ (.A(net207),
    .B(_00373_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _07243_ (.A(_04947_),
    .B(_05012_),
    .Y(_00375_));
 sky130_fd_sc_hd__o31a_2 _07244_ (.A1(_05241_),
    .A2(_00261_),
    .A3(_00375_),
    .B1(net190),
    .X(_00376_));
 sky130_fd_sc_hd__xnor2_4 _07245_ (.A(_05446_),
    .B(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__o22a_2 _07246_ (.A1(net247),
    .A2(net20),
    .B1(net18),
    .B2(net299),
    .X(_00378_));
 sky130_fd_sc_hd__xnor2_4 _07247_ (.A(net248),
    .B(_00378_),
    .Y(_00379_));
 sky130_fd_sc_hd__nor2_1 _07248_ (.A(_00374_),
    .B(_00379_),
    .Y(_00380_));
 sky130_fd_sc_hd__xor2_4 _07249_ (.A(_00374_),
    .B(_00379_),
    .X(_00381_));
 sky130_fd_sc_hd__xnor2_2 _07250_ (.A(_00372_),
    .B(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__o22a_1 _07251_ (.A1(net108),
    .A2(net98),
    .B1(net56),
    .B2(net104),
    .X(_00383_));
 sky130_fd_sc_hd__xnor2_1 _07252_ (.A(net129),
    .B(_00383_),
    .Y(_00384_));
 sky130_fd_sc_hd__o41a_2 _07253_ (.A1(reg1_val[13]),
    .A2(reg1_val[14]),
    .A3(reg1_val[15]),
    .A4(_06462_),
    .B1(net274),
    .X(_00385_));
 sky130_fd_sc_hd__o21ai_1 _07254_ (.A1(reg1_val[16]),
    .A2(_06463_),
    .B1(net274),
    .Y(_00386_));
 sky130_fd_sc_hd__xnor2_1 _07255_ (.A(reg1_val[17]),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_4 _07256_ (.A(net90),
    .Y(_00388_));
 sky130_fd_sc_hd__xnor2_4 _07257_ (.A(reg1_val[16]),
    .B(_00385_),
    .Y(_00389_));
 sky130_fd_sc_hd__or2_1 _07258_ (.A(net126),
    .B(_00389_),
    .X(_00390_));
 sky130_fd_sc_hd__nand2_2 _07259_ (.A(net126),
    .B(_00389_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_4 _07260_ (.A(_00390_),
    .B(_00391_),
    .Y(_00392_));
 sky130_fd_sc_hd__nor2_1 _07261_ (.A(net88),
    .B(_00390_),
    .Y(_00393_));
 sky130_fd_sc_hd__mux2_1 _07262_ (.A0(_00390_),
    .A1(_00391_),
    .S(net88),
    .X(_00394_));
 sky130_fd_sc_hd__o22a_1 _07263_ (.A1(net93),
    .A2(net52),
    .B1(net50),
    .B2(net91),
    .X(_00395_));
 sky130_fd_sc_hd__xnor2_1 _07264_ (.A(net89),
    .B(_00395_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2b_1 _07265_ (.A_N(_00384_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2b_1 _07266_ (.A_N(_00396_),
    .B(_00384_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_00397_),
    .B(_00398_),
    .Y(_00399_));
 sky130_fd_sc_hd__o22a_1 _07268_ (.A1(net100),
    .A2(net95),
    .B1(net54),
    .B2(net57),
    .X(_00400_));
 sky130_fd_sc_hd__xnor2_2 _07269_ (.A(net126),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__xnor2_2 _07270_ (.A(_00399_),
    .B(_00401_),
    .Y(_00402_));
 sky130_fd_sc_hd__nor2_1 _07271_ (.A(_00382_),
    .B(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__xnor2_2 _07272_ (.A(_00382_),
    .B(_00402_),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_2 _07273_ (.A(_00404_),
    .Y(_00405_));
 sky130_fd_sc_hd__xor2_2 _07274_ (.A(_00369_),
    .B(_00404_),
    .X(_00406_));
 sky130_fd_sc_hd__o21a_1 _07275_ (.A1(reg1_val[29]),
    .A2(_00219_),
    .B1(net274),
    .X(_00407_));
 sky130_fd_sc_hd__xnor2_4 _07276_ (.A(reg1_val[30]),
    .B(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__xnor2_4 _07277_ (.A(net67),
    .B(_00408_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2_2 _07278_ (.A(net214),
    .B(net16),
    .Y(_00410_));
 sky130_fd_sc_hd__xnor2_4 _07279_ (.A(_06322_),
    .B(_06488_),
    .Y(_00411_));
 sky130_fd_sc_hd__o22a_1 _07280_ (.A1(net168),
    .A2(net26),
    .B1(net159),
    .B2(net28),
    .X(_00412_));
 sky130_fd_sc_hd__xnor2_2 _07281_ (.A(net68),
    .B(_00412_),
    .Y(_00413_));
 sky130_fd_sc_hd__xor2_2 _07282_ (.A(_00410_),
    .B(_00413_),
    .X(_00414_));
 sky130_fd_sc_hd__o21ai_1 _07283_ (.A1(_00334_),
    .A2(_00336_),
    .B1(_00340_),
    .Y(_00415_));
 sky130_fd_sc_hd__o22a_1 _07284_ (.A1(net104),
    .A2(net98),
    .B1(net56),
    .B2(net100),
    .X(_00416_));
 sky130_fd_sc_hd__xnor2_1 _07285_ (.A(net129),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__o22a_1 _07286_ (.A1(_00311_),
    .A2(net95),
    .B1(net93),
    .B2(net54),
    .X(_00418_));
 sky130_fd_sc_hd__xnor2_1 _07287_ (.A(net126),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__nor2_1 _07288_ (.A(_00417_),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__a21oi_1 _07289_ (.A1(_00345_),
    .A2(_00353_),
    .B1(_00352_),
    .Y(_00421_));
 sky130_fd_sc_hd__and2b_1 _07290_ (.A_N(_00421_),
    .B(_00420_),
    .X(_00422_));
 sky130_fd_sc_hd__xnor2_1 _07291_ (.A(_00420_),
    .B(_00421_),
    .Y(_00423_));
 sky130_fd_sc_hd__and2_1 _07292_ (.A(_00415_),
    .B(_00423_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_1 _07293_ (.A(_00415_),
    .B(_00423_),
    .Y(_00425_));
 sky130_fd_sc_hd__or2_1 _07294_ (.A(_00424_),
    .B(_00425_),
    .X(_00426_));
 sky130_fd_sc_hd__xnor2_1 _07295_ (.A(_00406_),
    .B(_00414_),
    .Y(_00427_));
 sky130_fd_sc_hd__o32a_2 _07296_ (.A1(_00424_),
    .A2(_00425_),
    .A3(_00427_),
    .B1(_00414_),
    .B2(_00406_),
    .X(_00428_));
 sky130_fd_sc_hd__o21ai_2 _07297_ (.A1(_06463_),
    .A2(_06465_),
    .B1(net274),
    .Y(_00429_));
 sky130_fd_sc_hd__o31a_2 _07298_ (.A1(reg1_val[18]),
    .A2(_06463_),
    .A3(_06465_),
    .B1(net274),
    .X(_00430_));
 sky130_fd_sc_hd__xor2_4 _07299_ (.A(reg1_val[19]),
    .B(_00430_),
    .X(_00431_));
 sky130_fd_sc_hd__xnor2_4 _07300_ (.A(reg1_val[18]),
    .B(_00429_),
    .Y(_00432_));
 sky130_fd_sc_hd__xnor2_4 _07301_ (.A(net88),
    .B(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__a21o_1 _07302_ (.A1(net190),
    .A2(_00307_),
    .B1(_06194_),
    .X(_00434_));
 sky130_fd_sc_hd__nand3_2 _07303_ (.A(_06194_),
    .B(net190),
    .C(_00307_),
    .Y(_00435_));
 sky130_fd_sc_hd__and2_4 _07304_ (.A(_00434_),
    .B(_00435_),
    .X(_00436_));
 sky130_fd_sc_hd__nand2_4 _07305_ (.A(_00434_),
    .B(_00435_),
    .Y(_00437_));
 sky130_fd_sc_hd__or3b_4 _07306_ (.A(net89),
    .B(_00432_),
    .C_N(net85),
    .X(_00438_));
 sky130_fd_sc_hd__nand3b_4 _07307_ (.A_N(net85),
    .B(_00432_),
    .C(net89),
    .Y(_00439_));
 sky130_fd_sc_hd__and2_1 _07308_ (.A(_00438_),
    .B(_00439_),
    .X(_00440_));
 sky130_fd_sc_hd__o31a_4 _07309_ (.A1(_06476_),
    .A2(_06499_),
    .A3(_00147_),
    .B1(net190),
    .X(_00441_));
 sky130_fd_sc_hd__a211o_2 _07310_ (.A1(_06273_),
    .A2(_00148_),
    .B1(_06474_),
    .C1(_06238_),
    .X(_00442_));
 sky130_fd_sc_hd__a211o_2 _07311_ (.A1(_06272_),
    .A2(_06473_),
    .B1(_00441_),
    .C1(_06247_),
    .X(_00443_));
 sky130_fd_sc_hd__and2_2 _07312_ (.A(_00442_),
    .B(_00443_),
    .X(_00444_));
 sky130_fd_sc_hd__nand2_8 _07313_ (.A(_00442_),
    .B(_00443_),
    .Y(_00445_));
 sky130_fd_sc_hd__o22a_1 _07314_ (.A1(net48),
    .A2(net83),
    .B1(net13),
    .B2(net81),
    .X(_00446_));
 sky130_fd_sc_hd__xnor2_1 _07315_ (.A(net85),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__xnor2_4 _07316_ (.A(reg1_val[20]),
    .B(_06496_),
    .Y(_00448_));
 sky130_fd_sc_hd__xnor2_4 _07317_ (.A(net86),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__xnor2_4 _07318_ (.A(_06273_),
    .B(_00441_),
    .Y(_00450_));
 sky130_fd_sc_hd__xnor2_4 _07319_ (.A(_06272_),
    .B(_00441_),
    .Y(_00451_));
 sky130_fd_sc_hd__a21oi_4 _07320_ (.A1(net87),
    .A2(_00448_),
    .B1(_06504_),
    .Y(_00452_));
 sky130_fd_sc_hd__o21a_4 _07321_ (.A1(net86),
    .A2(_00448_),
    .B1(net112),
    .X(_00453_));
 sky130_fd_sc_hd__or2_2 _07322_ (.A(_00452_),
    .B(_00453_),
    .X(_00454_));
 sky130_fd_sc_hd__o31a_4 _07323_ (.A1(_06284_),
    .A2(_06476_),
    .A3(_06499_),
    .B1(net190),
    .X(_00455_));
 sky130_fd_sc_hd__xnor2_4 _07324_ (.A(_06278_),
    .B(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__xnor2_4 _07325_ (.A(_06279_),
    .B(_00455_),
    .Y(_00457_));
 sky130_fd_sc_hd__o22a_1 _07326_ (.A1(net46),
    .A2(net124),
    .B1(net11),
    .B2(net122),
    .X(_00458_));
 sky130_fd_sc_hd__xnor2_1 _07327_ (.A(net111),
    .B(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__and2_1 _07328_ (.A(_00447_),
    .B(_00459_),
    .X(_00460_));
 sky130_fd_sc_hd__nor2_1 _07329_ (.A(_00447_),
    .B(_00459_),
    .Y(_00461_));
 sky130_fd_sc_hd__nor2_1 _07330_ (.A(_00460_),
    .B(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__o22a_1 _07331_ (.A1(net80),
    .A2(net143),
    .B1(net33),
    .B2(net141),
    .X(_00463_));
 sky130_fd_sc_hd__xnor2_1 _07332_ (.A(net115),
    .B(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__o22a_1 _07333_ (.A1(net38),
    .A2(net174),
    .B1(net36),
    .B2(net159),
    .X(_00465_));
 sky130_fd_sc_hd__xnor2_1 _07334_ (.A(net121),
    .B(_00465_),
    .Y(_00466_));
 sky130_fd_sc_hd__xor2_1 _07335_ (.A(_00464_),
    .B(_00466_),
    .X(_00467_));
 sky130_fd_sc_hd__o22a_1 _07336_ (.A1(net31),
    .A2(net139),
    .B1(net30),
    .B2(net147),
    .X(_00468_));
 sky130_fd_sc_hd__xnor2_1 _07337_ (.A(net118),
    .B(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__and2_1 _07338_ (.A(_00467_),
    .B(_00469_),
    .X(_00470_));
 sky130_fd_sc_hd__a21o_1 _07339_ (.A1(_00464_),
    .A2(_00466_),
    .B1(_00470_),
    .X(_00471_));
 sky130_fd_sc_hd__o22a_1 _07340_ (.A1(net91),
    .A2(net52),
    .B1(net50),
    .B2(net83),
    .X(_00472_));
 sky130_fd_sc_hd__xnor2_1 _07341_ (.A(net89),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__o22a_1 _07342_ (.A1(net145),
    .A2(net11),
    .B1(net122),
    .B2(net46),
    .X(_00474_));
 sky130_fd_sc_hd__xnor2_1 _07343_ (.A(net111),
    .B(_00474_),
    .Y(_00475_));
 sky130_fd_sc_hd__xor2_1 _07344_ (.A(_00473_),
    .B(_00475_),
    .X(_00476_));
 sky130_fd_sc_hd__o22a_1 _07345_ (.A1(net48),
    .A2(net81),
    .B1(net124),
    .B2(net13),
    .X(_00477_));
 sky130_fd_sc_hd__xnor2_1 _07346_ (.A(net86),
    .B(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _07347_ (.A(_00476_),
    .B(_00478_),
    .Y(_00479_));
 sky130_fd_sc_hd__a21bo_1 _07348_ (.A1(_00473_),
    .A2(_00475_),
    .B1_N(_00479_),
    .X(_00480_));
 sky130_fd_sc_hd__xnor2_1 _07349_ (.A(_00462_),
    .B(_00471_),
    .Y(_00481_));
 sky130_fd_sc_hd__and2b_1 _07350_ (.A_N(_00481_),
    .B(_00480_),
    .X(_00482_));
 sky130_fd_sc_hd__a21oi_2 _07351_ (.A1(_00462_),
    .A2(_00471_),
    .B1(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__or2_1 _07352_ (.A(_00428_),
    .B(_00483_),
    .X(_00484_));
 sky130_fd_sc_hd__xor2_4 _07353_ (.A(_00428_),
    .B(_00483_),
    .X(_00485_));
 sky130_fd_sc_hd__xnor2_4 _07354_ (.A(_00359_),
    .B(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__and2_1 _07355_ (.A(_00417_),
    .B(_00419_),
    .X(_00487_));
 sky130_fd_sc_hd__nor2_1 _07356_ (.A(_00420_),
    .B(_00487_),
    .Y(_00488_));
 sky130_fd_sc_hd__o22a_1 _07357_ (.A1(net80),
    .A2(net140),
    .B1(net139),
    .B2(net34),
    .X(_00489_));
 sky130_fd_sc_hd__xor2_1 _07358_ (.A(net115),
    .B(_00489_),
    .X(_00490_));
 sky130_fd_sc_hd__o22a_1 _07359_ (.A1(net36),
    .A2(net168),
    .B1(net159),
    .B2(net38),
    .X(_00491_));
 sky130_fd_sc_hd__xnor2_1 _07360_ (.A(_06472_),
    .B(_00491_),
    .Y(_00492_));
 sky130_fd_sc_hd__nor2_1 _07361_ (.A(_00490_),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__xor2_1 _07362_ (.A(_00490_),
    .B(_00492_),
    .X(_00494_));
 sky130_fd_sc_hd__o22a_1 _07363_ (.A1(net147),
    .A2(net31),
    .B1(net30),
    .B2(net174),
    .X(_00495_));
 sky130_fd_sc_hd__xnor2_1 _07364_ (.A(_06482_),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__a21o_1 _07365_ (.A1(_00494_),
    .A2(_00496_),
    .B1(_00493_),
    .X(_00497_));
 sky130_fd_sc_hd__o22a_1 _07366_ (.A1(net52),
    .A2(net83),
    .B1(net81),
    .B2(net51),
    .X(_00498_));
 sky130_fd_sc_hd__xnor2_1 _07367_ (.A(net88),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__o22a_1 _07368_ (.A1(net144),
    .A2(net46),
    .B1(net11),
    .B2(net142),
    .X(_00500_));
 sky130_fd_sc_hd__xnor2_1 _07369_ (.A(net111),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__and2_1 _07370_ (.A(_00499_),
    .B(_00501_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_1 _07371_ (.A(_00499_),
    .B(_00501_),
    .Y(_00503_));
 sky130_fd_sc_hd__nor2_1 _07372_ (.A(_00502_),
    .B(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__o22a_1 _07373_ (.A1(net48),
    .A2(net124),
    .B1(net122),
    .B2(net14),
    .X(_00505_));
 sky130_fd_sc_hd__xnor2_1 _07374_ (.A(net86),
    .B(_00505_),
    .Y(_00506_));
 sky130_fd_sc_hd__a21o_1 _07375_ (.A1(_00504_),
    .A2(_00506_),
    .B1(_00502_),
    .X(_00507_));
 sky130_fd_sc_hd__xnor2_1 _07376_ (.A(_00488_),
    .B(_00497_),
    .Y(_00508_));
 sky130_fd_sc_hd__and2b_1 _07377_ (.A_N(_00508_),
    .B(_00507_),
    .X(_00509_));
 sky130_fd_sc_hd__a21oi_1 _07378_ (.A1(_00488_),
    .A2(_00497_),
    .B1(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__xnor2_1 _07379_ (.A(_00354_),
    .B(_00355_),
    .Y(_00511_));
 sky130_fd_sc_hd__nor2_1 _07380_ (.A(_00467_),
    .B(_00469_),
    .Y(_00512_));
 sky130_fd_sc_hd__nor2_1 _07381_ (.A(_00470_),
    .B(_00512_),
    .Y(_00513_));
 sky130_fd_sc_hd__and2b_1 _07382_ (.A_N(_00511_),
    .B(_00513_),
    .X(_00514_));
 sky130_fd_sc_hd__nor3_1 _07383_ (.A(_00274_),
    .B(_00293_),
    .C(_00294_),
    .Y(_00515_));
 sky130_fd_sc_hd__nor2_1 _07384_ (.A(_00295_),
    .B(_00515_),
    .Y(_00516_));
 sky130_fd_sc_hd__xnor2_1 _07385_ (.A(_00511_),
    .B(_00513_),
    .Y(_00517_));
 sky130_fd_sc_hd__a21oi_1 _07386_ (.A1(_00516_),
    .A2(_00517_),
    .B1(_00514_),
    .Y(_00518_));
 sky130_fd_sc_hd__or2_1 _07387_ (.A(_00476_),
    .B(_00478_),
    .X(_00519_));
 sky130_fd_sc_hd__nand2_2 _07388_ (.A(_00479_),
    .B(_00519_),
    .Y(_00520_));
 sky130_fd_sc_hd__nor2_1 _07389_ (.A(net214),
    .B(net28),
    .Y(_00521_));
 sky130_fd_sc_hd__a21o_1 _07390_ (.A1(_00267_),
    .A2(_00269_),
    .B1(net299),
    .X(_00522_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(_00265_),
    .B(_00284_),
    .Y(_00523_));
 sky130_fd_sc_hd__a21o_1 _07392_ (.A1(_00522_),
    .A2(_00523_),
    .B1(net248),
    .X(_00524_));
 sky130_fd_sc_hd__nand3_1 _07393_ (.A(net248),
    .B(_00522_),
    .C(_00523_),
    .Y(_00525_));
 sky130_fd_sc_hd__o22a_1 _07394_ (.A1(net77),
    .A2(net164),
    .B1(net62),
    .B2(net166),
    .X(_00526_));
 sky130_fd_sc_hd__xor2_1 _07395_ (.A(net206),
    .B(_00526_),
    .X(_00527_));
 sky130_fd_sc_hd__nand3_2 _07396_ (.A(_00524_),
    .B(_00525_),
    .C(_00527_),
    .Y(_00528_));
 sky130_fd_sc_hd__o22a_1 _07397_ (.A1(net65),
    .A2(net160),
    .B1(_00289_),
    .B2(net162),
    .X(_00529_));
 sky130_fd_sc_hd__xor2_1 _07398_ (.A(net204),
    .B(_00529_),
    .X(_00530_));
 sky130_fd_sc_hd__a21o_1 _07399_ (.A1(_00524_),
    .A2(_00525_),
    .B1(_00527_),
    .X(_00531_));
 sky130_fd_sc_hd__nand3_2 _07400_ (.A(_00528_),
    .B(_00530_),
    .C(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _07401_ (.A(_00528_),
    .B(_00532_),
    .Y(_00533_));
 sky130_fd_sc_hd__o21a_1 _07402_ (.A1(net214),
    .A2(net28),
    .B1(net68),
    .X(_00534_));
 sky130_fd_sc_hd__a31o_1 _07403_ (.A1(_00521_),
    .A2(_00528_),
    .A3(_00532_),
    .B1(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__o22a_1 _07404_ (.A1(net170),
    .A2(net76),
    .B1(net73),
    .B2(net136),
    .X(_00536_));
 sky130_fd_sc_hd__xnor2_1 _07405_ (.A(net184),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__o22a_1 _07406_ (.A1(net135),
    .A2(net69),
    .B1(net133),
    .B2(net109),
    .X(_00538_));
 sky130_fd_sc_hd__xnor2_1 _07407_ (.A(net186),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__or2_1 _07408_ (.A(_00537_),
    .B(_00539_),
    .X(_00540_));
 sky130_fd_sc_hd__xnor2_1 _07409_ (.A(_00198_),
    .B(_00216_),
    .Y(_00541_));
 sky130_fd_sc_hd__nor2_1 _07410_ (.A(_00540_),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__xor2_1 _07411_ (.A(_00291_),
    .B(_00292_),
    .X(_00543_));
 sky130_fd_sc_hd__xor2_1 _07412_ (.A(_00540_),
    .B(_00541_),
    .X(_00544_));
 sky130_fd_sc_hd__a21o_2 _07413_ (.A1(_00543_),
    .A2(_00544_),
    .B1(_00542_),
    .X(_00545_));
 sky130_fd_sc_hd__xnor2_2 _07414_ (.A(_00520_),
    .B(_00535_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2b_1 _07415_ (.A_N(_00546_),
    .B(_00545_),
    .Y(_00547_));
 sky130_fd_sc_hd__o21ai_2 _07416_ (.A1(_00520_),
    .A2(_00535_),
    .B1(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__xnor2_1 _07417_ (.A(_00510_),
    .B(_00518_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2b_1 _07418_ (.A_N(_00549_),
    .B(_00548_),
    .Y(_00550_));
 sky130_fd_sc_hd__o21a_2 _07419_ (.A1(_00510_),
    .A2(_00518_),
    .B1(_00550_),
    .X(_00551_));
 sky130_fd_sc_hd__xor2_1 _07420_ (.A(_00426_),
    .B(_00427_),
    .X(_00552_));
 sky130_fd_sc_hd__xnor2_1 _07421_ (.A(_00480_),
    .B(_00481_),
    .Y(_00553_));
 sky130_fd_sc_hd__and2_1 _07422_ (.A(_00552_),
    .B(_00553_),
    .X(_00554_));
 sky130_fd_sc_hd__xnor2_1 _07423_ (.A(_00356_),
    .B(_00357_),
    .Y(_00555_));
 sky130_fd_sc_hd__xor2_1 _07424_ (.A(_00552_),
    .B(_00553_),
    .X(_00556_));
 sky130_fd_sc_hd__a21o_1 _07425_ (.A1(_00555_),
    .A2(_00556_),
    .B1(_00554_),
    .X(_00557_));
 sky130_fd_sc_hd__xnor2_2 _07426_ (.A(_00486_),
    .B(_00551_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2b_1 _07427_ (.A_N(_00558_),
    .B(_00557_),
    .Y(_00559_));
 sky130_fd_sc_hd__o21ai_4 _07428_ (.A1(_00486_),
    .A2(_00551_),
    .B1(_00559_),
    .Y(_00560_));
 sky130_fd_sc_hd__o22a_1 _07429_ (.A1(net24),
    .A2(net160),
    .B1(net20),
    .B2(net162),
    .X(_00561_));
 sky130_fd_sc_hd__xnor2_1 _07430_ (.A(net204),
    .B(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _07431_ (.A(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__o22a_2 _07432_ (.A1(net166),
    .A2(net22),
    .B1(net61),
    .B2(net164),
    .X(_00564_));
 sky130_fd_sc_hd__xnor2_4 _07433_ (.A(net207),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__or4_2 _07434_ (.A(_05241_),
    .B(_05446_),
    .C(_00261_),
    .D(_00375_),
    .X(_00566_));
 sky130_fd_sc_hd__a21oi_4 _07435_ (.A1(net303),
    .A2(_00566_),
    .B1(_05382_),
    .Y(_00567_));
 sky130_fd_sc_hd__a21o_1 _07436_ (.A1(net303),
    .A2(_00566_),
    .B1(_05382_),
    .X(_00568_));
 sky130_fd_sc_hd__o22a_2 _07437_ (.A1(net247),
    .A2(_00377_),
    .B1(net9),
    .B2(net299),
    .X(_00569_));
 sky130_fd_sc_hd__xnor2_4 _07438_ (.A(net248),
    .B(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__nor2_1 _07439_ (.A(_00565_),
    .B(_00570_),
    .Y(_00571_));
 sky130_fd_sc_hd__xor2_4 _07440_ (.A(_00565_),
    .B(_00570_),
    .X(_00572_));
 sky130_fd_sc_hd__xnor2_4 _07441_ (.A(_00563_),
    .B(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__o22a_1 _07442_ (.A1(net69),
    .A2(net98),
    .B1(net56),
    .B2(net108),
    .X(_00574_));
 sky130_fd_sc_hd__xor2_1 _07443_ (.A(net129),
    .B(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__o22a_1 _07444_ (.A1(net57),
    .A2(net52),
    .B1(net50),
    .B2(net93),
    .X(_00576_));
 sky130_fd_sc_hd__xnor2_1 _07445_ (.A(net89),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(_00575_),
    .B(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__or2_1 _07447_ (.A(_00575_),
    .B(_00577_),
    .X(_00579_));
 sky130_fd_sc_hd__nand2_2 _07448_ (.A(_00578_),
    .B(_00579_),
    .Y(_00580_));
 sky130_fd_sc_hd__o22a_2 _07449_ (.A1(net104),
    .A2(net95),
    .B1(net54),
    .B2(net100),
    .X(_00581_));
 sky130_fd_sc_hd__xnor2_4 _07450_ (.A(net126),
    .B(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__xnor2_4 _07451_ (.A(_00580_),
    .B(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__or2_1 _07452_ (.A(_00573_),
    .B(_00583_),
    .X(_00584_));
 sky130_fd_sc_hd__o22a_1 _07453_ (.A1(net136),
    .A2(net65),
    .B1(net58),
    .B2(net170),
    .X(_00585_));
 sky130_fd_sc_hd__xnor2_1 _07454_ (.A(net183),
    .B(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__o22a_1 _07455_ (.A1(net107),
    .A2(net75),
    .B1(net72),
    .B2(net103),
    .X(_00587_));
 sky130_fd_sc_hd__xnor2_1 _07456_ (.A(net173),
    .B(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__nor2_1 _07457_ (.A(_00586_),
    .B(_00588_),
    .Y(_00589_));
 sky130_fd_sc_hd__and2_1 _07458_ (.A(_00586_),
    .B(_00588_),
    .X(_00590_));
 sky130_fd_sc_hd__nor2_1 _07459_ (.A(_00589_),
    .B(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__o22a_1 _07460_ (.A1(net77),
    .A2(net133),
    .B1(net62),
    .B2(net135),
    .X(_00592_));
 sky130_fd_sc_hd__xnor2_1 _07461_ (.A(net188),
    .B(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(_00591_),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__inv_2 _07463_ (.A(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__xnor2_4 _07464_ (.A(_00573_),
    .B(_00583_),
    .Y(_00596_));
 sky130_fd_sc_hd__o21ai_4 _07465_ (.A1(_00595_),
    .A2(_00596_),
    .B1(_00584_),
    .Y(_00597_));
 sky130_fd_sc_hd__o22a_1 _07466_ (.A1(net147),
    .A2(net28),
    .B1(net26),
    .B2(net174),
    .X(_00598_));
 sky130_fd_sc_hd__xnor2_1 _07467_ (.A(net68),
    .B(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__o22a_1 _07468_ (.A1(net145),
    .A2(net31),
    .B1(net30),
    .B2(net143),
    .X(_00600_));
 sky130_fd_sc_hd__xor2_1 _07469_ (.A(net118),
    .B(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__or2_1 _07470_ (.A(_00599_),
    .B(_00601_),
    .X(_00602_));
 sky130_fd_sc_hd__nand2_1 _07471_ (.A(_00599_),
    .B(_00601_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(_00602_),
    .B(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__o22a_1 _07473_ (.A1(net38),
    .A2(net141),
    .B1(net139),
    .B2(net36),
    .X(_00605_));
 sky130_fd_sc_hd__xnor2_1 _07474_ (.A(net119),
    .B(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__xnor2_1 _07475_ (.A(_00604_),
    .B(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__o21ba_1 _07476_ (.A1(_00365_),
    .A2(_00368_),
    .B1_N(_00364_),
    .X(_00608_));
 sky130_fd_sc_hd__nand2b_1 _07477_ (.A_N(_00608_),
    .B(_00460_),
    .Y(_00609_));
 sky130_fd_sc_hd__o21ai_1 _07478_ (.A1(_00399_),
    .A2(_00401_),
    .B1(_00397_),
    .Y(_00610_));
 sky130_fd_sc_hd__xnor2_1 _07479_ (.A(_00460_),
    .B(_00608_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _07480_ (.A(_00610_),
    .B(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__a21o_1 _07481_ (.A1(_00609_),
    .A2(_00612_),
    .B1(_00607_),
    .X(_00613_));
 sky130_fd_sc_hd__nand3_1 _07482_ (.A(_00607_),
    .B(_00609_),
    .C(_00612_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_2 _07483_ (.A(_00613_),
    .B(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2b_1 _07484_ (.A_N(_00615_),
    .B(_00597_),
    .Y(_00616_));
 sky130_fd_sc_hd__xnor2_4 _07485_ (.A(_00597_),
    .B(_00615_),
    .Y(_00617_));
 sky130_fd_sc_hd__o21ai_1 _07486_ (.A1(_00580_),
    .A2(_00582_),
    .B1(_00578_),
    .Y(_00618_));
 sky130_fd_sc_hd__o22a_1 _07487_ (.A1(net91),
    .A2(net48),
    .B1(net83),
    .B2(net13),
    .X(_00619_));
 sky130_fd_sc_hd__xnor2_1 _07488_ (.A(net85),
    .B(_00619_),
    .Y(_00620_));
 sky130_fd_sc_hd__o22a_1 _07489_ (.A1(net81),
    .A2(net46),
    .B1(net124),
    .B2(net11),
    .X(_00621_));
 sky130_fd_sc_hd__xnor2_1 _07490_ (.A(net111),
    .B(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__and2_1 _07491_ (.A(_00620_),
    .B(_00622_),
    .X(_00623_));
 sky130_fd_sc_hd__o21ba_1 _07492_ (.A1(_00590_),
    .A2(_00593_),
    .B1_N(_00589_),
    .X(_00624_));
 sky130_fd_sc_hd__and2b_1 _07493_ (.A_N(_00624_),
    .B(_00623_),
    .X(_00625_));
 sky130_fd_sc_hd__and2b_1 _07494_ (.A_N(_00623_),
    .B(_00624_),
    .X(_00626_));
 sky130_fd_sc_hd__nor2_1 _07495_ (.A(_00625_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__xor2_1 _07496_ (.A(_00618_),
    .B(_00627_),
    .X(_00628_));
 sky130_fd_sc_hd__o22a_1 _07497_ (.A1(net107),
    .A2(net77),
    .B1(net75),
    .B2(net103),
    .X(_00629_));
 sky130_fd_sc_hd__xnor2_2 _07498_ (.A(net173),
    .B(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__o22a_1 _07499_ (.A1(net170),
    .A2(net61),
    .B1(net58),
    .B2(net136),
    .X(_00631_));
 sky130_fd_sc_hd__xnor2_2 _07500_ (.A(net183),
    .B(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__nor2_1 _07501_ (.A(_00630_),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__xor2_2 _07502_ (.A(_00630_),
    .B(_00632_),
    .X(_00634_));
 sky130_fd_sc_hd__o22a_1 _07503_ (.A1(net135),
    .A2(net65),
    .B1(net62),
    .B2(net133),
    .X(_00635_));
 sky130_fd_sc_hd__xnor2_1 _07504_ (.A(net188),
    .B(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _07505_ (.A(_00636_),
    .Y(_00637_));
 sky130_fd_sc_hd__xnor2_1 _07506_ (.A(_00634_),
    .B(_00636_),
    .Y(_00638_));
 sky130_fd_sc_hd__o22a_1 _07507_ (.A1(net72),
    .A2(net98),
    .B1(net56),
    .B2(net69),
    .X(_00639_));
 sky130_fd_sc_hd__xnor2_1 _07508_ (.A(net129),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__o22a_1 _07509_ (.A1(net100),
    .A2(net52),
    .B1(net50),
    .B2(net57),
    .X(_00641_));
 sky130_fd_sc_hd__xnor2_1 _07510_ (.A(net89),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2b_1 _07511_ (.A_N(_00640_),
    .B(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__xor2_1 _07512_ (.A(_00640_),
    .B(_00642_),
    .X(_00644_));
 sky130_fd_sc_hd__o22a_1 _07513_ (.A1(net109),
    .A2(net95),
    .B1(net54),
    .B2(net104),
    .X(_00645_));
 sky130_fd_sc_hd__xnor2_1 _07514_ (.A(net128),
    .B(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__or2_1 _07515_ (.A(_00644_),
    .B(_00646_),
    .X(_00647_));
 sky130_fd_sc_hd__nand2_1 _07516_ (.A(_00644_),
    .B(_00646_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_00647_),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__o22a_1 _07518_ (.A1(net160),
    .A2(net20),
    .B1(net18),
    .B2(net162),
    .X(_00650_));
 sky130_fd_sc_hd__xor2_2 _07519_ (.A(net204),
    .B(_00650_),
    .X(_00651_));
 sky130_fd_sc_hd__o22a_1 _07520_ (.A1(net166),
    .A2(net24),
    .B1(net22),
    .B2(net164),
    .X(_00652_));
 sky130_fd_sc_hd__xor2_2 _07521_ (.A(net206),
    .B(_00652_),
    .X(_00653_));
 sky130_fd_sc_hd__a21oi_2 _07522_ (.A1(net299),
    .A2(net10),
    .B1(net248),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _07523_ (.A(_00653_),
    .B(_00654_),
    .Y(_00655_));
 sky130_fd_sc_hd__xor2_2 _07524_ (.A(_00653_),
    .B(_00654_),
    .X(_00656_));
 sky130_fd_sc_hd__xor2_2 _07525_ (.A(_00651_),
    .B(_00656_),
    .X(_00657_));
 sky130_fd_sc_hd__xnor2_1 _07526_ (.A(_00649_),
    .B(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__xor2_1 _07527_ (.A(_00638_),
    .B(_00658_),
    .X(_00659_));
 sky130_fd_sc_hd__or3_1 _07528_ (.A(reg1_val[29]),
    .B(reg1_val[30]),
    .C(_00219_),
    .X(_00660_));
 sky130_fd_sc_hd__a21oi_1 _07529_ (.A1(net303),
    .A2(_00660_),
    .B1(_04552_),
    .Y(_00661_));
 sky130_fd_sc_hd__a21o_1 _07530_ (.A1(net303),
    .A2(_00660_),
    .B1(_04552_),
    .X(_00662_));
 sky130_fd_sc_hd__nand2_1 _07531_ (.A(net213),
    .B(net43),
    .Y(_00663_));
 sky130_fd_sc_hd__a21oi_2 _07532_ (.A1(_00563_),
    .A2(_00572_),
    .B1(_00571_),
    .Y(_00664_));
 sky130_fd_sc_hd__a2111o_2 _07533_ (.A1(net303),
    .A2(_00219_),
    .B1(reg1_val[29]),
    .C1(reg1_val[30]),
    .D1(_04552_),
    .X(_00665_));
 sky130_fd_sc_hd__o41a_1 _07534_ (.A1(_00220_),
    .A2(_00221_),
    .A3(_00408_),
    .A4(net43),
    .B1(_00665_),
    .X(_00666_));
 sky130_fd_sc_hd__o22a_1 _07535_ (.A1(net16),
    .A2(net159),
    .B1(net7),
    .B2(net168),
    .X(_00667_));
 sky130_fd_sc_hd__xnor2_2 _07536_ (.A(net43),
    .B(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__and2b_1 _07537_ (.A_N(_00664_),
    .B(_00668_),
    .X(_00669_));
 sky130_fd_sc_hd__xnor2_2 _07538_ (.A(_00664_),
    .B(_00668_),
    .Y(_00670_));
 sky130_fd_sc_hd__xnor2_2 _07539_ (.A(_00663_),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__and2_1 _07540_ (.A(_00659_),
    .B(_00671_),
    .X(_00672_));
 sky130_fd_sc_hd__xor2_1 _07541_ (.A(_00659_),
    .B(_00671_),
    .X(_00673_));
 sky130_fd_sc_hd__xnor2_1 _07542_ (.A(_00628_),
    .B(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__o22a_1 _07543_ (.A1(net147),
    .A2(net36),
    .B1(net139),
    .B2(net38),
    .X(_00675_));
 sky130_fd_sc_hd__xnor2_1 _07544_ (.A(net121),
    .B(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__o22a_1 _07545_ (.A1(net145),
    .A2(net34),
    .B1(net122),
    .B2(net80),
    .X(_00677_));
 sky130_fd_sc_hd__xnor2_1 _07546_ (.A(net114),
    .B(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__and2_1 _07547_ (.A(_00676_),
    .B(_00678_),
    .X(_00679_));
 sky130_fd_sc_hd__nor2_1 _07548_ (.A(_00676_),
    .B(_00678_),
    .Y(_00680_));
 sky130_fd_sc_hd__nor2_1 _07549_ (.A(_00679_),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__o22a_1 _07550_ (.A1(net143),
    .A2(net31),
    .B1(net30),
    .B2(net141),
    .X(_00682_));
 sky130_fd_sc_hd__xor2_2 _07551_ (.A(net118),
    .B(_00682_),
    .X(_00683_));
 sky130_fd_sc_hd__o21bai_2 _07552_ (.A1(_00680_),
    .A2(_00683_),
    .B1_N(_00679_),
    .Y(_00684_));
 sky130_fd_sc_hd__or2_1 _07553_ (.A(net93),
    .B(net49),
    .X(_00685_));
 sky130_fd_sc_hd__a21o_1 _07554_ (.A1(_00438_),
    .A2(_00439_),
    .B1(net91),
    .X(_00686_));
 sky130_fd_sc_hd__and3_1 _07555_ (.A(net85),
    .B(_00685_),
    .C(_00686_),
    .X(_00687_));
 sky130_fd_sc_hd__a21oi_1 _07556_ (.A1(_00685_),
    .A2(_00686_),
    .B1(net85),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(_06508_),
    .B(_00450_),
    .Y(_00689_));
 sky130_fd_sc_hd__a21o_1 _07558_ (.A1(_06514_),
    .A2(_06515_),
    .B1(net122),
    .X(_00690_));
 sky130_fd_sc_hd__and3_1 _07559_ (.A(net114),
    .B(_00689_),
    .C(_00690_),
    .X(_00691_));
 sky130_fd_sc_hd__a21oi_1 _07560_ (.A1(_00689_),
    .A2(_00690_),
    .B1(net114),
    .Y(_00692_));
 sky130_fd_sc_hd__o22a_1 _07561_ (.A1(_00687_),
    .A2(_00688_),
    .B1(_00691_),
    .B2(_00692_),
    .X(_00693_));
 sky130_fd_sc_hd__or4_1 _07562_ (.A(_00687_),
    .B(_00688_),
    .C(_00691_),
    .D(_00692_),
    .X(_00694_));
 sky130_fd_sc_hd__and2b_1 _07563_ (.A_N(_00693_),
    .B(_00694_),
    .X(_00695_));
 sky130_fd_sc_hd__o22a_1 _07564_ (.A1(net83),
    .A2(net46),
    .B1(net12),
    .B2(net81),
    .X(_00696_));
 sky130_fd_sc_hd__xnor2_2 _07565_ (.A(net111),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__xor2_2 _07566_ (.A(_00695_),
    .B(_00697_),
    .X(_00698_));
 sky130_fd_sc_hd__a21oi_4 _07567_ (.A1(_00372_),
    .A2(_00381_),
    .B1(_00380_),
    .Y(_00699_));
 sky130_fd_sc_hd__o22a_2 _07568_ (.A1(net174),
    .A2(net28),
    .B1(net26),
    .B2(net159),
    .X(_00700_));
 sky130_fd_sc_hd__xor2_4 _07569_ (.A(net68),
    .B(_00700_),
    .X(_00701_));
 sky130_fd_sc_hd__and2b_1 _07570_ (.A_N(_00699_),
    .B(_00701_),
    .X(_00702_));
 sky130_fd_sc_hd__o22a_2 _07571_ (.A1(net168),
    .A2(net16),
    .B1(net7),
    .B2(net214),
    .X(_00703_));
 sky130_fd_sc_hd__xnor2_4 _07572_ (.A(net44),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__xnor2_4 _07573_ (.A(_00699_),
    .B(_00701_),
    .Y(_00705_));
 sky130_fd_sc_hd__a21o_1 _07574_ (.A1(_00704_),
    .A2(_00705_),
    .B1(_00702_),
    .X(_00706_));
 sky130_fd_sc_hd__and2_1 _07575_ (.A(_00698_),
    .B(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__xor2_1 _07576_ (.A(_00698_),
    .B(_00706_),
    .X(_00708_));
 sky130_fd_sc_hd__xnor2_1 _07577_ (.A(_00684_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__nor2_1 _07578_ (.A(_00674_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _07579_ (.A(_00674_),
    .B(_00709_),
    .Y(_00711_));
 sky130_fd_sc_hd__and2b_1 _07580_ (.A_N(_00710_),
    .B(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__xor2_4 _07581_ (.A(_00617_),
    .B(_00712_),
    .X(_00713_));
 sky130_fd_sc_hd__or2_1 _07582_ (.A(_00610_),
    .B(_00611_),
    .X(_00714_));
 sky130_fd_sc_hd__and2_2 _07583_ (.A(_00612_),
    .B(_00714_),
    .X(_00715_));
 sky130_fd_sc_hd__xnor2_4 _07584_ (.A(_00595_),
    .B(_00596_),
    .Y(_00716_));
 sky130_fd_sc_hd__xnor2_4 _07585_ (.A(_00704_),
    .B(_00705_),
    .Y(_00717_));
 sky130_fd_sc_hd__nor2_1 _07586_ (.A(_00716_),
    .B(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__xor2_4 _07587_ (.A(_00716_),
    .B(_00717_),
    .X(_00719_));
 sky130_fd_sc_hd__xor2_4 _07588_ (.A(_00715_),
    .B(_00719_),
    .X(_00720_));
 sky130_fd_sc_hd__nor2_1 _07589_ (.A(_00620_),
    .B(_00622_),
    .Y(_00721_));
 sky130_fd_sc_hd__nor2_2 _07590_ (.A(_00623_),
    .B(_00721_),
    .Y(_00722_));
 sky130_fd_sc_hd__nor2_1 _07591_ (.A(_00410_),
    .B(net44),
    .Y(_00723_));
 sky130_fd_sc_hd__a21oi_2 _07592_ (.A1(_00410_),
    .A2(_00413_),
    .B1(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__xor2_1 _07593_ (.A(_00722_),
    .B(_00724_),
    .X(_00725_));
 sky130_fd_sc_hd__o21a_1 _07594_ (.A1(_06519_),
    .A2(_00141_),
    .B1(_00725_),
    .X(_00726_));
 sky130_fd_sc_hd__nor3_1 _07595_ (.A(_06519_),
    .B(_00141_),
    .C(_00725_),
    .Y(_00727_));
 sky130_fd_sc_hd__or2_2 _07596_ (.A(_00726_),
    .B(_00727_),
    .X(_00728_));
 sky130_fd_sc_hd__inv_2 _07597_ (.A(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__a21o_2 _07598_ (.A1(_00369_),
    .A2(_00405_),
    .B1(_00403_),
    .X(_00730_));
 sky130_fd_sc_hd__xnor2_1 _07599_ (.A(_00681_),
    .B(_00683_),
    .Y(_00731_));
 sky130_fd_sc_hd__o21a_1 _07600_ (.A1(_00422_),
    .A2(_00424_),
    .B1(_00731_),
    .X(_00732_));
 sky130_fd_sc_hd__or3_1 _07601_ (.A(_00422_),
    .B(_00424_),
    .C(_00731_),
    .X(_00733_));
 sky130_fd_sc_hd__and2b_1 _07602_ (.A_N(_00732_),
    .B(_00733_),
    .X(_00734_));
 sky130_fd_sc_hd__xnor2_4 _07603_ (.A(_00730_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__xnor2_4 _07604_ (.A(_00720_),
    .B(_00728_),
    .Y(_00736_));
 sky130_fd_sc_hd__and2b_1 _07605_ (.A_N(_00735_),
    .B(_00736_),
    .X(_00737_));
 sky130_fd_sc_hd__a21oi_4 _07606_ (.A1(_00720_),
    .A2(_00729_),
    .B1(_00737_),
    .Y(_00738_));
 sky130_fd_sc_hd__a21o_2 _07607_ (.A1(_00730_),
    .A2(_00733_),
    .B1(_00732_),
    .X(_00739_));
 sky130_fd_sc_hd__a21oi_4 _07608_ (.A1(_00715_),
    .A2(_00719_),
    .B1(_00718_),
    .Y(_00740_));
 sky130_fd_sc_hd__a21oi_4 _07609_ (.A1(_00722_),
    .A2(_00724_),
    .B1(_00726_),
    .Y(_00741_));
 sky130_fd_sc_hd__nor2_1 _07610_ (.A(_00740_),
    .B(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__xor2_4 _07611_ (.A(_00740_),
    .B(_00741_),
    .X(_00743_));
 sky130_fd_sc_hd__xnor2_4 _07612_ (.A(_00739_),
    .B(_00743_),
    .Y(_00744_));
 sky130_fd_sc_hd__a21bo_2 _07613_ (.A1(_00359_),
    .A2(_00485_),
    .B1_N(_00484_),
    .X(_00745_));
 sky130_fd_sc_hd__nand2b_1 _07614_ (.A_N(_00744_),
    .B(_00745_),
    .Y(_00746_));
 sky130_fd_sc_hd__xnor2_4 _07615_ (.A(_00744_),
    .B(_00745_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand2b_1 _07616_ (.A_N(_00738_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__xnor2_4 _07617_ (.A(_00738_),
    .B(_00747_),
    .Y(_00749_));
 sky130_fd_sc_hd__and2_1 _07618_ (.A(_00713_),
    .B(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__xor2_4 _07619_ (.A(_00713_),
    .B(_00749_),
    .X(_00751_));
 sky130_fd_sc_hd__xnor2_4 _07620_ (.A(_00560_),
    .B(_00751_),
    .Y(_00752_));
 sky130_fd_sc_hd__xnor2_4 _07621_ (.A(_00735_),
    .B(_00736_),
    .Y(_00753_));
 sky130_fd_sc_hd__xnor2_2 _07622_ (.A(_00557_),
    .B(_00558_),
    .Y(_00754_));
 sky130_fd_sc_hd__and2_1 _07623_ (.A(_00753_),
    .B(_00754_),
    .X(_00755_));
 sky130_fd_sc_hd__xor2_2 _07624_ (.A(_00548_),
    .B(_00549_),
    .X(_00756_));
 sky130_fd_sc_hd__xnor2_1 _07625_ (.A(_00543_),
    .B(_00544_),
    .Y(_00757_));
 sky130_fd_sc_hd__xor2_1 _07626_ (.A(_00494_),
    .B(_00496_),
    .X(_00758_));
 sky130_fd_sc_hd__and2b_1 _07627_ (.A_N(_00757_),
    .B(_00758_),
    .X(_00759_));
 sky130_fd_sc_hd__xnor2_1 _07628_ (.A(_00757_),
    .B(_00758_),
    .Y(_00760_));
 sky130_fd_sc_hd__xor2_2 _07629_ (.A(_00521_),
    .B(_00533_),
    .X(_00761_));
 sky130_fd_sc_hd__a21oi_2 _07630_ (.A1(_00760_),
    .A2(_00761_),
    .B1(_00759_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(_00316_),
    .B(_00331_),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _07632_ (.A(_00332_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__o22a_1 _07633_ (.A1(_00392_),
    .A2(net81),
    .B1(net124),
    .B2(net51),
    .X(_00765_));
 sky130_fd_sc_hd__xnor2_1 _07634_ (.A(net90),
    .B(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__o32a_1 _07635_ (.A1(net140),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net46),
    .B2(net142),
    .X(_00767_));
 sky130_fd_sc_hd__xnor2_1 _07636_ (.A(net112),
    .B(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__xor2_1 _07637_ (.A(_00766_),
    .B(_00768_),
    .X(_00769_));
 sky130_fd_sc_hd__o22a_1 _07638_ (.A1(net144),
    .A2(net14),
    .B1(net123),
    .B2(net49),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_1 _07639_ (.A(net86),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _07640_ (.A(_00769_),
    .B(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__a21bo_1 _07641_ (.A1(_00766_),
    .A2(_00768_),
    .B1_N(_00772_),
    .X(_00773_));
 sky130_fd_sc_hd__o22a_1 _07642_ (.A1(net107),
    .A2(_00166_),
    .B1(net102),
    .B2(net101),
    .X(_00774_));
 sky130_fd_sc_hd__xnor2_1 _07643_ (.A(_00145_),
    .B(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__o22a_1 _07644_ (.A1(net96),
    .A2(net92),
    .B1(net84),
    .B2(net55),
    .X(_00776_));
 sky130_fd_sc_hd__xnor2_1 _07645_ (.A(net127),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__a22o_1 _07646_ (.A1(_00305_),
    .A2(net97),
    .B1(_00314_),
    .B2(_00323_),
    .X(_00778_));
 sky130_fd_sc_hd__xor2_1 _07647_ (.A(net131),
    .B(_00778_),
    .X(_00779_));
 sky130_fd_sc_hd__xnor2_1 _07648_ (.A(_00775_),
    .B(_00777_),
    .Y(_00780_));
 sky130_fd_sc_hd__or2_1 _07649_ (.A(_00779_),
    .B(_00780_),
    .X(_00781_));
 sky130_fd_sc_hd__o21ai_1 _07650_ (.A1(_00775_),
    .A2(_00777_),
    .B1(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__xor2_1 _07651_ (.A(_00764_),
    .B(_00773_),
    .X(_00783_));
 sky130_fd_sc_hd__and2b_1 _07652_ (.A_N(_00783_),
    .B(_00782_),
    .X(_00784_));
 sky130_fd_sc_hd__a31oi_4 _07653_ (.A1(_00332_),
    .A2(_00763_),
    .A3(_00773_),
    .B1(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__nor2_1 _07654_ (.A(_00762_),
    .B(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hd__xor2_1 _07655_ (.A(_00504_),
    .B(_00506_),
    .X(_00787_));
 sky130_fd_sc_hd__o22a_1 _07656_ (.A1(net214),
    .A2(net36),
    .B1(net168),
    .B2(net38),
    .X(_00788_));
 sky130_fd_sc_hd__xnor2_1 _07657_ (.A(net121),
    .B(_00788_),
    .Y(_00789_));
 sky130_fd_sc_hd__o22a_1 _07658_ (.A1(net147),
    .A2(net34),
    .B1(net138),
    .B2(net80),
    .X(_00790_));
 sky130_fd_sc_hd__xnor2_1 _07659_ (.A(net115),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__and2_1 _07660_ (.A(_00789_),
    .B(_00791_),
    .X(_00792_));
 sky130_fd_sc_hd__nor2_1 _07661_ (.A(_00789_),
    .B(_00791_),
    .Y(_00793_));
 sky130_fd_sc_hd__nor2_1 _07662_ (.A(_00792_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__o22a_1 _07663_ (.A1(net174),
    .A2(net31),
    .B1(net30),
    .B2(net159),
    .X(_00795_));
 sky130_fd_sc_hd__xnor2_1 _07664_ (.A(net118),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__and2_1 _07665_ (.A(_00794_),
    .B(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__o21ai_1 _07666_ (.A1(_00792_),
    .A2(_00797_),
    .B1(_00787_),
    .Y(_00798_));
 sky130_fd_sc_hd__a21o_1 _07667_ (.A1(_00528_),
    .A2(_00531_),
    .B1(_00530_),
    .X(_00799_));
 sky130_fd_sc_hd__o22a_1 _07668_ (.A1(net77),
    .A2(net166),
    .B1(net164),
    .B2(net76),
    .X(_00800_));
 sky130_fd_sc_hd__xnor2_2 _07669_ (.A(net207),
    .B(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__o22a_1 _07670_ (.A1(net299),
    .A2(net61),
    .B1(_00289_),
    .B2(net247),
    .X(_00802_));
 sky130_fd_sc_hd__xnor2_1 _07671_ (.A(net248),
    .B(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_1 _07672_ (.A(_00801_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hd__o22a_1 _07673_ (.A1(net65),
    .A2(net162),
    .B1(net160),
    .B2(_00251_),
    .X(_00805_));
 sky130_fd_sc_hd__xor2_2 _07674_ (.A(net204),
    .B(_00805_),
    .X(_00806_));
 sky130_fd_sc_hd__nand2_1 _07675_ (.A(_00801_),
    .B(_00803_),
    .Y(_00807_));
 sky130_fd_sc_hd__xnor2_1 _07676_ (.A(_00801_),
    .B(_00803_),
    .Y(_00808_));
 sky130_fd_sc_hd__a21o_1 _07677_ (.A1(_00806_),
    .A2(_00807_),
    .B1(_00804_),
    .X(_00809_));
 sky130_fd_sc_hd__nand3_2 _07678_ (.A(_00532_),
    .B(_00799_),
    .C(_00809_),
    .Y(_00810_));
 sky130_fd_sc_hd__o22a_1 _07679_ (.A1(net171),
    .A2(net73),
    .B1(net69),
    .B2(net136),
    .X(_00811_));
 sky130_fd_sc_hd__xnor2_1 _07680_ (.A(_00171_),
    .B(_00811_),
    .Y(_00812_));
 sky130_fd_sc_hd__o22a_1 _07681_ (.A1(_00155_),
    .A2(net135),
    .B1(net133),
    .B2(_00166_),
    .X(_00813_));
 sky130_fd_sc_hd__xnor2_1 _07682_ (.A(net188),
    .B(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__nor2_1 _07683_ (.A(_00812_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__a21o_1 _07684_ (.A1(_00532_),
    .A2(_00799_),
    .B1(_00809_),
    .X(_00816_));
 sky130_fd_sc_hd__nand3_2 _07685_ (.A(_00810_),
    .B(_00815_),
    .C(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_2 _07686_ (.A(_00810_),
    .B(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__or3_1 _07687_ (.A(_00787_),
    .B(_00792_),
    .C(_00797_),
    .X(_00819_));
 sky130_fd_sc_hd__and2_1 _07688_ (.A(_00798_),
    .B(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__a21bo_1 _07689_ (.A1(_00818_),
    .A2(_00819_),
    .B1_N(_00798_),
    .X(_00821_));
 sky130_fd_sc_hd__xor2_2 _07690_ (.A(_00762_),
    .B(_00785_),
    .X(_00822_));
 sky130_fd_sc_hd__a21oi_2 _07691_ (.A1(_00821_),
    .A2(_00822_),
    .B1(_00786_),
    .Y(_00823_));
 sky130_fd_sc_hd__and2b_1 _07692_ (.A_N(_00507_),
    .B(_00508_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _07693_ (.A(_00509_),
    .B(_00824_),
    .X(_00825_));
 sky130_fd_sc_hd__xnor2_1 _07694_ (.A(_00516_),
    .B(_00517_),
    .Y(_00826_));
 sky130_fd_sc_hd__nor2_1 _07695_ (.A(_00825_),
    .B(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__xnor2_4 _07696_ (.A(_00545_),
    .B(_00546_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(_00825_),
    .B(_00826_),
    .Y(_00829_));
 sky130_fd_sc_hd__and2b_1 _07698_ (.A_N(_00827_),
    .B(_00829_),
    .X(_00830_));
 sky130_fd_sc_hd__a21o_1 _07699_ (.A1(_00828_),
    .A2(_00829_),
    .B1(_00827_),
    .X(_00831_));
 sky130_fd_sc_hd__xnor2_1 _07700_ (.A(_00756_),
    .B(_00823_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2b_1 _07701_ (.A_N(_00832_),
    .B(_00831_),
    .Y(_00833_));
 sky130_fd_sc_hd__o21ai_4 _07702_ (.A1(_00756_),
    .A2(_00823_),
    .B1(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__xor2_4 _07703_ (.A(_00753_),
    .B(_00754_),
    .X(_00835_));
 sky130_fd_sc_hd__a21oi_4 _07704_ (.A1(_00834_),
    .A2(_00835_),
    .B1(_00755_),
    .Y(_00836_));
 sky130_fd_sc_hd__or2_1 _07705_ (.A(_00752_),
    .B(_00836_),
    .X(_00837_));
 sky130_fd_sc_hd__and2_1 _07706_ (.A(_00752_),
    .B(_00836_),
    .X(_00838_));
 sky130_fd_sc_hd__xnor2_4 _07707_ (.A(_00752_),
    .B(_00836_),
    .Y(_00839_));
 sky130_fd_sc_hd__or2_1 _07708_ (.A(net146),
    .B(net49),
    .X(_00840_));
 sky130_fd_sc_hd__a21o_1 _07709_ (.A1(_00438_),
    .A2(_00439_),
    .B1(net175),
    .X(_00841_));
 sky130_fd_sc_hd__nand3_1 _07710_ (.A(net86),
    .B(_00840_),
    .C(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__a21o_1 _07711_ (.A1(_00840_),
    .A2(_00841_),
    .B1(net86),
    .X(_00843_));
 sky130_fd_sc_hd__o32a_1 _07712_ (.A1(net169),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net158),
    .B2(net46),
    .X(_00844_));
 sky130_fd_sc_hd__xnor2_1 _07713_ (.A(_06505_),
    .B(_00844_),
    .Y(_00845_));
 sky130_fd_sc_hd__a21o_1 _07714_ (.A1(_00842_),
    .A2(_00843_),
    .B1(_00845_),
    .X(_00846_));
 sky130_fd_sc_hd__inv_2 _07715_ (.A(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__nand3_1 _07716_ (.A(_00842_),
    .B(_00843_),
    .C(_00845_),
    .Y(_00848_));
 sky130_fd_sc_hd__o22a_1 _07717_ (.A1(net106),
    .A2(net84),
    .B1(net81),
    .B2(net102),
    .X(_00849_));
 sky130_fd_sc_hd__xnor2_2 _07718_ (.A(net172),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__a22o_1 _07719_ (.A1(_00180_),
    .A2(net99),
    .B1(net97),
    .B2(_00190_),
    .X(_00851_));
 sky130_fd_sc_hd__xor2_2 _07720_ (.A(net185),
    .B(_00851_),
    .X(_00852_));
 sky130_fd_sc_hd__nor2_1 _07721_ (.A(_00850_),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__xor2_2 _07722_ (.A(_00850_),
    .B(_00852_),
    .X(_00854_));
 sky130_fd_sc_hd__o22a_1 _07723_ (.A1(_00205_),
    .A2(net94),
    .B1(net92),
    .B2(net133),
    .X(_00855_));
 sky130_fd_sc_hd__xnor2_1 _07724_ (.A(net187),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__inv_2 _07725_ (.A(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__xnor2_1 _07726_ (.A(_00854_),
    .B(_00856_),
    .Y(_00858_));
 sky130_fd_sc_hd__and3_1 _07727_ (.A(_00846_),
    .B(_00848_),
    .C(_00858_),
    .X(_00859_));
 sky130_fd_sc_hd__a21oi_1 _07728_ (.A1(_00846_),
    .A2(_00848_),
    .B1(_00858_),
    .Y(_00860_));
 sky130_fd_sc_hd__a22o_1 _07729_ (.A1(_00305_),
    .A2(_00450_),
    .B1(_00457_),
    .B2(_00314_),
    .X(_00861_));
 sky130_fd_sc_hd__xor2_1 _07730_ (.A(net131),
    .B(_00861_),
    .X(_00862_));
 sky130_fd_sc_hd__o22a_1 _07731_ (.A1(net140),
    .A2(net53),
    .B1(net51),
    .B2(net139),
    .X(_00863_));
 sky130_fd_sc_hd__xnor2_1 _07732_ (.A(_00388_),
    .B(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__or2_1 _07733_ (.A(_00862_),
    .B(_00864_),
    .X(_00865_));
 sky130_fd_sc_hd__xnor2_1 _07734_ (.A(_00862_),
    .B(_00864_),
    .Y(_00866_));
 sky130_fd_sc_hd__o22a_1 _07735_ (.A1(net144),
    .A2(net96),
    .B1(net55),
    .B2(net142),
    .X(_00867_));
 sky130_fd_sc_hd__xnor2_1 _07736_ (.A(net127),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__xnor2_1 _07737_ (.A(_00866_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__or3_1 _07738_ (.A(_00859_),
    .B(_00860_),
    .C(_00869_),
    .X(_00870_));
 sky130_fd_sc_hd__o21ai_1 _07739_ (.A1(_00859_),
    .A2(_00860_),
    .B1(_00869_),
    .Y(_00871_));
 sky130_fd_sc_hd__nor2_1 _07740_ (.A(net215),
    .B(net79),
    .Y(_00872_));
 sky130_fd_sc_hd__a21oi_1 _07741_ (.A1(_00192_),
    .A2(_00193_),
    .B1(net300),
    .Y(_00873_));
 sky130_fd_sc_hd__and3_1 _07742_ (.A(_00199_),
    .B(_00200_),
    .C(_00265_),
    .X(_00874_));
 sky130_fd_sc_hd__o21ai_1 _07743_ (.A1(_00873_),
    .A2(_00874_),
    .B1(net250),
    .Y(_00875_));
 sky130_fd_sc_hd__or3_1 _07744_ (.A(net250),
    .B(_00873_),
    .C(_00874_),
    .X(_00876_));
 sky130_fd_sc_hd__o22a_1 _07745_ (.A1(net105),
    .A2(net167),
    .B1(net165),
    .B2(net101),
    .X(_00877_));
 sky130_fd_sc_hd__xor2_1 _07746_ (.A(net208),
    .B(_00877_),
    .X(_00878_));
 sky130_fd_sc_hd__and3_1 _07747_ (.A(_00875_),
    .B(_00876_),
    .C(_00878_),
    .X(_00879_));
 sky130_fd_sc_hd__o22a_1 _07748_ (.A1(net70),
    .A2(net163),
    .B1(net161),
    .B2(net109),
    .X(_00880_));
 sky130_fd_sc_hd__xor2_1 _07749_ (.A(net205),
    .B(_00880_),
    .X(_00881_));
 sky130_fd_sc_hd__a21oi_1 _07750_ (.A1(_00875_),
    .A2(_00876_),
    .B1(_00878_),
    .Y(_00882_));
 sky130_fd_sc_hd__or3b_1 _07751_ (.A(_00879_),
    .B(_00882_),
    .C_N(_00881_),
    .X(_00883_));
 sky130_fd_sc_hd__and2b_1 _07752_ (.A_N(_00879_),
    .B(_00883_),
    .X(_00884_));
 sky130_fd_sc_hd__xnor2_1 _07753_ (.A(_00872_),
    .B(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__and3_1 _07754_ (.A(_00870_),
    .B(_00871_),
    .C(_00885_),
    .X(_00886_));
 sky130_fd_sc_hd__a21oi_1 _07755_ (.A1(_00870_),
    .A2(_00871_),
    .B1(_00885_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_2 _07756_ (.A(_00886_),
    .B(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__a22o_1 _07757_ (.A1(_06502_),
    .A2(_00314_),
    .B1(_00457_),
    .B2(_00305_),
    .X(_00889_));
 sky130_fd_sc_hd__xor2_2 _07758_ (.A(net131),
    .B(_00889_),
    .X(_00890_));
 sky130_fd_sc_hd__o22a_1 _07759_ (.A1(net142),
    .A2(net96),
    .B1(net55),
    .B2(net140),
    .X(_00891_));
 sky130_fd_sc_hd__xnor2_2 _07760_ (.A(net127),
    .B(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__or2_2 _07761_ (.A(_00890_),
    .B(_00892_),
    .X(_00893_));
 sky130_fd_sc_hd__o22a_2 _07762_ (.A1(_00155_),
    .A2(net167),
    .B1(net165),
    .B2(net105),
    .X(_00894_));
 sky130_fd_sc_hd__xnor2_4 _07763_ (.A(_00173_),
    .B(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__o22a_2 _07764_ (.A1(net300),
    .A2(net77),
    .B1(net76),
    .B2(_00266_),
    .X(_00896_));
 sky130_fd_sc_hd__xnor2_4 _07765_ (.A(net249),
    .B(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__nor2_1 _07766_ (.A(_00895_),
    .B(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__xor2_4 _07767_ (.A(_00895_),
    .B(_00897_),
    .X(_00899_));
 sky130_fd_sc_hd__o22a_2 _07768_ (.A1(net73),
    .A2(net163),
    .B1(net161),
    .B2(net70),
    .X(_00900_));
 sky130_fd_sc_hd__xor2_4 _07769_ (.A(net205),
    .B(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__xnor2_4 _07770_ (.A(_00899_),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__o22a_1 _07771_ (.A1(net106),
    .A2(net82),
    .B1(net124),
    .B2(net102),
    .X(_00903_));
 sky130_fd_sc_hd__xnor2_1 _07772_ (.A(net172),
    .B(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__a22o_1 _07773_ (.A1(_00180_),
    .A2(net97),
    .B1(_00323_),
    .B2(_00190_),
    .X(_00905_));
 sky130_fd_sc_hd__xor2_1 _07774_ (.A(_00171_),
    .B(_00905_),
    .X(_00906_));
 sky130_fd_sc_hd__xor2_1 _07775_ (.A(_00904_),
    .B(_00906_),
    .X(_00907_));
 sky130_fd_sc_hd__o22a_1 _07776_ (.A1(net134),
    .A2(net92),
    .B1(net84),
    .B2(net132),
    .X(_00908_));
 sky130_fd_sc_hd__xnor2_1 _07777_ (.A(net188),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__and2b_1 _07778_ (.A_N(_00909_),
    .B(_00907_),
    .X(_00910_));
 sky130_fd_sc_hd__o21ba_2 _07779_ (.A1(_00904_),
    .A2(_00906_),
    .B1_N(_00910_),
    .X(_00911_));
 sky130_fd_sc_hd__xnor2_4 _07780_ (.A(_00902_),
    .B(_00911_),
    .Y(_00912_));
 sky130_fd_sc_hd__xnor2_4 _07781_ (.A(_00893_),
    .B(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_4 _07782_ (.A(_00888_),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hd__xor2_1 _07783_ (.A(_00890_),
    .B(_00892_),
    .X(_00915_));
 sky130_fd_sc_hd__o21bai_1 _07784_ (.A1(_00879_),
    .A2(_00882_),
    .B1_N(_00881_),
    .Y(_00916_));
 sky130_fd_sc_hd__and3_1 _07785_ (.A(_00883_),
    .B(_00915_),
    .C(_00916_),
    .X(_00917_));
 sky130_fd_sc_hd__inv_2 _07786_ (.A(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hd__a21oi_1 _07787_ (.A1(_00883_),
    .A2(_00916_),
    .B1(_00915_),
    .Y(_00919_));
 sky130_fd_sc_hd__and2b_1 _07788_ (.A_N(_00907_),
    .B(_00909_),
    .X(_00920_));
 sky130_fd_sc_hd__or2_1 _07789_ (.A(_00910_),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__or3_1 _07790_ (.A(_00917_),
    .B(_00919_),
    .C(_00921_),
    .X(_00922_));
 sky130_fd_sc_hd__o21ai_1 _07791_ (.A1(_00917_),
    .A2(_00919_),
    .B1(_00921_),
    .Y(_00923_));
 sky130_fd_sc_hd__o22a_1 _07792_ (.A1(net138),
    .A2(net53),
    .B1(net51),
    .B2(net146),
    .X(_00924_));
 sky130_fd_sc_hd__xnor2_1 _07793_ (.A(net90),
    .B(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hd__o32a_1 _07794_ (.A1(net215),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net169),
    .B2(net47),
    .X(_00926_));
 sky130_fd_sc_hd__xnor2_1 _07795_ (.A(net112),
    .B(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__and2_1 _07796_ (.A(_00925_),
    .B(_00927_),
    .X(_00928_));
 sky130_fd_sc_hd__nor2_1 _07797_ (.A(_00925_),
    .B(_00927_),
    .Y(_00929_));
 sky130_fd_sc_hd__nor2_1 _07798_ (.A(_00928_),
    .B(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__o22a_1 _07799_ (.A1(net175),
    .A2(net49),
    .B1(net14),
    .B2(net158),
    .X(_00931_));
 sky130_fd_sc_hd__xnor2_1 _07800_ (.A(net86),
    .B(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__xor2_1 _07801_ (.A(_00930_),
    .B(_00932_),
    .X(_00933_));
 sky130_fd_sc_hd__and3_1 _07802_ (.A(_00922_),
    .B(_00923_),
    .C(_00933_),
    .X(_00934_));
 sky130_fd_sc_hd__a21oi_1 _07803_ (.A1(_00922_),
    .A2(_00923_),
    .B1(_00933_),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_2 _07804_ (.A(_00934_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__o22a_1 _07805_ (.A1(net106),
    .A2(net124),
    .B1(net123),
    .B2(net102),
    .X(_00937_));
 sky130_fd_sc_hd__xnor2_2 _07806_ (.A(net172),
    .B(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__o22a_1 _07807_ (.A1(net171),
    .A2(net94),
    .B1(net92),
    .B2(net137),
    .X(_00939_));
 sky130_fd_sc_hd__xnor2_2 _07808_ (.A(net185),
    .B(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__xor2_1 _07809_ (.A(_00938_),
    .B(_00940_),
    .X(_00941_));
 sky130_fd_sc_hd__o22a_1 _07810_ (.A1(net134),
    .A2(net84),
    .B1(net82),
    .B2(net132),
    .X(_00942_));
 sky130_fd_sc_hd__xnor2_1 _07811_ (.A(net187),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__and2b_1 _07812_ (.A_N(_00943_),
    .B(_00941_),
    .X(_00944_));
 sky130_fd_sc_hd__o21bai_4 _07813_ (.A1(_00938_),
    .A2(_00940_),
    .B1_N(_00944_),
    .Y(_00945_));
 sky130_fd_sc_hd__a22o_2 _07814_ (.A1(_06502_),
    .A2(_00305_),
    .B1(_00314_),
    .B2(_06513_),
    .X(_00946_));
 sky130_fd_sc_hd__xor2_4 _07815_ (.A(net130),
    .B(_00946_),
    .X(_00947_));
 sky130_fd_sc_hd__o22a_2 _07816_ (.A1(net140),
    .A2(net96),
    .B1(net55),
    .B2(net138),
    .X(_00948_));
 sky130_fd_sc_hd__xnor2_4 _07817_ (.A(net127),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__nor2_2 _07818_ (.A(_00947_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__a22o_1 _07819_ (.A1(_00241_),
    .A2(_00300_),
    .B1(_00310_),
    .B2(_00249_),
    .X(_00951_));
 sky130_fd_sc_hd__xnor2_1 _07820_ (.A(net208),
    .B(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__and3_1 _07821_ (.A(net302),
    .B(_00199_),
    .C(_00200_),
    .X(_00953_));
 sky130_fd_sc_hd__a21oi_1 _07822_ (.A1(_00208_),
    .A2(_00209_),
    .B1(net247),
    .Y(_00954_));
 sky130_fd_sc_hd__o21ai_1 _07823_ (.A1(_00953_),
    .A2(_00954_),
    .B1(net250),
    .Y(_00955_));
 sky130_fd_sc_hd__or3_1 _07824_ (.A(net250),
    .B(_00953_),
    .C(_00954_),
    .X(_00956_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_00952_),
    .B(_00955_),
    .C(_00956_),
    .Y(_00957_));
 sky130_fd_sc_hd__o22a_1 _07826_ (.A1(net109),
    .A2(net163),
    .B1(net161),
    .B2(net105),
    .X(_00958_));
 sky130_fd_sc_hd__xor2_2 _07827_ (.A(net205),
    .B(_00958_),
    .X(_00959_));
 sky130_fd_sc_hd__a21o_1 _07828_ (.A1(_00955_),
    .A2(_00956_),
    .B1(_00952_),
    .X(_00960_));
 sky130_fd_sc_hd__nand3_1 _07829_ (.A(_00957_),
    .B(_00959_),
    .C(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hd__a21boi_4 _07830_ (.A1(_00959_),
    .A2(_00960_),
    .B1_N(_00957_),
    .Y(_00962_));
 sky130_fd_sc_hd__xnor2_4 _07831_ (.A(_00950_),
    .B(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _07832_ (.A(_00945_),
    .B(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__xnor2_4 _07833_ (.A(_00945_),
    .B(_00963_),
    .Y(_00965_));
 sky130_fd_sc_hd__o21ba_2 _07834_ (.A1(_00935_),
    .A2(_00965_),
    .B1_N(_00934_),
    .X(_00966_));
 sky130_fd_sc_hd__o31ai_4 _07835_ (.A1(_00947_),
    .A2(_00949_),
    .A3(_00962_),
    .B1(_00964_),
    .Y(_00967_));
 sky130_fd_sc_hd__o21bai_2 _07836_ (.A1(_00919_),
    .A2(_00921_),
    .B1_N(_00917_),
    .Y(_00968_));
 sky130_fd_sc_hd__a21oi_2 _07837_ (.A1(_00930_),
    .A2(_00932_),
    .B1(_00928_),
    .Y(_00969_));
 sky130_fd_sc_hd__a21o_1 _07838_ (.A1(_00918_),
    .A2(_00922_),
    .B1(_00969_),
    .X(_00970_));
 sky130_fd_sc_hd__nand2b_1 _07839_ (.A_N(_00968_),
    .B(_00969_),
    .Y(_00971_));
 sky130_fd_sc_hd__xor2_2 _07840_ (.A(_00968_),
    .B(_00969_),
    .X(_00972_));
 sky130_fd_sc_hd__xnor2_4 _07841_ (.A(_00967_),
    .B(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__xor2_2 _07842_ (.A(_00947_),
    .B(_00949_),
    .X(_00974_));
 sky130_fd_sc_hd__a21o_1 _07843_ (.A1(_00957_),
    .A2(_00960_),
    .B1(_00959_),
    .X(_00975_));
 sky130_fd_sc_hd__and3_1 _07844_ (.A(_00961_),
    .B(_00974_),
    .C(_00975_),
    .X(_00976_));
 sky130_fd_sc_hd__a21oi_2 _07845_ (.A1(_00961_),
    .A2(_00975_),
    .B1(_00974_),
    .Y(_00977_));
 sky130_fd_sc_hd__and2b_1 _07846_ (.A_N(_00941_),
    .B(_00943_),
    .X(_00978_));
 sky130_fd_sc_hd__or2_1 _07847_ (.A(_00944_),
    .B(_00978_),
    .X(_00979_));
 sky130_fd_sc_hd__or3_1 _07848_ (.A(_00976_),
    .B(_00977_),
    .C(_00979_),
    .X(_00980_));
 sky130_fd_sc_hd__o21ba_2 _07849_ (.A1(_00977_),
    .A2(_00979_),
    .B1_N(_00976_),
    .X(_00981_));
 sky130_fd_sc_hd__o22a_1 _07850_ (.A1(net146),
    .A2(net53),
    .B1(net51),
    .B2(net174),
    .X(_00982_));
 sky130_fd_sc_hd__xnor2_1 _07851_ (.A(net90),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__nor2_1 _07852_ (.A(net215),
    .B(_00449_),
    .Y(_00984_));
 sky130_fd_sc_hd__xnor2_2 _07853_ (.A(net111),
    .B(_00984_),
    .Y(_00985_));
 sky130_fd_sc_hd__and2b_1 _07854_ (.A_N(_00985_),
    .B(_00983_),
    .X(_00986_));
 sky130_fd_sc_hd__xor2_1 _07855_ (.A(_00983_),
    .B(_00985_),
    .X(_00987_));
 sky130_fd_sc_hd__inv_2 _07856_ (.A(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__o22a_1 _07857_ (.A1(net158),
    .A2(net49),
    .B1(net14),
    .B2(net169),
    .X(_00989_));
 sky130_fd_sc_hd__xnor2_2 _07858_ (.A(net86),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__a21oi_2 _07859_ (.A1(_00988_),
    .A2(_00990_),
    .B1(_00986_),
    .Y(_00991_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(_00981_),
    .B(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__o22a_1 _07861_ (.A1(net171),
    .A2(net92),
    .B1(net84),
    .B2(net137),
    .X(_00993_));
 sky130_fd_sc_hd__xnor2_1 _07862_ (.A(net185),
    .B(_00993_),
    .Y(_00994_));
 sky130_fd_sc_hd__o22a_1 _07863_ (.A1(net134),
    .A2(net82),
    .B1(net125),
    .B2(net132),
    .X(_00995_));
 sky130_fd_sc_hd__xnor2_1 _07864_ (.A(net187),
    .B(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__or2_2 _07865_ (.A(_00994_),
    .B(_00996_),
    .X(_00997_));
 sky130_fd_sc_hd__a22o_1 _07866_ (.A1(_00241_),
    .A2(_00310_),
    .B1(_00323_),
    .B2(_00249_),
    .X(_00998_));
 sky130_fd_sc_hd__xor2_1 _07867_ (.A(net208),
    .B(_00998_),
    .X(_00999_));
 sky130_fd_sc_hd__a21o_1 _07868_ (.A1(_00208_),
    .A2(_00209_),
    .B1(net300),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _07869_ (.A(net109),
    .B(_00266_),
    .X(_01001_));
 sky130_fd_sc_hd__a21oi_1 _07870_ (.A1(_01000_),
    .A2(_01001_),
    .B1(_00256_),
    .Y(_01002_));
 sky130_fd_sc_hd__and3_1 _07871_ (.A(net249),
    .B(_01000_),
    .C(_01001_),
    .X(_01003_));
 sky130_fd_sc_hd__or3_2 _07872_ (.A(_00999_),
    .B(_01002_),
    .C(_01003_),
    .X(_01004_));
 sky130_fd_sc_hd__o22a_1 _07873_ (.A1(net105),
    .A2(net163),
    .B1(net161),
    .B2(net101),
    .X(_01005_));
 sky130_fd_sc_hd__xnor2_1 _07874_ (.A(net205),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__o21ai_1 _07875_ (.A1(_01002_),
    .A2(_01003_),
    .B1(_00999_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand3b_2 _07876_ (.A_N(_01006_),
    .B(_01007_),
    .C(_01004_),
    .Y(_01008_));
 sky130_fd_sc_hd__xnor2_1 _07877_ (.A(_06505_),
    .B(_00997_),
    .Y(_01009_));
 sky130_fd_sc_hd__a21o_1 _07878_ (.A1(_01004_),
    .A2(_01008_),
    .B1(_01009_),
    .X(_01010_));
 sky130_fd_sc_hd__o21ai_4 _07879_ (.A1(_06505_),
    .A2(_00997_),
    .B1(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__xor2_4 _07880_ (.A(_00981_),
    .B(_00991_),
    .X(_01012_));
 sky130_fd_sc_hd__a21oi_4 _07881_ (.A1(_01011_),
    .A2(_01012_),
    .B1(_00992_),
    .Y(_01013_));
 sky130_fd_sc_hd__and2b_1 _07882_ (.A_N(_01013_),
    .B(_00973_),
    .X(_01014_));
 sky130_fd_sc_hd__xnor2_4 _07883_ (.A(_00973_),
    .B(_01013_),
    .Y(_01015_));
 sky130_fd_sc_hd__and2b_1 _07884_ (.A_N(_00966_),
    .B(_01015_),
    .X(_01016_));
 sky130_fd_sc_hd__xnor2_4 _07885_ (.A(_00966_),
    .B(_01015_),
    .Y(_01017_));
 sky130_fd_sc_hd__and2_1 _07886_ (.A(_00914_),
    .B(_01017_),
    .X(_01018_));
 sky130_fd_sc_hd__xor2_4 _07887_ (.A(_00914_),
    .B(_01017_),
    .X(_01019_));
 sky130_fd_sc_hd__xnor2_2 _07888_ (.A(_01011_),
    .B(_01012_),
    .Y(_01020_));
 sky130_fd_sc_hd__o22a_1 _07889_ (.A1(net144),
    .A2(net102),
    .B1(net123),
    .B2(net106),
    .X(_01021_));
 sky130_fd_sc_hd__nor2_1 _07890_ (.A(net172),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__and2_1 _07891_ (.A(net172),
    .B(_01021_),
    .X(_01023_));
 sky130_fd_sc_hd__or2_1 _07892_ (.A(_01022_),
    .B(_01023_),
    .X(_01024_));
 sky130_fd_sc_hd__o22a_1 _07893_ (.A1(_00136_),
    .A2(net96),
    .B1(net55),
    .B2(net146),
    .X(_01025_));
 sky130_fd_sc_hd__xnor2_1 _07894_ (.A(_00320_),
    .B(_01025_),
    .Y(_01026_));
 sky130_fd_sc_hd__a22o_1 _07895_ (.A1(_06513_),
    .A2(_00305_),
    .B1(_00314_),
    .B2(_06522_),
    .X(_01027_));
 sky130_fd_sc_hd__xor2_1 _07896_ (.A(net130),
    .B(_01027_),
    .X(_01028_));
 sky130_fd_sc_hd__xnor2_1 _07897_ (.A(_01024_),
    .B(_01026_),
    .Y(_01029_));
 sky130_fd_sc_hd__o32a_1 _07898_ (.A1(_01022_),
    .A2(_01023_),
    .A3(_01026_),
    .B1(_01028_),
    .B2(_01029_),
    .X(_01030_));
 sky130_fd_sc_hd__o22a_1 _07899_ (.A1(net171),
    .A2(net84),
    .B1(net82),
    .B2(net137),
    .X(_01031_));
 sky130_fd_sc_hd__xnor2_2 _07900_ (.A(net185),
    .B(_01031_),
    .Y(_01032_));
 sky130_fd_sc_hd__o22a_1 _07901_ (.A1(net134),
    .A2(net125),
    .B1(net122),
    .B2(net132),
    .X(_01033_));
 sky130_fd_sc_hd__xnor2_2 _07902_ (.A(net188),
    .B(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__or2_1 _07903_ (.A(_01032_),
    .B(_01034_),
    .X(_01035_));
 sky130_fd_sc_hd__xnor2_1 _07904_ (.A(_00994_),
    .B(_00996_),
    .Y(_01036_));
 sky130_fd_sc_hd__nor2_1 _07905_ (.A(_01035_),
    .B(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__a21bo_1 _07906_ (.A1(_01004_),
    .A2(_01007_),
    .B1_N(_01006_),
    .X(_01038_));
 sky130_fd_sc_hd__xor2_1 _07907_ (.A(_01035_),
    .B(_01036_),
    .X(_01039_));
 sky130_fd_sc_hd__and3_1 _07908_ (.A(_01008_),
    .B(_01038_),
    .C(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__a31o_1 _07909_ (.A1(_01008_),
    .A2(_01038_),
    .A3(_01039_),
    .B1(_01037_),
    .X(_01041_));
 sky130_fd_sc_hd__nand2b_1 _07910_ (.A_N(_01030_),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__o22a_1 _07911_ (.A1(net300),
    .A2(net109),
    .B1(net105),
    .B2(_00266_),
    .X(_01043_));
 sky130_fd_sc_hd__xnor2_2 _07912_ (.A(net249),
    .B(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__o22a_1 _07913_ (.A1(net167),
    .A2(net94),
    .B1(net92),
    .B2(net165),
    .X(_01045_));
 sky130_fd_sc_hd__xnor2_2 _07914_ (.A(net208),
    .B(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__nor2_1 _07915_ (.A(_01044_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__a22o_1 _07916_ (.A1(_00281_),
    .A2(_00300_),
    .B1(net97),
    .B2(_00287_),
    .X(_01048_));
 sky130_fd_sc_hd__xor2_2 _07917_ (.A(net205),
    .B(_01048_),
    .X(_01049_));
 sky130_fd_sc_hd__inv_2 _07918_ (.A(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__xor2_2 _07919_ (.A(_01044_),
    .B(_01046_),
    .X(_01051_));
 sky130_fd_sc_hd__a21oi_1 _07920_ (.A1(_01050_),
    .A2(_01051_),
    .B1(_01047_),
    .Y(_01052_));
 sky130_fd_sc_hd__o22a_1 _07921_ (.A1(net175),
    .A2(net53),
    .B1(net51),
    .B2(net158),
    .X(_01053_));
 sky130_fd_sc_hd__xnor2_1 _07922_ (.A(net90),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2b_1 _07923_ (.A_N(_01052_),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__xnor2_1 _07924_ (.A(_01052_),
    .B(_01054_),
    .Y(_01056_));
 sky130_fd_sc_hd__o22a_1 _07925_ (.A1(net169),
    .A2(net49),
    .B1(net14),
    .B2(net215),
    .X(_01057_));
 sky130_fd_sc_hd__xnor2_1 _07926_ (.A(net87),
    .B(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__a21boi_2 _07927_ (.A1(_01056_),
    .A2(_01058_),
    .B1_N(_01055_),
    .Y(_01059_));
 sky130_fd_sc_hd__xor2_2 _07928_ (.A(_01030_),
    .B(_01041_),
    .X(_01060_));
 sky130_fd_sc_hd__o21ai_2 _07929_ (.A1(_01059_),
    .A2(_01060_),
    .B1(_01042_),
    .Y(_01061_));
 sky130_fd_sc_hd__and2b_1 _07930_ (.A_N(_01020_),
    .B(_01061_),
    .X(_01062_));
 sky130_fd_sc_hd__o21ai_1 _07931_ (.A1(_00976_),
    .A2(_00977_),
    .B1(_00979_),
    .Y(_01063_));
 sky130_fd_sc_hd__xnor2_1 _07932_ (.A(_00987_),
    .B(_00990_),
    .Y(_01064_));
 sky130_fd_sc_hd__and3_1 _07933_ (.A(_00980_),
    .B(_01063_),
    .C(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__a21oi_1 _07934_ (.A1(_00980_),
    .A2(_01063_),
    .B1(_01064_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand3_1 _07935_ (.A(_01004_),
    .B(_01008_),
    .C(_01009_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _07936_ (.A(_01010_),
    .B(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__or3_2 _07937_ (.A(_01065_),
    .B(_01066_),
    .C(_01068_),
    .X(_01069_));
 sky130_fd_sc_hd__and2b_1 _07938_ (.A_N(_01065_),
    .B(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__xnor2_2 _07939_ (.A(_01020_),
    .B(_01061_),
    .Y(_01071_));
 sky130_fd_sc_hd__and2b_1 _07940_ (.A_N(_01070_),
    .B(_01071_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_4 _07941_ (.A(_01062_),
    .B(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__a21oi_4 _07942_ (.A1(_01019_),
    .A2(_01073_),
    .B1(_01018_),
    .Y(_01074_));
 sky130_fd_sc_hd__a21o_1 _07943_ (.A1(_00899_),
    .A2(_00901_),
    .B1(_00898_),
    .X(_01075_));
 sky130_fd_sc_hd__a21oi_2 _07944_ (.A1(_00854_),
    .A2(_00857_),
    .B1(_00853_),
    .Y(_01076_));
 sky130_fd_sc_hd__o22a_1 _07945_ (.A1(net215),
    .A2(net34),
    .B1(net168),
    .B2(net80),
    .X(_01077_));
 sky130_fd_sc_hd__xnor2_2 _07946_ (.A(net115),
    .B(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__and2b_1 _07947_ (.A_N(_01076_),
    .B(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__xnor2_2 _07948_ (.A(_01076_),
    .B(_01078_),
    .Y(_01080_));
 sky130_fd_sc_hd__xor2_1 _07949_ (.A(_01075_),
    .B(_01080_),
    .X(_01081_));
 sky130_fd_sc_hd__a22o_1 _07950_ (.A1(_00305_),
    .A2(_00445_),
    .B1(_00450_),
    .B2(_00314_),
    .X(_01082_));
 sky130_fd_sc_hd__xor2_1 _07951_ (.A(net131),
    .B(_01082_),
    .X(_01083_));
 sky130_fd_sc_hd__o22a_1 _07952_ (.A1(net142),
    .A2(net53),
    .B1(net51),
    .B2(net141),
    .X(_01084_));
 sky130_fd_sc_hd__xnor2_1 _07953_ (.A(_00388_),
    .B(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__or2_1 _07954_ (.A(_01083_),
    .B(_01085_),
    .X(_01086_));
 sky130_fd_sc_hd__xnor2_1 _07955_ (.A(_01083_),
    .B(_01085_),
    .Y(_01087_));
 sky130_fd_sc_hd__o22a_1 _07956_ (.A1(net144),
    .A2(net55),
    .B1(net123),
    .B2(net96),
    .X(_01088_));
 sky130_fd_sc_hd__xnor2_1 _07957_ (.A(net127),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__xnor2_1 _07958_ (.A(_01087_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__o22a_1 _07959_ (.A1(net106),
    .A2(net92),
    .B1(net84),
    .B2(net102),
    .X(_01091_));
 sky130_fd_sc_hd__xnor2_2 _07960_ (.A(_00145_),
    .B(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__o22a_1 _07961_ (.A1(_00166_),
    .A2(net171),
    .B1(net137),
    .B2(net101),
    .X(_01093_));
 sky130_fd_sc_hd__xnor2_2 _07962_ (.A(net185),
    .B(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hd__nor2_1 _07963_ (.A(_01092_),
    .B(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__xor2_2 _07964_ (.A(_01092_),
    .B(_01094_),
    .X(_01096_));
 sky130_fd_sc_hd__o2bb2a_1 _07965_ (.A1_N(_00206_),
    .A2_N(net97),
    .B1(net94),
    .B2(net132),
    .X(_01097_));
 sky130_fd_sc_hd__xnor2_1 _07966_ (.A(net187),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__inv_2 _07967_ (.A(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__xnor2_1 _07968_ (.A(_01096_),
    .B(_01098_),
    .Y(_01100_));
 sky130_fd_sc_hd__or2_1 _07969_ (.A(net138),
    .B(net49),
    .X(_01101_));
 sky130_fd_sc_hd__a21o_1 _07970_ (.A1(_00438_),
    .A2(_00439_),
    .B1(net147),
    .X(_01102_));
 sky130_fd_sc_hd__nand3_1 _07971_ (.A(net86),
    .B(_01101_),
    .C(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__a21o_1 _07972_ (.A1(_01101_),
    .A2(_01102_),
    .B1(net86),
    .X(_01104_));
 sky130_fd_sc_hd__o32a_1 _07973_ (.A1(net158),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net47),
    .B2(net175),
    .X(_01105_));
 sky130_fd_sc_hd__xnor2_1 _07974_ (.A(_06505_),
    .B(_01105_),
    .Y(_01106_));
 sky130_fd_sc_hd__a21o_1 _07975_ (.A1(_01103_),
    .A2(_01104_),
    .B1(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__inv_2 _07976_ (.A(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand3_1 _07977_ (.A(_01103_),
    .B(_01104_),
    .C(_01106_),
    .Y(_01109_));
 sky130_fd_sc_hd__and3_1 _07978_ (.A(_01100_),
    .B(_01107_),
    .C(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__a21oi_1 _07979_ (.A1(_01107_),
    .A2(_01109_),
    .B1(_01100_),
    .Y(_01111_));
 sky130_fd_sc_hd__or3_1 _07980_ (.A(_01090_),
    .B(_01110_),
    .C(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__o21ai_1 _07981_ (.A1(_01110_),
    .A2(_01111_),
    .B1(_01090_),
    .Y(_01113_));
 sky130_fd_sc_hd__and3_1 _07982_ (.A(_01081_),
    .B(_01112_),
    .C(_01113_),
    .X(_01114_));
 sky130_fd_sc_hd__a21oi_1 _07983_ (.A1(_01112_),
    .A2(_01113_),
    .B1(_01081_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_2 _07984_ (.A(_01114_),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__o21a_2 _07985_ (.A1(_00866_),
    .A2(_00868_),
    .B1(_00865_),
    .X(_01117_));
 sky130_fd_sc_hd__o22a_2 _07986_ (.A1(net76),
    .A2(net163),
    .B1(net161),
    .B2(net73),
    .X(_01118_));
 sky130_fd_sc_hd__xnor2_4 _07987_ (.A(net205),
    .B(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__inv_2 _07988_ (.A(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__o22a_2 _07989_ (.A1(net300),
    .A2(net62),
    .B1(_00266_),
    .B2(_00187_),
    .X(_01121_));
 sky130_fd_sc_hd__xnor2_4 _07990_ (.A(net249),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__o22a_2 _07991_ (.A1(net70),
    .A2(net167),
    .B1(net165),
    .B2(net109),
    .X(_01123_));
 sky130_fd_sc_hd__xnor2_4 _07992_ (.A(net208),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _07993_ (.A(_01122_),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__xor2_4 _07994_ (.A(_01122_),
    .B(_01124_),
    .X(_01126_));
 sky130_fd_sc_hd__xnor2_4 _07995_ (.A(_01119_),
    .B(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__and2b_1 _07996_ (.A_N(_01117_),
    .B(_01127_),
    .X(_01128_));
 sky130_fd_sc_hd__xnor2_4 _07997_ (.A(_01117_),
    .B(_01127_),
    .Y(_01129_));
 sky130_fd_sc_hd__xnor2_4 _07998_ (.A(_00847_),
    .B(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__xnor2_4 _07999_ (.A(_01116_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__o21ba_2 _08000_ (.A1(_00887_),
    .A2(_00913_),
    .B1_N(_00886_),
    .X(_01132_));
 sky130_fd_sc_hd__a21boi_4 _08001_ (.A1(_00967_),
    .A2(_00971_),
    .B1_N(_00970_),
    .Y(_01133_));
 sky130_fd_sc_hd__o32ai_4 _08002_ (.A1(_00890_),
    .A2(_00892_),
    .A3(_00912_),
    .B1(_00911_),
    .B2(_00902_),
    .Y(_01134_));
 sky130_fd_sc_hd__o21ba_2 _08003_ (.A1(_00860_),
    .A2(_00869_),
    .B1_N(_00859_),
    .X(_01135_));
 sky130_fd_sc_hd__nor2_1 _08004_ (.A(net115),
    .B(_00872_),
    .Y(_01136_));
 sky130_fd_sc_hd__a21o_1 _08005_ (.A1(_00872_),
    .A2(_00884_),
    .B1(_01136_),
    .X(_01137_));
 sky130_fd_sc_hd__nor2_1 _08006_ (.A(_01135_),
    .B(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__xor2_4 _08007_ (.A(_01135_),
    .B(_01137_),
    .X(_01139_));
 sky130_fd_sc_hd__xnor2_4 _08008_ (.A(_01134_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__xor2_4 _08009_ (.A(_01133_),
    .B(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__nand2b_1 _08010_ (.A_N(_01132_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__xnor2_4 _08011_ (.A(_01132_),
    .B(_01141_),
    .Y(_01143_));
 sky130_fd_sc_hd__nand2_1 _08012_ (.A(_01131_),
    .B(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__xor2_4 _08013_ (.A(_01131_),
    .B(_01143_),
    .X(_01145_));
 sky130_fd_sc_hd__or2_2 _08014_ (.A(_01014_),
    .B(_01016_),
    .X(_01146_));
 sky130_fd_sc_hd__nand2_1 _08015_ (.A(_01145_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__xor2_4 _08016_ (.A(_01145_),
    .B(_01146_),
    .X(_01148_));
 sky130_fd_sc_hd__and2b_1 _08017_ (.A_N(_01148_),
    .B(_01074_),
    .X(_01149_));
 sky130_fd_sc_hd__nand2b_1 _08018_ (.A_N(_01074_),
    .B(_01148_),
    .Y(_01150_));
 sky130_fd_sc_hd__xor2_4 _08019_ (.A(_01019_),
    .B(_01073_),
    .X(_01151_));
 sky130_fd_sc_hd__xnor2_4 _08020_ (.A(_00936_),
    .B(_00965_),
    .Y(_01152_));
 sky130_fd_sc_hd__xnor2_2 _08021_ (.A(_01070_),
    .B(_01071_),
    .Y(_01153_));
 sky130_fd_sc_hd__and2_1 _08022_ (.A(_01152_),
    .B(_01153_),
    .X(_01154_));
 sky130_fd_sc_hd__xor2_4 _08023_ (.A(_01152_),
    .B(_01153_),
    .X(_01155_));
 sky130_fd_sc_hd__xor2_2 _08024_ (.A(_01059_),
    .B(_01060_),
    .X(_01156_));
 sky130_fd_sc_hd__o22a_1 _08025_ (.A1(net300),
    .A2(net105),
    .B1(_00266_),
    .B2(net101),
    .X(_01157_));
 sky130_fd_sc_hd__xnor2_2 _08026_ (.A(net249),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__a22o_1 _08027_ (.A1(_00281_),
    .A2(net97),
    .B1(_00323_),
    .B2(_00287_),
    .X(_01159_));
 sky130_fd_sc_hd__xor2_2 _08028_ (.A(net205),
    .B(_01159_),
    .X(_01160_));
 sky130_fd_sc_hd__or2_1 _08029_ (.A(_01158_),
    .B(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__xnor2_2 _08030_ (.A(_01032_),
    .B(_01034_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_1 _08031_ (.A(_01161_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _08032_ (.A(_01161_),
    .B(_01162_),
    .Y(_01164_));
 sky130_fd_sc_hd__xnor2_1 _08033_ (.A(_01161_),
    .B(_01162_),
    .Y(_01165_));
 sky130_fd_sc_hd__xnor2_2 _08034_ (.A(_01049_),
    .B(_01051_),
    .Y(_01166_));
 sky130_fd_sc_hd__a21o_1 _08035_ (.A1(_01164_),
    .A2(_01166_),
    .B1(_01163_),
    .X(_01167_));
 sky130_fd_sc_hd__o22a_1 _08036_ (.A1(net144),
    .A2(net106),
    .B1(net102),
    .B2(net142),
    .X(_01168_));
 sky130_fd_sc_hd__xnor2_2 _08037_ (.A(net172),
    .B(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__o22a_1 _08038_ (.A1(net146),
    .A2(net96),
    .B1(net55),
    .B2(net175),
    .X(_01170_));
 sky130_fd_sc_hd__xnor2_2 _08039_ (.A(net127),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__or2_1 _08040_ (.A(_01169_),
    .B(_01171_),
    .X(_01172_));
 sky130_fd_sc_hd__o22a_1 _08041_ (.A1(net140),
    .A2(_00306_),
    .B1(_00313_),
    .B2(net138),
    .X(_01173_));
 sky130_fd_sc_hd__xnor2_2 _08042_ (.A(net131),
    .B(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__xnor2_2 _08043_ (.A(_01169_),
    .B(_01171_),
    .Y(_01175_));
 sky130_fd_sc_hd__o21ai_2 _08044_ (.A1(_01174_),
    .A2(_01175_),
    .B1(_01172_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_1 _08045_ (.A(_01167_),
    .B(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor2_1 _08046_ (.A(net215),
    .B(net49),
    .Y(_01178_));
 sky130_fd_sc_hd__o22a_1 _08047_ (.A1(net169),
    .A2(net51),
    .B1(net158),
    .B2(net53),
    .X(_01179_));
 sky130_fd_sc_hd__xnor2_1 _08048_ (.A(net90),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__mux2_2 _08049_ (.A0(net87),
    .A1(_01180_),
    .S(_01178_),
    .X(_01181_));
 sky130_fd_sc_hd__xor2_2 _08050_ (.A(_01167_),
    .B(_01176_),
    .X(_01182_));
 sky130_fd_sc_hd__a21boi_2 _08051_ (.A1(_01181_),
    .A2(_01182_),
    .B1_N(_01177_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2b_1 _08052_ (.A_N(_01183_),
    .B(_01156_),
    .Y(_01184_));
 sky130_fd_sc_hd__xnor2_1 _08053_ (.A(_01028_),
    .B(_01029_),
    .Y(_01185_));
 sky130_fd_sc_hd__a21oi_1 _08054_ (.A1(_01008_),
    .A2(_01038_),
    .B1(_01039_),
    .Y(_01186_));
 sky130_fd_sc_hd__or3_1 _08055_ (.A(_01040_),
    .B(_01185_),
    .C(_01186_),
    .X(_01187_));
 sky130_fd_sc_hd__xor2_1 _08056_ (.A(_01056_),
    .B(_01058_),
    .X(_01188_));
 sky130_fd_sc_hd__o21ai_1 _08057_ (.A1(_01040_),
    .A2(_01186_),
    .B1(_01185_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand3_1 _08058_ (.A(_01187_),
    .B(_01188_),
    .C(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_2 _08059_ (.A(_01187_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__xor2_2 _08060_ (.A(_01156_),
    .B(_01183_),
    .X(_01192_));
 sky130_fd_sc_hd__nand2b_1 _08061_ (.A_N(_01192_),
    .B(_01191_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_2 _08062_ (.A(_01184_),
    .B(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__a21o_2 _08063_ (.A1(_01155_),
    .A2(_01194_),
    .B1(_01154_),
    .X(_01195_));
 sky130_fd_sc_hd__nand2_1 _08064_ (.A(_01151_),
    .B(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__a21oi_1 _08065_ (.A1(_01150_),
    .A2(_01196_),
    .B1(_01149_),
    .Y(_01197_));
 sky130_fd_sc_hd__xor2_4 _08066_ (.A(_01155_),
    .B(_01194_),
    .X(_01198_));
 sky130_fd_sc_hd__o21ai_1 _08067_ (.A1(_01065_),
    .A2(_01066_),
    .B1(_01068_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_4 _08068_ (.A(_01069_),
    .B(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__xor2_4 _08069_ (.A(_01191_),
    .B(_01192_),
    .X(_01201_));
 sky130_fd_sc_hd__xnor2_4 _08070_ (.A(_01200_),
    .B(_01201_),
    .Y(_01202_));
 sky130_fd_sc_hd__xor2_2 _08071_ (.A(_01158_),
    .B(_01160_),
    .X(_01203_));
 sky130_fd_sc_hd__o22a_1 _08072_ (.A1(net169),
    .A2(net53),
    .B1(net51),
    .B2(net215),
    .X(_01204_));
 sky130_fd_sc_hd__xnor2_1 _08073_ (.A(net90),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__and2_1 _08074_ (.A(_01203_),
    .B(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__a22o_1 _08075_ (.A1(net302),
    .A2(_00300_),
    .B1(net97),
    .B2(_00265_),
    .X(_01207_));
 sky130_fd_sc_hd__xnor2_2 _08076_ (.A(net250),
    .B(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__o22a_1 _08077_ (.A1(net163),
    .A2(net94),
    .B1(net92),
    .B2(net161),
    .X(_01209_));
 sky130_fd_sc_hd__xnor2_1 _08078_ (.A(net205),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_1 _08079_ (.A(_01208_),
    .B(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__xor2_1 _08080_ (.A(_01203_),
    .B(_01205_),
    .X(_01212_));
 sky130_fd_sc_hd__a21o_1 _08081_ (.A1(_01211_),
    .A2(_01212_),
    .B1(_01206_),
    .X(_01213_));
 sky130_fd_sc_hd__o22a_1 _08082_ (.A1(net167),
    .A2(net92),
    .B1(net84),
    .B2(net165),
    .X(_01214_));
 sky130_fd_sc_hd__xnor2_1 _08083_ (.A(net208),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__o22a_1 _08084_ (.A1(net144),
    .A2(net132),
    .B1(net122),
    .B2(net134),
    .X(_01216_));
 sky130_fd_sc_hd__xnor2_1 _08085_ (.A(net187),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__or2_1 _08086_ (.A(_01215_),
    .B(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__o22a_1 _08087_ (.A1(net171),
    .A2(net82),
    .B1(net125),
    .B2(net137),
    .X(_01219_));
 sky130_fd_sc_hd__xnor2_1 _08088_ (.A(net185),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__xnor2_1 _08089_ (.A(_01215_),
    .B(_01217_),
    .Y(_01221_));
 sky130_fd_sc_hd__or2_1 _08090_ (.A(_01220_),
    .B(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__and2_1 _08091_ (.A(_01218_),
    .B(_01222_),
    .X(_01223_));
 sky130_fd_sc_hd__a21boi_1 _08092_ (.A1(_01218_),
    .A2(_01222_),
    .B1_N(_01213_),
    .Y(_01224_));
 sky130_fd_sc_hd__o22a_1 _08093_ (.A1(net142),
    .A2(net106),
    .B1(net102),
    .B2(net140),
    .X(_01225_));
 sky130_fd_sc_hd__xnor2_2 _08094_ (.A(net172),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__o22a_1 _08095_ (.A1(net175),
    .A2(net96),
    .B1(net55),
    .B2(net158),
    .X(_01227_));
 sky130_fd_sc_hd__xnor2_2 _08096_ (.A(net127),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__o22a_1 _08097_ (.A1(net138),
    .A2(_00306_),
    .B1(net56),
    .B2(net146),
    .X(_01229_));
 sky130_fd_sc_hd__xnor2_1 _08098_ (.A(net131),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__xnor2_1 _08099_ (.A(_01226_),
    .B(_01228_),
    .Y(_01231_));
 sky130_fd_sc_hd__or2_1 _08100_ (.A(_01230_),
    .B(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__o21ai_4 _08101_ (.A1(_01226_),
    .A2(_01228_),
    .B1(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2b_1 _08102_ (.A_N(_01213_),
    .B(_01223_),
    .Y(_01234_));
 sky130_fd_sc_hd__xor2_2 _08103_ (.A(_01213_),
    .B(_01223_),
    .X(_01235_));
 sky130_fd_sc_hd__a21o_1 _08104_ (.A1(_01233_),
    .A2(_01234_),
    .B1(_01224_),
    .X(_01236_));
 sky130_fd_sc_hd__xor2_2 _08105_ (.A(_01181_),
    .B(_01182_),
    .X(_01237_));
 sky130_fd_sc_hd__xnor2_1 _08106_ (.A(_01165_),
    .B(_01166_),
    .Y(_01238_));
 sky130_fd_sc_hd__xor2_1 _08107_ (.A(_01174_),
    .B(_01175_),
    .X(_01239_));
 sky130_fd_sc_hd__xnor2_1 _08108_ (.A(_01238_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__xnor2_1 _08109_ (.A(_01178_),
    .B(_01180_),
    .Y(_01241_));
 sky130_fd_sc_hd__or2_1 _08110_ (.A(_01240_),
    .B(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__a21bo_1 _08111_ (.A1(_01238_),
    .A2(_01239_),
    .B1_N(_01242_),
    .X(_01243_));
 sky130_fd_sc_hd__xnor2_2 _08112_ (.A(_01236_),
    .B(_01237_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand2b_1 _08113_ (.A_N(_01244_),
    .B(_01243_),
    .Y(_01245_));
 sky130_fd_sc_hd__a21bo_2 _08114_ (.A1(_01236_),
    .A2(_01237_),
    .B1_N(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__and2b_1 _08115_ (.A_N(_01202_),
    .B(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__o21bai_4 _08116_ (.A1(_01200_),
    .A2(_01201_),
    .B1_N(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__or2_1 _08117_ (.A(_01198_),
    .B(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__xnor2_4 _08118_ (.A(_01202_),
    .B(_01246_),
    .Y(_01250_));
 sky130_fd_sc_hd__a21o_1 _08119_ (.A1(_01187_),
    .A2(_01189_),
    .B1(_01188_),
    .X(_01251_));
 sky130_fd_sc_hd__and2_2 _08120_ (.A(_01190_),
    .B(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__xnor2_2 _08121_ (.A(_01243_),
    .B(_01244_),
    .Y(_01253_));
 sky130_fd_sc_hd__and2_1 _08122_ (.A(_01252_),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__xnor2_4 _08123_ (.A(_01233_),
    .B(_01235_),
    .Y(_01255_));
 sky130_fd_sc_hd__o22a_1 _08124_ (.A1(net167),
    .A2(net84),
    .B1(net82),
    .B2(net165),
    .X(_01256_));
 sky130_fd_sc_hd__xnor2_1 _08125_ (.A(net208),
    .B(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__o22a_1 _08126_ (.A1(net144),
    .A2(net134),
    .B1(net132),
    .B2(net142),
    .X(_01258_));
 sky130_fd_sc_hd__xnor2_1 _08127_ (.A(net187),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__or2_1 _08128_ (.A(_01257_),
    .B(_01259_),
    .X(_01260_));
 sky130_fd_sc_hd__xnor2_1 _08129_ (.A(_01257_),
    .B(_01259_),
    .Y(_01261_));
 sky130_fd_sc_hd__o22a_1 _08130_ (.A1(net171),
    .A2(net125),
    .B1(net123),
    .B2(net137),
    .X(_01262_));
 sky130_fd_sc_hd__xnor2_1 _08131_ (.A(net185),
    .B(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__o21ai_2 _08132_ (.A1(_01261_),
    .A2(_01263_),
    .B1(_01260_),
    .Y(_01264_));
 sky130_fd_sc_hd__xor2_1 _08133_ (.A(_01208_),
    .B(_01210_),
    .X(_01265_));
 sky130_fd_sc_hd__nor2_1 _08134_ (.A(net215),
    .B(net53),
    .Y(_01266_));
 sky130_fd_sc_hd__mux2_1 _08135_ (.A0(net90),
    .A1(_01265_),
    .S(_01266_),
    .X(_01267_));
 sky130_fd_sc_hd__and2_1 _08136_ (.A(_01264_),
    .B(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__o22a_1 _08137_ (.A1(net140),
    .A2(net106),
    .B1(net102),
    .B2(net138),
    .X(_01269_));
 sky130_fd_sc_hd__xnor2_2 _08138_ (.A(net172),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__o22a_1 _08139_ (.A1(net169),
    .A2(net55),
    .B1(net158),
    .B2(net96),
    .X(_01271_));
 sky130_fd_sc_hd__xnor2_2 _08140_ (.A(net127),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__or2_1 _08141_ (.A(_01270_),
    .B(_01272_),
    .X(_01273_));
 sky130_fd_sc_hd__o22a_1 _08142_ (.A1(net146),
    .A2(_00306_),
    .B1(_00313_),
    .B2(net175),
    .X(_01274_));
 sky130_fd_sc_hd__xnor2_2 _08143_ (.A(net131),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__xnor2_2 _08144_ (.A(_01270_),
    .B(_01272_),
    .Y(_01276_));
 sky130_fd_sc_hd__o21ai_2 _08145_ (.A1(_01275_),
    .A2(_01276_),
    .B1(_01273_),
    .Y(_01277_));
 sky130_fd_sc_hd__xor2_2 _08146_ (.A(_01264_),
    .B(_01267_),
    .X(_01278_));
 sky130_fd_sc_hd__a21oi_2 _08147_ (.A1(_01277_),
    .A2(_01278_),
    .B1(_01268_),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2b_1 _08148_ (.A_N(_01279_),
    .B(_01255_),
    .Y(_01280_));
 sky130_fd_sc_hd__xnor2_1 _08149_ (.A(_01211_),
    .B(_01212_),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_1 _08150_ (.A(_01220_),
    .B(_01221_),
    .Y(_01282_));
 sky130_fd_sc_hd__and2_1 _08151_ (.A(_01222_),
    .B(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__nand2b_1 _08152_ (.A_N(_01281_),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__xnor2_1 _08153_ (.A(_01281_),
    .B(_01283_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(_01230_),
    .B(_01231_),
    .Y(_01286_));
 sky130_fd_sc_hd__and2_1 _08155_ (.A(_01232_),
    .B(_01286_),
    .X(_01287_));
 sky130_fd_sc_hd__nand2_1 _08156_ (.A(_01285_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_2 _08157_ (.A(_01284_),
    .B(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__xor2_4 _08158_ (.A(_01255_),
    .B(_01279_),
    .X(_01290_));
 sky130_fd_sc_hd__nand2b_1 _08159_ (.A_N(_01290_),
    .B(_01289_),
    .Y(_01291_));
 sky130_fd_sc_hd__nand2_4 _08160_ (.A(_01280_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__xor2_4 _08161_ (.A(_01252_),
    .B(_01253_),
    .X(_01293_));
 sky130_fd_sc_hd__a21oi_4 _08162_ (.A1(_01292_),
    .A2(_01293_),
    .B1(_01254_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2b_1 _08163_ (.A_N(_01294_),
    .B(_01250_),
    .Y(_01295_));
 sky130_fd_sc_hd__a21bo_1 _08164_ (.A1(_01198_),
    .A2(_01248_),
    .B1_N(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__nand2_1 _08165_ (.A(_01240_),
    .B(_01241_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_2 _08166_ (.A(_01242_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__xor2_4 _08167_ (.A(_01289_),
    .B(_01290_),
    .X(_01299_));
 sky130_fd_sc_hd__nor2_1 _08168_ (.A(_01298_),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__xnor2_2 _08169_ (.A(_01277_),
    .B(_01278_),
    .Y(_01301_));
 sky130_fd_sc_hd__o22a_1 _08170_ (.A1(net175),
    .A2(_00306_),
    .B1(_00313_),
    .B2(net158),
    .X(_01302_));
 sky130_fd_sc_hd__xnor2_1 _08171_ (.A(net130),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__o22a_1 _08172_ (.A1(net169),
    .A2(net96),
    .B1(net55),
    .B2(net215),
    .X(_01304_));
 sky130_fd_sc_hd__xnor2_1 _08173_ (.A(net127),
    .B(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__or2_1 _08174_ (.A(_01303_),
    .B(_01305_),
    .X(_01306_));
 sky130_fd_sc_hd__o22a_1 _08175_ (.A1(net167),
    .A2(net82),
    .B1(net125),
    .B2(net165),
    .X(_01307_));
 sky130_fd_sc_hd__xnor2_1 _08176_ (.A(net208),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__a22o_1 _08177_ (.A1(net302),
    .A2(net97),
    .B1(_00323_),
    .B2(_00265_),
    .X(_01309_));
 sky130_fd_sc_hd__xnor2_1 _08178_ (.A(net250),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_1 _08179_ (.A(_01308_),
    .B(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__o22a_1 _08180_ (.A1(net163),
    .A2(net92),
    .B1(net84),
    .B2(net161),
    .X(_01312_));
 sky130_fd_sc_hd__xnor2_2 _08181_ (.A(net205),
    .B(_01312_),
    .Y(_01313_));
 sky130_fd_sc_hd__inv_2 _08182_ (.A(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__xor2_1 _08183_ (.A(_01308_),
    .B(_01310_),
    .X(_01315_));
 sky130_fd_sc_hd__a21oi_1 _08184_ (.A1(_01314_),
    .A2(_01315_),
    .B1(_01311_),
    .Y(_01316_));
 sky130_fd_sc_hd__or2_1 _08185_ (.A(_01306_),
    .B(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__o22a_1 _08186_ (.A1(net138),
    .A2(net106),
    .B1(net102),
    .B2(net146),
    .X(_01318_));
 sky130_fd_sc_hd__xnor2_2 _08187_ (.A(net172),
    .B(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__o22a_1 _08188_ (.A1(net144),
    .A2(net137),
    .B1(net123),
    .B2(net171),
    .X(_01320_));
 sky130_fd_sc_hd__xnor2_1 _08189_ (.A(net185),
    .B(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__xor2_1 _08190_ (.A(_01319_),
    .B(_01321_),
    .X(_01322_));
 sky130_fd_sc_hd__o22a_1 _08191_ (.A1(net142),
    .A2(net134),
    .B1(net132),
    .B2(net140),
    .X(_01323_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(net188),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2b_1 _08193_ (.A_N(_01324_),
    .B(_01322_),
    .Y(_01325_));
 sky130_fd_sc_hd__o21ai_2 _08194_ (.A1(_01319_),
    .A2(_01321_),
    .B1(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__xor2_1 _08195_ (.A(_01306_),
    .B(_01316_),
    .X(_01327_));
 sky130_fd_sc_hd__a21boi_2 _08196_ (.A1(_01326_),
    .A2(_01327_),
    .B1_N(_01317_),
    .Y(_01328_));
 sky130_fd_sc_hd__or2_1 _08197_ (.A(_01301_),
    .B(_01328_),
    .X(_01329_));
 sky130_fd_sc_hd__xnor2_1 _08198_ (.A(_01261_),
    .B(_01263_),
    .Y(_01330_));
 sky130_fd_sc_hd__xnor2_1 _08199_ (.A(_01265_),
    .B(_01266_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2_1 _08200_ (.A(_01330_),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__and2_1 _08201_ (.A(_01330_),
    .B(_01331_),
    .X(_01333_));
 sky130_fd_sc_hd__nor2_1 _08202_ (.A(_01332_),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__xor2_2 _08203_ (.A(_01275_),
    .B(_01276_),
    .X(_01335_));
 sky130_fd_sc_hd__a21oi_2 _08204_ (.A1(_01334_),
    .A2(_01335_),
    .B1(_01332_),
    .Y(_01336_));
 sky130_fd_sc_hd__xnor2_2 _08205_ (.A(_01301_),
    .B(_01328_),
    .Y(_01337_));
 sky130_fd_sc_hd__o21ai_4 _08206_ (.A1(_01336_),
    .A2(_01337_),
    .B1(_01329_),
    .Y(_01338_));
 sky130_fd_sc_hd__xor2_4 _08207_ (.A(_01298_),
    .B(_01299_),
    .X(_01339_));
 sky130_fd_sc_hd__a21oi_4 _08208_ (.A1(_01338_),
    .A2(_01339_),
    .B1(_01300_),
    .Y(_01340_));
 sky130_fd_sc_hd__xnor2_4 _08209_ (.A(_01292_),
    .B(_01293_),
    .Y(_01341_));
 sky130_fd_sc_hd__and2_1 _08210_ (.A(_01340_),
    .B(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__or2_1 _08211_ (.A(_01285_),
    .B(_01287_),
    .X(_01343_));
 sky130_fd_sc_hd__nand2_1 _08212_ (.A(_01288_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__xnor2_1 _08213_ (.A(_01336_),
    .B(_01337_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _08214_ (.A(_01344_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__o22a_1 _08215_ (.A1(net169),
    .A2(_00313_),
    .B1(net158),
    .B2(net98),
    .X(_01347_));
 sky130_fd_sc_hd__xnor2_1 _08216_ (.A(net131),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__nor2_1 _08217_ (.A(net215),
    .B(net96),
    .Y(_01349_));
 sky130_fd_sc_hd__xnor2_1 _08218_ (.A(net127),
    .B(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__and2b_1 _08219_ (.A_N(_01348_),
    .B(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__o22a_1 _08220_ (.A1(net167),
    .A2(net125),
    .B1(net123),
    .B2(net165),
    .X(_01352_));
 sky130_fd_sc_hd__xnor2_1 _08221_ (.A(net208),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__o22a_1 _08222_ (.A1(net300),
    .A2(net94),
    .B1(net92),
    .B2(net247),
    .X(_01354_));
 sky130_fd_sc_hd__xnor2_1 _08223_ (.A(net249),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _08224_ (.A(_01353_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__o22a_1 _08225_ (.A1(net163),
    .A2(net84),
    .B1(net82),
    .B2(net161),
    .X(_01357_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_00236_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__inv_2 _08227_ (.A(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__xor2_1 _08228_ (.A(_01353_),
    .B(_01355_),
    .X(_01360_));
 sky130_fd_sc_hd__a21o_1 _08229_ (.A1(_01359_),
    .A2(_01360_),
    .B1(_01356_),
    .X(_01361_));
 sky130_fd_sc_hd__nand2_1 _08230_ (.A(_01351_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__o22a_1 _08231_ (.A1(net146),
    .A2(net106),
    .B1(_00167_),
    .B2(net175),
    .X(_01363_));
 sky130_fd_sc_hd__xnor2_2 _08232_ (.A(_00145_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__o22a_1 _08233_ (.A1(net144),
    .A2(net171),
    .B1(net137),
    .B2(net142),
    .X(_01365_));
 sky130_fd_sc_hd__xnor2_1 _08234_ (.A(net185),
    .B(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__xor2_1 _08235_ (.A(_01364_),
    .B(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__o22a_1 _08236_ (.A1(net141),
    .A2(net134),
    .B1(net132),
    .B2(net139),
    .X(_01368_));
 sky130_fd_sc_hd__xnor2_1 _08237_ (.A(net188),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__nand2b_1 _08238_ (.A_N(_01369_),
    .B(_01367_),
    .Y(_01370_));
 sky130_fd_sc_hd__o21ai_2 _08239_ (.A1(_01364_),
    .A2(_01366_),
    .B1(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__xor2_2 _08240_ (.A(_01351_),
    .B(_01361_),
    .X(_01372_));
 sky130_fd_sc_hd__a21bo_1 _08241_ (.A1(_01371_),
    .A2(_01372_),
    .B1_N(_01362_),
    .X(_01373_));
 sky130_fd_sc_hd__xor2_1 _08242_ (.A(_01326_),
    .B(_01327_),
    .X(_01374_));
 sky130_fd_sc_hd__nand2_1 _08243_ (.A(_01303_),
    .B(_01305_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _08244_ (.A(_01306_),
    .B(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__xnor2_1 _08245_ (.A(_01313_),
    .B(_01315_),
    .Y(_01377_));
 sky130_fd_sc_hd__xnor2_1 _08246_ (.A(_01376_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__xnor2_1 _08247_ (.A(_01322_),
    .B(_01324_),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _08248_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__a32o_1 _08249_ (.A1(_01306_),
    .A2(_01375_),
    .A3(_01377_),
    .B1(_01378_),
    .B2(_01379_),
    .X(_01381_));
 sky130_fd_sc_hd__xnor2_1 _08250_ (.A(_01373_),
    .B(_01374_),
    .Y(_01382_));
 sky130_fd_sc_hd__and2b_1 _08251_ (.A_N(_01382_),
    .B(_01381_),
    .X(_01383_));
 sky130_fd_sc_hd__a21o_1 _08252_ (.A1(_01373_),
    .A2(_01374_),
    .B1(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__xor2_1 _08253_ (.A(_01344_),
    .B(_01345_),
    .X(_01385_));
 sky130_fd_sc_hd__a21o_2 _08254_ (.A1(_01384_),
    .A2(_01385_),
    .B1(_01346_),
    .X(_01386_));
 sky130_fd_sc_hd__xor2_4 _08255_ (.A(_01338_),
    .B(_01339_),
    .X(_01387_));
 sky130_fd_sc_hd__nor2_1 _08256_ (.A(_01386_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__and2_1 _08257_ (.A(_01386_),
    .B(_01387_),
    .X(_01389_));
 sky130_fd_sc_hd__nand2_1 _08258_ (.A(_01386_),
    .B(_01387_),
    .Y(_01390_));
 sky130_fd_sc_hd__xor2_4 _08259_ (.A(_01386_),
    .B(_01387_),
    .X(_01391_));
 sky130_fd_sc_hd__xnor2_2 _08260_ (.A(_01334_),
    .B(_01335_),
    .Y(_01392_));
 sky130_fd_sc_hd__xor2_1 _08261_ (.A(_01381_),
    .B(_01382_),
    .X(_01393_));
 sky130_fd_sc_hd__or2_1 _08262_ (.A(_01392_),
    .B(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__xor2_2 _08263_ (.A(_01392_),
    .B(_01393_),
    .X(_01395_));
 sky130_fd_sc_hd__xnor2_2 _08264_ (.A(_01371_),
    .B(_01372_),
    .Y(_01396_));
 sky130_fd_sc_hd__o22a_1 _08265_ (.A1(net142),
    .A2(net171),
    .B1(net137),
    .B2(net141),
    .X(_01397_));
 sky130_fd_sc_hd__xnor2_1 _08266_ (.A(net185),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__o22a_1 _08267_ (.A1(_00136_),
    .A2(net134),
    .B1(net132),
    .B2(net146),
    .X(_01399_));
 sky130_fd_sc_hd__xnor2_1 _08268_ (.A(net187),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_1 _08269_ (.A(_01398_),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__and2_1 _08270_ (.A(_00319_),
    .B(_01401_),
    .X(_01402_));
 sky130_fd_sc_hd__o22a_1 _08271_ (.A1(net145),
    .A2(net165),
    .B1(net123),
    .B2(net167),
    .X(_01403_));
 sky130_fd_sc_hd__xnor2_1 _08272_ (.A(net208),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__o22a_1 _08273_ (.A1(net300),
    .A2(net92),
    .B1(net84),
    .B2(net247),
    .X(_01405_));
 sky130_fd_sc_hd__xnor2_1 _08274_ (.A(net249),
    .B(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _08275_ (.A(_01404_),
    .B(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__o22a_1 _08276_ (.A1(net163),
    .A2(net82),
    .B1(net125),
    .B2(net161),
    .X(_01408_));
 sky130_fd_sc_hd__xor2_1 _08277_ (.A(net205),
    .B(_01408_),
    .X(_01409_));
 sky130_fd_sc_hd__xor2_1 _08278_ (.A(_01404_),
    .B(_01406_),
    .X(_01410_));
 sky130_fd_sc_hd__a21o_1 _08279_ (.A1(_01409_),
    .A2(_01410_),
    .B1(_01407_),
    .X(_01411_));
 sky130_fd_sc_hd__or2_1 _08280_ (.A(_00319_),
    .B(_01401_),
    .X(_01412_));
 sky130_fd_sc_hd__nand2b_1 _08281_ (.A_N(_01402_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__a21oi_2 _08282_ (.A1(_01411_),
    .A2(_01412_),
    .B1(_01402_),
    .Y(_01414_));
 sky130_fd_sc_hd__xnor2_1 _08283_ (.A(_01348_),
    .B(_01350_),
    .Y(_01415_));
 sky130_fd_sc_hd__xnor2_1 _08284_ (.A(_01358_),
    .B(_01360_),
    .Y(_01416_));
 sky130_fd_sc_hd__xnor2_1 _08285_ (.A(_01367_),
    .B(_01369_),
    .Y(_01417_));
 sky130_fd_sc_hd__inv_2 _08286_ (.A(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__xnor2_1 _08287_ (.A(_01415_),
    .B(_01416_),
    .Y(_01419_));
 sky130_fd_sc_hd__or2_1 _08288_ (.A(_01418_),
    .B(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__a21bo_2 _08289_ (.A1(_01415_),
    .A2(_01416_),
    .B1_N(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__xnor2_2 _08290_ (.A(_01396_),
    .B(_01414_),
    .Y(_01422_));
 sky130_fd_sc_hd__and2b_1 _08291_ (.A_N(_01422_),
    .B(_01421_),
    .X(_01423_));
 sky130_fd_sc_hd__o21bai_2 _08292_ (.A1(_01396_),
    .A2(_01414_),
    .B1_N(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _08293_ (.A(_01395_),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__xnor2_1 _08294_ (.A(_01384_),
    .B(_01385_),
    .Y(_01426_));
 sky130_fd_sc_hd__and3_1 _08295_ (.A(_01394_),
    .B(_01425_),
    .C(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__xnor2_2 _08296_ (.A(_01395_),
    .B(_01424_),
    .Y(_01428_));
 sky130_fd_sc_hd__or2_1 _08297_ (.A(_01378_),
    .B(_01379_),
    .X(_01429_));
 sky130_fd_sc_hd__nand2_2 _08298_ (.A(_01380_),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__xor2_4 _08299_ (.A(_01421_),
    .B(_01422_),
    .X(_01431_));
 sky130_fd_sc_hd__nor2_1 _08300_ (.A(_01430_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__xor2_4 _08301_ (.A(_01430_),
    .B(_01431_),
    .X(_01433_));
 sky130_fd_sc_hd__xnor2_2 _08302_ (.A(_01411_),
    .B(_01413_),
    .Y(_01434_));
 sky130_fd_sc_hd__a22o_1 _08303_ (.A1(_06502_),
    .A2(_00241_),
    .B1(_00249_),
    .B2(_06513_),
    .X(_01435_));
 sky130_fd_sc_hd__xnor2_1 _08304_ (.A(net208),
    .B(_01435_),
    .Y(_01436_));
 sky130_fd_sc_hd__and3_1 _08305_ (.A(net302),
    .B(_00434_),
    .C(_00435_),
    .X(_01437_));
 sky130_fd_sc_hd__a21oi_1 _08306_ (.A1(_00442_),
    .A2(_00443_),
    .B1(net247),
    .Y(_01438_));
 sky130_fd_sc_hd__o21ai_1 _08307_ (.A1(_01437_),
    .A2(_01438_),
    .B1(net250),
    .Y(_01439_));
 sky130_fd_sc_hd__or3_1 _08308_ (.A(net250),
    .B(_01437_),
    .C(_01438_),
    .X(_01440_));
 sky130_fd_sc_hd__and3_1 _08309_ (.A(_01436_),
    .B(_01439_),
    .C(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__a22o_1 _08310_ (.A1(_00281_),
    .A2(_00450_),
    .B1(_00457_),
    .B2(_00287_),
    .X(_01442_));
 sky130_fd_sc_hd__xnor2_1 _08311_ (.A(_00236_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__a21o_1 _08312_ (.A1(_01439_),
    .A2(_01440_),
    .B1(_01436_),
    .X(_01444_));
 sky130_fd_sc_hd__nand2b_1 _08313_ (.A_N(_01441_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__a21o_1 _08314_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01441_),
    .X(_01446_));
 sky130_fd_sc_hd__o22a_1 _08315_ (.A1(net174),
    .A2(net106),
    .B1(net102),
    .B2(net158),
    .X(_01447_));
 sky130_fd_sc_hd__xnor2_2 _08316_ (.A(_00146_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _08317_ (.A(_01446_),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__a22o_1 _08318_ (.A1(_00224_),
    .A2(_00305_),
    .B1(_00314_),
    .B2(net213),
    .X(_01450_));
 sky130_fd_sc_hd__xor2_2 _08319_ (.A(net130),
    .B(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__xnor2_2 _08320_ (.A(_01446_),
    .B(_01448_),
    .Y(_01452_));
 sky130_fd_sc_hd__o21a_1 _08321_ (.A1(_01451_),
    .A2(_01452_),
    .B1(_01449_),
    .X(_01453_));
 sky130_fd_sc_hd__nand2b_1 _08322_ (.A_N(_01453_),
    .B(_01434_),
    .Y(_01454_));
 sky130_fd_sc_hd__o22a_1 _08323_ (.A1(net141),
    .A2(net171),
    .B1(net137),
    .B2(net138),
    .X(_01455_));
 sky130_fd_sc_hd__xnor2_1 _08324_ (.A(net185),
    .B(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__o22a_1 _08325_ (.A1(net146),
    .A2(net134),
    .B1(net132),
    .B2(net175),
    .X(_01457_));
 sky130_fd_sc_hd__xnor2_1 _08326_ (.A(net187),
    .B(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__or2_2 _08327_ (.A(_01456_),
    .B(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__and2_1 _08328_ (.A(_01398_),
    .B(_01400_),
    .X(_01460_));
 sky130_fd_sc_hd__or2_1 _08329_ (.A(_01401_),
    .B(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__xnor2_1 _08330_ (.A(_01459_),
    .B(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__xnor2_1 _08331_ (.A(_01409_),
    .B(_01410_),
    .Y(_01463_));
 sky130_fd_sc_hd__or2_1 _08332_ (.A(_01462_),
    .B(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__o21ai_2 _08333_ (.A1(_01459_),
    .A2(_01461_),
    .B1(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__xor2_2 _08334_ (.A(_01434_),
    .B(_01453_),
    .X(_01466_));
 sky130_fd_sc_hd__nand2b_1 _08335_ (.A_N(_01466_),
    .B(_01465_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_2 _08336_ (.A(_01454_),
    .B(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__a21oi_2 _08337_ (.A1(_01433_),
    .A2(_01468_),
    .B1(_01432_),
    .Y(_01469_));
 sky130_fd_sc_hd__or2_1 _08338_ (.A(_01428_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__xnor2_1 _08339_ (.A(_01428_),
    .B(_01469_),
    .Y(_01471_));
 sky130_fd_sc_hd__inv_2 _08340_ (.A(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__xor2_4 _08341_ (.A(_01433_),
    .B(_01468_),
    .X(_01473_));
 sky130_fd_sc_hd__nand2_1 _08342_ (.A(_01418_),
    .B(_01419_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_2 _08343_ (.A(_01420_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__xor2_2 _08344_ (.A(_01465_),
    .B(_01466_),
    .X(_01476_));
 sky130_fd_sc_hd__xor2_2 _08345_ (.A(_01451_),
    .B(_01452_),
    .X(_01477_));
 sky130_fd_sc_hd__o22a_1 _08346_ (.A1(net102),
    .A2(net169),
    .B1(net158),
    .B2(net106),
    .X(_01478_));
 sky130_fd_sc_hd__xnor2_1 _08347_ (.A(net172),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _08348_ (.A(net215),
    .B(_00306_),
    .Y(_01480_));
 sky130_fd_sc_hd__mux2_1 _08349_ (.A0(net131),
    .A1(_01479_),
    .S(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__inv_2 _08350_ (.A(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__and2_1 _08351_ (.A(_01477_),
    .B(_01482_),
    .X(_01483_));
 sky130_fd_sc_hd__a21o_1 _08352_ (.A1(_00442_),
    .A2(_00443_),
    .B1(net300),
    .X(_01484_));
 sky130_fd_sc_hd__nand2_1 _08353_ (.A(_00265_),
    .B(_00450_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21oi_1 _08354_ (.A1(_01484_),
    .A2(_01485_),
    .B1(_00256_),
    .Y(_01486_));
 sky130_fd_sc_hd__and3_1 _08355_ (.A(_00256_),
    .B(_01484_),
    .C(_01485_),
    .X(_01487_));
 sky130_fd_sc_hd__o22a_1 _08356_ (.A1(net145),
    .A2(net161),
    .B1(net123),
    .B2(net163),
    .X(_01488_));
 sky130_fd_sc_hd__xnor2_1 _08357_ (.A(net205),
    .B(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__or3_2 _08358_ (.A(_01486_),
    .B(_01487_),
    .C(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _08359_ (.A(_01456_),
    .B(_01458_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _08360_ (.A(_01459_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _08361_ (.A(_01490_),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__xnor2_1 _08362_ (.A(_01443_),
    .B(_01445_),
    .Y(_01494_));
 sky130_fd_sc_hd__xor2_1 _08363_ (.A(_01490_),
    .B(_01492_),
    .X(_01495_));
 sky130_fd_sc_hd__a21o_1 _08364_ (.A1(_01494_),
    .A2(_01495_),
    .B1(_01493_),
    .X(_01496_));
 sky130_fd_sc_hd__xnor2_2 _08365_ (.A(_01477_),
    .B(_01481_),
    .Y(_01497_));
 sky130_fd_sc_hd__a21o_1 _08366_ (.A1(_01496_),
    .A2(_01497_),
    .B1(_01483_),
    .X(_01498_));
 sky130_fd_sc_hd__xnor2_1 _08367_ (.A(_01475_),
    .B(_01476_),
    .Y(_01499_));
 sky130_fd_sc_hd__and2b_1 _08368_ (.A_N(_01499_),
    .B(_01498_),
    .X(_01500_));
 sky130_fd_sc_hd__o21bai_4 _08369_ (.A1(_01475_),
    .A2(_01476_),
    .B1_N(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__nor2_1 _08370_ (.A(_01473_),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_1 _08371_ (.A(_01462_),
    .B(_01463_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_1 _08372_ (.A(_01464_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__xnor2_2 _08373_ (.A(_01496_),
    .B(_01497_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _08374_ (.A(_01504_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__xor2_2 _08375_ (.A(_01504_),
    .B(_01505_),
    .X(_01507_));
 sky130_fd_sc_hd__o22a_1 _08376_ (.A1(net143),
    .A2(net167),
    .B1(net165),
    .B2(net140),
    .X(_01508_));
 sky130_fd_sc_hd__xnor2_1 _08377_ (.A(net208),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__o22a_1 _08378_ (.A1(net175),
    .A2(net134),
    .B1(net132),
    .B2(net158),
    .X(_01510_));
 sky130_fd_sc_hd__xnor2_1 _08379_ (.A(net187),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__or2_1 _08380_ (.A(_01509_),
    .B(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__o22a_1 _08381_ (.A1(net138),
    .A2(net171),
    .B1(net137),
    .B2(net146),
    .X(_01513_));
 sky130_fd_sc_hd__xnor2_1 _08382_ (.A(net185),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__xnor2_1 _08383_ (.A(_01509_),
    .B(_01511_),
    .Y(_01515_));
 sky130_fd_sc_hd__o21a_1 _08384_ (.A1(_01514_),
    .A2(_01515_),
    .B1(_01512_),
    .X(_01516_));
 sky130_fd_sc_hd__xnor2_1 _08385_ (.A(_01479_),
    .B(_01480_),
    .Y(_01517_));
 sky130_fd_sc_hd__and2b_1 _08386_ (.A_N(_01516_),
    .B(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__o21ai_1 _08387_ (.A1(_01486_),
    .A2(_01487_),
    .B1(_01489_),
    .Y(_01519_));
 sky130_fd_sc_hd__o22a_1 _08388_ (.A1(net215),
    .A2(net102),
    .B1(net169),
    .B2(net106),
    .X(_01520_));
 sky130_fd_sc_hd__xnor2_1 _08389_ (.A(_00146_),
    .B(_01520_),
    .Y(_01521_));
 sky130_fd_sc_hd__and3_1 _08390_ (.A(_01490_),
    .B(_01519_),
    .C(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__o22a_1 _08391_ (.A1(net144),
    .A2(net162),
    .B1(net160),
    .B2(net142),
    .X(_01523_));
 sky130_fd_sc_hd__xnor2_1 _08392_ (.A(net203),
    .B(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__a22o_1 _08393_ (.A1(net302),
    .A2(_00450_),
    .B1(_00457_),
    .B2(_00265_),
    .X(_01525_));
 sky130_fd_sc_hd__xnor2_1 _08394_ (.A(net250),
    .B(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__nor2_1 _08395_ (.A(_01524_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__a21o_1 _08396_ (.A1(_01490_),
    .A2(_01519_),
    .B1(_01521_),
    .X(_01528_));
 sky130_fd_sc_hd__nand2b_1 _08397_ (.A_N(_01522_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__a21oi_1 _08398_ (.A1(_01527_),
    .A2(_01528_),
    .B1(_01522_),
    .Y(_01530_));
 sky130_fd_sc_hd__xnor2_1 _08399_ (.A(_01516_),
    .B(_01517_),
    .Y(_01531_));
 sky130_fd_sc_hd__and2b_1 _08400_ (.A_N(_01530_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__or2_1 _08401_ (.A(_01518_),
    .B(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__and2_1 _08402_ (.A(_01507_),
    .B(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__xnor2_1 _08403_ (.A(_01498_),
    .B(_01499_),
    .Y(_01535_));
 sky130_fd_sc_hd__o21a_1 _08404_ (.A1(_01506_),
    .A2(_01534_),
    .B1(_01535_),
    .X(_01536_));
 sky130_fd_sc_hd__a21oi_1 _08405_ (.A1(_01473_),
    .A2(_01501_),
    .B1(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__xor2_1 _08406_ (.A(_01494_),
    .B(_01495_),
    .X(_01538_));
 sky130_fd_sc_hd__xnor2_1 _08407_ (.A(_01530_),
    .B(_01531_),
    .Y(_01539_));
 sky130_fd_sc_hd__o22a_1 _08408_ (.A1(net140),
    .A2(net166),
    .B1(net164),
    .B2(net138),
    .X(_01540_));
 sky130_fd_sc_hd__xnor2_2 _08409_ (.A(net208),
    .B(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__o22a_1 _08410_ (.A1(net132),
    .A2(net169),
    .B1(net158),
    .B2(net134),
    .X(_01542_));
 sky130_fd_sc_hd__xnor2_2 _08411_ (.A(net188),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__or2_1 _08412_ (.A(_01541_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__xnor2_2 _08413_ (.A(_01541_),
    .B(_01543_),
    .Y(_01545_));
 sky130_fd_sc_hd__o22a_1 _08414_ (.A1(net146),
    .A2(net170),
    .B1(net136),
    .B2(net175),
    .X(_01546_));
 sky130_fd_sc_hd__xor2_2 _08415_ (.A(_00171_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__inv_2 _08416_ (.A(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__o21a_1 _08417_ (.A1(_01545_),
    .A2(_01548_),
    .B1(_01544_),
    .X(_01549_));
 sky130_fd_sc_hd__xnor2_1 _08418_ (.A(_01514_),
    .B(_01515_),
    .Y(_01550_));
 sky130_fd_sc_hd__xnor2_1 _08419_ (.A(_01549_),
    .B(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2_1 _08420_ (.A(net214),
    .B(net106),
    .Y(_01552_));
 sky130_fd_sc_hd__and2_1 _08421_ (.A(_01524_),
    .B(_01526_),
    .X(_01553_));
 sky130_fd_sc_hd__nor2_1 _08422_ (.A(_01527_),
    .B(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__or2_1 _08423_ (.A(_00146_),
    .B(_01552_),
    .X(_01555_));
 sky130_fd_sc_hd__o31ai_2 _08424_ (.A1(net214),
    .A2(net106),
    .A3(_01554_),
    .B1(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _08425_ (.A(_01551_),
    .B(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__o21bai_1 _08426_ (.A1(_01549_),
    .A2(_01550_),
    .B1_N(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__xnor2_1 _08427_ (.A(_01538_),
    .B(_01539_),
    .Y(_01559_));
 sky130_fd_sc_hd__and2b_1 _08428_ (.A_N(_01559_),
    .B(_01558_),
    .X(_01560_));
 sky130_fd_sc_hd__a21o_1 _08429_ (.A1(_01538_),
    .A2(_01539_),
    .B1(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__xor2_2 _08430_ (.A(_01507_),
    .B(_01533_),
    .X(_01562_));
 sky130_fd_sc_hd__nor2_1 _08431_ (.A(_01561_),
    .B(_01562_),
    .Y(_01563_));
 sky130_fd_sc_hd__xor2_1 _08432_ (.A(_01527_),
    .B(_01529_),
    .X(_01564_));
 sky130_fd_sc_hd__xnor2_1 _08433_ (.A(_01551_),
    .B(_01556_),
    .Y(_01565_));
 sky130_fd_sc_hd__or2_1 _08434_ (.A(_01564_),
    .B(_01565_),
    .X(_01566_));
 sky130_fd_sc_hd__xnor2_1 _08435_ (.A(_01564_),
    .B(_01565_),
    .Y(_01567_));
 sky130_fd_sc_hd__xnor2_2 _08436_ (.A(_01545_),
    .B(_01547_),
    .Y(_01568_));
 sky130_fd_sc_hd__o22a_1 _08437_ (.A1(net138),
    .A2(net166),
    .B1(net164),
    .B2(net146),
    .X(_01569_));
 sky130_fd_sc_hd__xnor2_2 _08438_ (.A(net206),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__o22a_1 _08439_ (.A1(net144),
    .A2(net247),
    .B1(net123),
    .B2(net299),
    .X(_01571_));
 sky130_fd_sc_hd__xnor2_2 _08440_ (.A(net249),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_1 _08441_ (.A(_01570_),
    .B(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__a22o_1 _08442_ (.A1(_06513_),
    .A2(_00281_),
    .B1(_00287_),
    .B2(_06522_),
    .X(_01574_));
 sky130_fd_sc_hd__xnor2_2 _08443_ (.A(net205),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_01570_),
    .B(_01572_),
    .Y(_01576_));
 sky130_fd_sc_hd__xnor2_1 _08445_ (.A(_01570_),
    .B(_01572_),
    .Y(_01577_));
 sky130_fd_sc_hd__a21o_1 _08446_ (.A1(_01575_),
    .A2(_01576_),
    .B1(_01573_),
    .X(_01578_));
 sky130_fd_sc_hd__and2_1 _08447_ (.A(_01568_),
    .B(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__o22a_1 _08448_ (.A1(net174),
    .A2(net170),
    .B1(net136),
    .B2(net159),
    .X(_01580_));
 sky130_fd_sc_hd__xnor2_1 _08449_ (.A(net185),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__o22a_1 _08450_ (.A1(net214),
    .A2(net132),
    .B1(net168),
    .B2(net134),
    .X(_01582_));
 sky130_fd_sc_hd__xnor2_1 _08451_ (.A(net187),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__nor2_1 _08452_ (.A(_01581_),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__xor2_2 _08453_ (.A(_01568_),
    .B(_01578_),
    .X(_01585_));
 sky130_fd_sc_hd__a21o_1 _08454_ (.A1(_01584_),
    .A2(_01585_),
    .B1(_01579_),
    .X(_01586_));
 sky130_fd_sc_hd__nand2b_1 _08455_ (.A_N(_01567_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__xor2_1 _08456_ (.A(_01558_),
    .B(_01559_),
    .X(_01588_));
 sky130_fd_sc_hd__and3_1 _08457_ (.A(_01566_),
    .B(_01587_),
    .C(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__a21o_1 _08458_ (.A1(_01566_),
    .A2(_01587_),
    .B1(_01588_),
    .X(_01590_));
 sky130_fd_sc_hd__nand2b_1 _08459_ (.A_N(_01589_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__xnor2_2 _08460_ (.A(_01584_),
    .B(_01585_),
    .Y(_01592_));
 sky130_fd_sc_hd__xnor2_2 _08461_ (.A(_01552_),
    .B(_01554_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _08462_ (.A(_01592_),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__o22a_1 _08463_ (.A1(net147),
    .A2(net166),
    .B1(net164),
    .B2(net174),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_2 _08464_ (.A(net207),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__o22a_1 _08465_ (.A1(net299),
    .A2(net144),
    .B1(net142),
    .B2(net247),
    .X(_01597_));
 sky130_fd_sc_hd__xnor2_2 _08466_ (.A(net248),
    .B(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__nor2_1 _08467_ (.A(_01596_),
    .B(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__o22a_1 _08468_ (.A1(net140),
    .A2(net162),
    .B1(net160),
    .B2(net138),
    .X(_01600_));
 sky130_fd_sc_hd__xnor2_1 _08469_ (.A(net203),
    .B(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__inv_2 _08470_ (.A(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__xor2_2 _08471_ (.A(_01596_),
    .B(_01598_),
    .X(_01603_));
 sky130_fd_sc_hd__a21oi_2 _08472_ (.A1(_01602_),
    .A2(_01603_),
    .B1(_01599_),
    .Y(_01604_));
 sky130_fd_sc_hd__xnor2_2 _08473_ (.A(_01575_),
    .B(_01577_),
    .Y(_01605_));
 sky130_fd_sc_hd__nand2b_1 _08474_ (.A_N(_01604_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__o22a_1 _08475_ (.A1(net136),
    .A2(net168),
    .B1(net159),
    .B2(net170),
    .X(_01607_));
 sky130_fd_sc_hd__xnor2_1 _08476_ (.A(net183),
    .B(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _08477_ (.A(net214),
    .B(net134),
    .Y(_01609_));
 sky130_fd_sc_hd__xnor2_1 _08478_ (.A(net187),
    .B(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__and2b_1 _08479_ (.A_N(_01608_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__xnor2_2 _08480_ (.A(_01604_),
    .B(_01605_),
    .Y(_01612_));
 sky130_fd_sc_hd__a21bo_1 _08481_ (.A1(_01611_),
    .A2(_01612_),
    .B1_N(_01606_),
    .X(_01613_));
 sky130_fd_sc_hd__xnor2_2 _08482_ (.A(_01592_),
    .B(_01593_),
    .Y(_01614_));
 sky130_fd_sc_hd__and2b_1 _08483_ (.A_N(_01614_),
    .B(_01613_),
    .X(_01615_));
 sky130_fd_sc_hd__xnor2_1 _08484_ (.A(_01567_),
    .B(_01586_),
    .Y(_01616_));
 sky130_fd_sc_hd__or3_1 _08485_ (.A(_01594_),
    .B(_01615_),
    .C(_01616_),
    .X(_01617_));
 sky130_fd_sc_hd__inv_2 _08486_ (.A(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__and2_1 _08487_ (.A(_01581_),
    .B(_01583_),
    .X(_01619_));
 sky130_fd_sc_hd__or2_1 _08488_ (.A(_01584_),
    .B(_01619_),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_2 _08489_ (.A(_01611_),
    .B(_01612_),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_1 _08490_ (.A(_01620_),
    .B(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__xor2_2 _08491_ (.A(_01620_),
    .B(_01621_),
    .X(_01623_));
 sky130_fd_sc_hd__xnor2_1 _08492_ (.A(_01601_),
    .B(_01603_),
    .Y(_01624_));
 sky130_fd_sc_hd__and2b_1 _08493_ (.A_N(net186),
    .B(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__o22a_1 _08494_ (.A1(net299),
    .A2(net142),
    .B1(net140),
    .B2(net247),
    .X(_01626_));
 sky130_fd_sc_hd__xnor2_1 _08495_ (.A(net249),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__o22a_1 _08496_ (.A1(net138),
    .A2(net163),
    .B1(net160),
    .B2(net147),
    .X(_01628_));
 sky130_fd_sc_hd__xnor2_1 _08497_ (.A(net203),
    .B(_01628_),
    .Y(_01629_));
 sky130_fd_sc_hd__nor2_1 _08498_ (.A(_01627_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__xnor2_1 _08499_ (.A(net186),
    .B(_01624_),
    .Y(_01631_));
 sky130_fd_sc_hd__a21o_1 _08500_ (.A1(_01630_),
    .A2(_01631_),
    .B1(_01625_),
    .X(_01632_));
 sky130_fd_sc_hd__a21oi_2 _08501_ (.A1(_01623_),
    .A2(_01632_),
    .B1(_01622_),
    .Y(_01633_));
 sky130_fd_sc_hd__xor2_2 _08502_ (.A(_01613_),
    .B(_01614_),
    .X(_01634_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(_01633_),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__or2_1 _08504_ (.A(_01633_),
    .B(_01634_),
    .X(_01636_));
 sky130_fd_sc_hd__xnor2_2 _08505_ (.A(_01633_),
    .B(_01634_),
    .Y(_01637_));
 sky130_fd_sc_hd__xor2_1 _08506_ (.A(_01608_),
    .B(_01610_),
    .X(_01638_));
 sky130_fd_sc_hd__xnor2_1 _08507_ (.A(_01630_),
    .B(_01631_),
    .Y(_01639_));
 sky130_fd_sc_hd__or2_1 _08508_ (.A(_01638_),
    .B(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__xnor2_1 _08509_ (.A(_01638_),
    .B(_01639_),
    .Y(_01641_));
 sky130_fd_sc_hd__o22a_1 _08510_ (.A1(net147),
    .A2(net162),
    .B1(net160),
    .B2(net174),
    .X(_01642_));
 sky130_fd_sc_hd__xor2_2 _08511_ (.A(net204),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__o22a_1 _08512_ (.A1(net299),
    .A2(net141),
    .B1(net139),
    .B2(net247),
    .X(_01644_));
 sky130_fd_sc_hd__xnor2_2 _08513_ (.A(_00255_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__o22a_1 _08514_ (.A1(net174),
    .A2(net166),
    .B1(net164),
    .B2(net159),
    .X(_01646_));
 sky130_fd_sc_hd__xor2_1 _08515_ (.A(net207),
    .B(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__nand3_1 _08516_ (.A(_01643_),
    .B(_01645_),
    .C(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__o22a_1 _08517_ (.A1(net214),
    .A2(net136),
    .B1(net168),
    .B2(net170),
    .X(_01649_));
 sky130_fd_sc_hd__xor2_1 _08518_ (.A(net183),
    .B(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__a21o_1 _08519_ (.A1(_01643_),
    .A2(_01645_),
    .B1(_01647_),
    .X(_01651_));
 sky130_fd_sc_hd__nand3_1 _08520_ (.A(_01648_),
    .B(_01650_),
    .C(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _08521_ (.A(_01648_),
    .B(_01652_),
    .Y(_01653_));
 sky130_fd_sc_hd__inv_2 _08522_ (.A(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__o21ai_2 _08523_ (.A1(_01641_),
    .A2(_01654_),
    .B1(_01640_),
    .Y(_01655_));
 sky130_fd_sc_hd__xor2_2 _08524_ (.A(_01623_),
    .B(_01632_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_1 _08525_ (.A(_01655_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(_01655_),
    .B(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__xnor2_1 _08527_ (.A(_01641_),
    .B(_01654_),
    .Y(_01659_));
 sky130_fd_sc_hd__and2_1 _08528_ (.A(_01627_),
    .B(_01629_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_1 _08529_ (.A(_01630_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21o_1 _08530_ (.A1(_01648_),
    .A2(_01651_),
    .B1(_01650_),
    .X(_01662_));
 sky130_fd_sc_hd__and3_1 _08531_ (.A(_01652_),
    .B(_01661_),
    .C(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__nor2_1 _08532_ (.A(net214),
    .B(net170),
    .Y(_01664_));
 sky130_fd_sc_hd__o22a_1 _08533_ (.A1(net168),
    .A2(net164),
    .B1(net159),
    .B2(net166),
    .X(_01665_));
 sky130_fd_sc_hd__xnor2_1 _08534_ (.A(net206),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__mux2_1 _08535_ (.A0(net183),
    .A1(_01666_),
    .S(_01664_),
    .X(_01667_));
 sky130_fd_sc_hd__a21oi_1 _08536_ (.A1(_01652_),
    .A2(_01662_),
    .B1(_01661_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor3_1 _08537_ (.A(_01663_),
    .B(_01667_),
    .C(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_1 _08538_ (.A(_01663_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__or2_1 _08539_ (.A(_01659_),
    .B(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__xor2_1 _08540_ (.A(_01643_),
    .B(_01645_),
    .X(_01672_));
 sky130_fd_sc_hd__xor2_1 _08541_ (.A(_01664_),
    .B(_01666_),
    .X(_01673_));
 sky130_fd_sc_hd__nand2b_1 _08542_ (.A_N(_01673_),
    .B(_01672_),
    .Y(_01674_));
 sky130_fd_sc_hd__a21o_1 _08543_ (.A1(_06529_),
    .A2(_06530_),
    .B1(net299),
    .X(_01675_));
 sky130_fd_sc_hd__nand3_1 _08544_ (.A(_06477_),
    .B(_06478_),
    .C(_00265_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21oi_1 _08545_ (.A1(_01675_),
    .A2(_01676_),
    .B1(net248),
    .Y(_01677_));
 sky130_fd_sc_hd__and3_1 _08546_ (.A(net248),
    .B(_01675_),
    .C(_01676_),
    .X(_01678_));
 sky130_fd_sc_hd__o22a_1 _08547_ (.A1(net174),
    .A2(net162),
    .B1(net160),
    .B2(net159),
    .X(_01679_));
 sky130_fd_sc_hd__xnor2_1 _08548_ (.A(net203),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__or3_2 _08549_ (.A(_01677_),
    .B(_01678_),
    .C(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__xor2_1 _08550_ (.A(_01672_),
    .B(_01673_),
    .X(_01682_));
 sky130_fd_sc_hd__or2_1 _08551_ (.A(_01681_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__o21a_1 _08552_ (.A1(_01663_),
    .A2(_01668_),
    .B1(_01667_),
    .X(_01684_));
 sky130_fd_sc_hd__o211a_1 _08553_ (.A1(_01669_),
    .A2(_01684_),
    .B1(_01683_),
    .C1(_01674_),
    .X(_01685_));
 sky130_fd_sc_hd__a211o_1 _08554_ (.A1(_01674_),
    .A2(_01683_),
    .B1(_01684_),
    .C1(_01669_),
    .X(_01686_));
 sky130_fd_sc_hd__xor2_1 _08555_ (.A(_01681_),
    .B(_01682_),
    .X(_01687_));
 sky130_fd_sc_hd__o21ai_1 _08556_ (.A1(_01677_),
    .A2(_01678_),
    .B1(_01680_),
    .Y(_01688_));
 sky130_fd_sc_hd__o22a_1 _08557_ (.A1(net168),
    .A2(net166),
    .B1(net164),
    .B2(net214),
    .X(_01689_));
 sky130_fd_sc_hd__xor2_1 _08558_ (.A(net206),
    .B(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__and3_1 _08559_ (.A(_01681_),
    .B(_01688_),
    .C(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__o22a_1 _08560_ (.A1(net168),
    .A2(net160),
    .B1(net159),
    .B2(net162),
    .X(_01692_));
 sky130_fd_sc_hd__xnor2_2 _08561_ (.A(net203),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__a32o_1 _08562_ (.A1(reg1_val[0]),
    .A2(_06477_),
    .A3(_06478_),
    .B1(_06491_),
    .B2(_00265_),
    .X(_01694_));
 sky130_fd_sc_hd__xnor2_2 _08563_ (.A(_00255_),
    .B(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__or2_1 _08564_ (.A(_01693_),
    .B(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__a21oi_1 _08565_ (.A1(_01681_),
    .A2(_01688_),
    .B1(_01690_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor3_1 _08566_ (.A(_01691_),
    .B(_01696_),
    .C(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__or3_1 _08567_ (.A(_01691_),
    .B(_01696_),
    .C(_01697_),
    .X(_01699_));
 sky130_fd_sc_hd__nor3_1 _08568_ (.A(_01687_),
    .B(_01691_),
    .C(_01698_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21ai_1 _08569_ (.A1(_01691_),
    .A2(_01698_),
    .B1(_01687_),
    .Y(_01701_));
 sky130_fd_sc_hd__xnor2_2 _08570_ (.A(_01693_),
    .B(_01695_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(net213),
    .B(_00241_),
    .Y(_01703_));
 sky130_fd_sc_hd__and3_1 _08572_ (.A(net213),
    .B(_00241_),
    .C(_01702_),
    .X(_01704_));
 sky130_fd_sc_hd__a21oi_1 _08573_ (.A1(net206),
    .A2(_01703_),
    .B1(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__o21ai_1 _08574_ (.A1(_01691_),
    .A2(_01697_),
    .B1(_01696_),
    .Y(_01706_));
 sky130_fd_sc_hd__nand2_1 _08575_ (.A(_01699_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__a21o_1 _08576_ (.A1(_01699_),
    .A2(_01706_),
    .B1(_01705_),
    .X(_01708_));
 sky130_fd_sc_hd__and3_1 _08577_ (.A(_01699_),
    .B(_01705_),
    .C(_01706_),
    .X(_01709_));
 sky130_fd_sc_hd__o22a_1 _08578_ (.A1(net299),
    .A2(net174),
    .B1(net247),
    .B2(net159),
    .X(_01710_));
 sky130_fd_sc_hd__xnor2_1 _08579_ (.A(net248),
    .B(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__o22a_1 _08580_ (.A1(net168),
    .A2(net162),
    .B1(net160),
    .B2(net214),
    .X(_01712_));
 sky130_fd_sc_hd__xnor2_1 _08581_ (.A(net203),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__nor2_1 _08582_ (.A(_01711_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__xnor2_2 _08583_ (.A(_01702_),
    .B(_01703_),
    .Y(_01715_));
 sky130_fd_sc_hd__and2b_1 _08584_ (.A_N(_01715_),
    .B(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__xnor2_2 _08585_ (.A(_01714_),
    .B(_01715_),
    .Y(_01717_));
 sky130_fd_sc_hd__o22a_1 _08586_ (.A1(net168),
    .A2(net247),
    .B1(net159),
    .B2(net299),
    .X(_01718_));
 sky130_fd_sc_hd__xnor2_2 _08587_ (.A(net248),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__nor2_1 _08588_ (.A(net214),
    .B(net162),
    .Y(_01720_));
 sky130_fd_sc_hd__xor2_1 _08589_ (.A(net203),
    .B(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__nor2_1 _08590_ (.A(_01719_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__and2_1 _08591_ (.A(_01719_),
    .B(_01721_),
    .X(_01723_));
 sky130_fd_sc_hd__xor2_1 _08592_ (.A(_01719_),
    .B(_01720_),
    .X(_01724_));
 sky130_fd_sc_hd__a22o_1 _08593_ (.A1(reg1_val[0]),
    .A2(_00224_),
    .B1(_00265_),
    .B2(net213),
    .X(_01725_));
 sky130_fd_sc_hd__nand2b_1 _08594_ (.A_N(_01725_),
    .B(_06411_),
    .Y(_01726_));
 sky130_fd_sc_hd__or3_1 _08595_ (.A(net248),
    .B(_01724_),
    .C(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__xor2_1 _08596_ (.A(_01711_),
    .B(_01713_),
    .X(_01728_));
 sky130_fd_sc_hd__xnor2_1 _08597_ (.A(_01722_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__mux2_1 _08598_ (.A0(net203),
    .A1(_01719_),
    .S(_01720_),
    .X(_01730_));
 sky130_fd_sc_hd__inv_2 _08599_ (.A(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__a2bb2o_1 _08600_ (.A1_N(_01727_),
    .A2_N(_01729_),
    .B1(_01731_),
    .B2(_01728_),
    .X(_01732_));
 sky130_fd_sc_hd__a21o_1 _08601_ (.A1(_01717_),
    .A2(_01732_),
    .B1(_01716_),
    .X(_01733_));
 sky130_fd_sc_hd__xnor2_1 _08602_ (.A(_01705_),
    .B(_01707_),
    .Y(_01734_));
 sky130_fd_sc_hd__a21oi_2 _08603_ (.A1(_01708_),
    .A2(_01733_),
    .B1(_01709_),
    .Y(_01735_));
 sky130_fd_sc_hd__a21o_1 _08604_ (.A1(_01701_),
    .A2(_01735_),
    .B1(_01700_),
    .X(_01736_));
 sky130_fd_sc_hd__and2b_1 _08605_ (.A_N(_01700_),
    .B(_01701_),
    .X(_01737_));
 sky130_fd_sc_hd__a21o_1 _08606_ (.A1(_01686_),
    .A2(_01736_),
    .B1(_01685_),
    .X(_01738_));
 sky130_fd_sc_hd__a21o_1 _08607_ (.A1(_01659_),
    .A2(_01670_),
    .B1(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__and2b_1 _08608_ (.A_N(_01685_),
    .B(_01686_),
    .X(_01740_));
 sky130_fd_sc_hd__xnor2_1 _08609_ (.A(_01659_),
    .B(_01670_),
    .Y(_01741_));
 sky130_fd_sc_hd__a31o_1 _08610_ (.A1(_01658_),
    .A2(_01671_),
    .A3(_01739_),
    .B1(_01657_),
    .X(_01742_));
 sky130_fd_sc_hd__a311o_1 _08611_ (.A1(_01658_),
    .A2(_01671_),
    .A3(_01739_),
    .B1(_01657_),
    .C1(_01637_),
    .X(_01743_));
 sky130_fd_sc_hd__o21ai_1 _08612_ (.A1(_01594_),
    .A2(_01615_),
    .B1(_01616_),
    .Y(_01744_));
 sky130_fd_sc_hd__and2_1 _08613_ (.A(_01636_),
    .B(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__and2_1 _08614_ (.A(_01617_),
    .B(_01744_),
    .X(_01746_));
 sky130_fd_sc_hd__a21o_1 _08615_ (.A1(_01743_),
    .A2(_01745_),
    .B1(_01618_),
    .X(_01747_));
 sky130_fd_sc_hd__a211o_1 _08616_ (.A1(_01743_),
    .A2(_01745_),
    .B1(_01591_),
    .C1(_01618_),
    .X(_01748_));
 sky130_fd_sc_hd__nand2_1 _08617_ (.A(_01561_),
    .B(_01562_),
    .Y(_01749_));
 sky130_fd_sc_hd__a31o_2 _08618_ (.A1(_01590_),
    .A2(_01748_),
    .A3(_01749_),
    .B1(_01563_),
    .X(_01750_));
 sky130_fd_sc_hd__xnor2_4 _08619_ (.A(_01473_),
    .B(_01501_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor3_1 _08620_ (.A(_01506_),
    .B(_01534_),
    .C(_01535_),
    .Y(_01752_));
 sky130_fd_sc_hd__or2_2 _08621_ (.A(_01536_),
    .B(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__o32ai_4 _08622_ (.A1(_01750_),
    .A2(_01751_),
    .A3(_01753_),
    .B1(_01537_),
    .B2(_01502_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21o_1 _08623_ (.A1(_01394_),
    .A2(_01425_),
    .B1(_01426_),
    .X(_01755_));
 sky130_fd_sc_hd__a21oi_1 _08624_ (.A1(_01470_),
    .A2(_01755_),
    .B1(_01427_),
    .Y(_01756_));
 sky130_fd_sc_hd__and2b_1 _08625_ (.A_N(_01427_),
    .B(_01755_),
    .X(_01757_));
 sky130_fd_sc_hd__nand2b_2 _08626_ (.A_N(_01427_),
    .B(_01755_),
    .Y(_01758_));
 sky130_fd_sc_hd__a31o_2 _08627_ (.A1(_01472_),
    .A2(_01754_),
    .A3(_01757_),
    .B1(_01756_),
    .X(_01759_));
 sky130_fd_sc_hd__or2_1 _08628_ (.A(_01340_),
    .B(_01341_),
    .X(_01760_));
 sky130_fd_sc_hd__a21oi_1 _08629_ (.A1(_01390_),
    .A2(_01760_),
    .B1(_01342_),
    .Y(_01761_));
 sky130_fd_sc_hd__xor2_4 _08630_ (.A(_01340_),
    .B(_01341_),
    .X(_01762_));
 sky130_fd_sc_hd__a31o_4 _08631_ (.A1(_01391_),
    .A2(_01759_),
    .A3(_01762_),
    .B1(_01761_),
    .X(_01763_));
 sky130_fd_sc_hd__xor2_4 _08632_ (.A(_01198_),
    .B(_01248_),
    .X(_01764_));
 sky130_fd_sc_hd__xnor2_1 _08633_ (.A(_01198_),
    .B(_01248_),
    .Y(_01765_));
 sky130_fd_sc_hd__and2b_1 _08634_ (.A_N(_01250_),
    .B(_01294_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_4 _08635_ (.A(_01250_),
    .B(_01294_),
    .Y(_01767_));
 sky130_fd_sc_hd__and2_2 _08636_ (.A(_01764_),
    .B(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__a22oi_4 _08637_ (.A1(_01249_),
    .A2(_01296_),
    .B1(_01763_),
    .B2(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__xnor2_4 _08638_ (.A(_01074_),
    .B(_01148_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_1 _08639_ (.A(_01151_),
    .B(_01195_),
    .Y(_01771_));
 sky130_fd_sc_hd__xor2_4 _08640_ (.A(_01151_),
    .B(_01195_),
    .X(_01772_));
 sky130_fd_sc_hd__xnor2_1 _08641_ (.A(_01151_),
    .B(_01195_),
    .Y(_01773_));
 sky130_fd_sc_hd__and2_1 _08642_ (.A(_01770_),
    .B(_01772_),
    .X(_01774_));
 sky130_fd_sc_hd__and4_1 _08643_ (.A(_01249_),
    .B(_01296_),
    .C(_01770_),
    .D(_01772_),
    .X(_01775_));
 sky130_fd_sc_hd__a311oi_4 _08644_ (.A1(_01763_),
    .A2(_01768_),
    .A3(_01774_),
    .B1(_01775_),
    .C1(_01197_),
    .Y(_01776_));
 sky130_fd_sc_hd__o22a_1 _08645_ (.A1(net73),
    .A2(net167),
    .B1(net165),
    .B2(net70),
    .X(_01777_));
 sky130_fd_sc_hd__xnor2_1 _08646_ (.A(net208),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__o22a_1 _08647_ (.A1(net135),
    .A2(net101),
    .B1(_00311_),
    .B2(net132),
    .X(_01779_));
 sky130_fd_sc_hd__xnor2_1 _08648_ (.A(net187),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _08649_ (.A(_01778_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__xnor2_1 _08650_ (.A(_01778_),
    .B(_01780_),
    .Y(_01782_));
 sky130_fd_sc_hd__o22a_1 _08651_ (.A1(net109),
    .A2(net171),
    .B1(net137),
    .B2(net105),
    .X(_01783_));
 sky130_fd_sc_hd__xnor2_1 _08652_ (.A(net185),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _08653_ (.A(_01782_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__xor2_1 _08654_ (.A(_01782_),
    .B(_01784_),
    .X(_01786_));
 sky130_fd_sc_hd__o21a_1 _08655_ (.A1(_01087_),
    .A2(_01089_),
    .B1(_01086_),
    .X(_01787_));
 sky130_fd_sc_hd__and2b_1 _08656_ (.A_N(_01787_),
    .B(_01786_),
    .X(_01788_));
 sky130_fd_sc_hd__xnor2_1 _08657_ (.A(_01786_),
    .B(_01787_),
    .Y(_01789_));
 sky130_fd_sc_hd__xnor2_1 _08658_ (.A(_01107_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__o22a_1 _08659_ (.A1(net144),
    .A2(net53),
    .B1(net51),
    .B2(net142),
    .X(_01791_));
 sky130_fd_sc_hd__xnor2_2 _08660_ (.A(net90),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__o32a_1 _08661_ (.A1(net175),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net47),
    .B2(_06479_),
    .X(_01793_));
 sky130_fd_sc_hd__xnor2_2 _08662_ (.A(net111),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__and2_1 _08663_ (.A(_01792_),
    .B(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__xor2_2 _08664_ (.A(_01792_),
    .B(_01794_),
    .X(_01796_));
 sky130_fd_sc_hd__o22a_1 _08665_ (.A1(net140),
    .A2(net49),
    .B1(net14),
    .B2(net139),
    .X(_01797_));
 sky130_fd_sc_hd__xnor2_2 _08666_ (.A(net86),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__xor2_2 _08667_ (.A(_01796_),
    .B(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__a22o_1 _08668_ (.A1(_00305_),
    .A2(_00436_),
    .B1(_00445_),
    .B2(_00314_),
    .X(_01800_));
 sky130_fd_sc_hd__xnor2_1 _08669_ (.A(net131),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__o22a_1 _08670_ (.A1(net106),
    .A2(net94),
    .B1(net92),
    .B2(net102),
    .X(_01802_));
 sky130_fd_sc_hd__xnor2_1 _08671_ (.A(net172),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__nor2_1 _08672_ (.A(_00322_),
    .B(net125),
    .Y(_01804_));
 sky130_fd_sc_hd__a21oi_2 _08673_ (.A1(_00325_),
    .A2(_00326_),
    .B1(net123),
    .Y(_01805_));
 sky130_fd_sc_hd__or3_1 _08674_ (.A(net127),
    .B(_01804_),
    .C(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__o21ai_1 _08675_ (.A1(_01804_),
    .A2(_01805_),
    .B1(net127),
    .Y(_01807_));
 sky130_fd_sc_hd__a21o_1 _08676_ (.A1(_01806_),
    .A2(_01807_),
    .B1(_01803_),
    .X(_01808_));
 sky130_fd_sc_hd__nand3_1 _08677_ (.A(_01803_),
    .B(_01806_),
    .C(_01807_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand3_1 _08678_ (.A(_01801_),
    .B(_01808_),
    .C(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__a21o_1 _08679_ (.A1(_01808_),
    .A2(_01809_),
    .B1(_01801_),
    .X(_01811_));
 sky130_fd_sc_hd__nor2_1 _08680_ (.A(net215),
    .B(net31),
    .Y(_01812_));
 sky130_fd_sc_hd__or2_1 _08681_ (.A(net80),
    .B(_00411_),
    .X(_01813_));
 sky130_fd_sc_hd__a21o_1 _08682_ (.A1(_06514_),
    .A2(_06515_),
    .B1(net169),
    .X(_01814_));
 sky130_fd_sc_hd__nand3_1 _08683_ (.A(net115),
    .B(_01813_),
    .C(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__a21o_1 _08684_ (.A1(_01813_),
    .A2(_01814_),
    .B1(net115),
    .X(_01816_));
 sky130_fd_sc_hd__and3_1 _08685_ (.A(_01812_),
    .B(_01815_),
    .C(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__a21oi_1 _08686_ (.A1(_01815_),
    .A2(_01816_),
    .B1(_01812_),
    .Y(_01818_));
 sky130_fd_sc_hd__o211ai_2 _08687_ (.A1(_01817_),
    .A2(_01818_),
    .B1(_01810_),
    .C1(_01811_),
    .Y(_01819_));
 sky130_fd_sc_hd__a211o_1 _08688_ (.A1(_01810_),
    .A2(_01811_),
    .B1(_01817_),
    .C1(_01818_),
    .X(_01820_));
 sky130_fd_sc_hd__and3_1 _08689_ (.A(_01799_),
    .B(_01819_),
    .C(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__a21oi_1 _08690_ (.A1(_01819_),
    .A2(_01820_),
    .B1(_01799_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21o_1 _08691_ (.A1(_01120_),
    .A2(_01126_),
    .B1(_01125_),
    .X(_01823_));
 sky130_fd_sc_hd__o22a_1 _08692_ (.A1(net78),
    .A2(net163),
    .B1(net161),
    .B2(net76),
    .X(_01824_));
 sky130_fd_sc_hd__xnor2_2 _08693_ (.A(net204),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__o22a_1 _08694_ (.A1(net300),
    .A2(net65),
    .B1(_00251_),
    .B2(_00266_),
    .X(_01826_));
 sky130_fd_sc_hd__xnor2_2 _08695_ (.A(_00256_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__xor2_2 _08696_ (.A(_01825_),
    .B(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__a21oi_2 _08697_ (.A1(_01096_),
    .A2(_01099_),
    .B1(_01095_),
    .Y(_01829_));
 sky130_fd_sc_hd__and2b_1 _08698_ (.A_N(_01829_),
    .B(_01828_),
    .X(_01830_));
 sky130_fd_sc_hd__xnor2_2 _08699_ (.A(_01828_),
    .B(_01829_),
    .Y(_01831_));
 sky130_fd_sc_hd__xnor2_1 _08700_ (.A(_01823_),
    .B(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__or3_1 _08701_ (.A(_01821_),
    .B(_01822_),
    .C(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__o21ai_1 _08702_ (.A1(_01821_),
    .A2(_01822_),
    .B1(_01832_),
    .Y(_01834_));
 sky130_fd_sc_hd__and3_1 _08703_ (.A(_01790_),
    .B(_01833_),
    .C(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__a21oi_1 _08704_ (.A1(_01833_),
    .A2(_01834_),
    .B1(_01790_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _08705_ (.A(_01835_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__o21ba_1 _08706_ (.A1(_01115_),
    .A2(_01130_),
    .B1_N(_01114_),
    .X(_01838_));
 sky130_fd_sc_hd__a21o_1 _08707_ (.A1(_01134_),
    .A2(_01139_),
    .B1(_01138_),
    .X(_01839_));
 sky130_fd_sc_hd__a21o_1 _08708_ (.A1(_00847_),
    .A2(_01129_),
    .B1(_01128_),
    .X(_01840_));
 sky130_fd_sc_hd__a21oi_2 _08709_ (.A1(_01075_),
    .A2(_01080_),
    .B1(_01079_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21ba_1 _08710_ (.A1(_01090_),
    .A2(_01111_),
    .B1_N(_01110_),
    .X(_01842_));
 sky130_fd_sc_hd__nor2_1 _08711_ (.A(_01841_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__xor2_2 _08712_ (.A(_01841_),
    .B(_01842_),
    .X(_01844_));
 sky130_fd_sc_hd__xnor2_1 _08713_ (.A(_01840_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand2b_1 _08714_ (.A_N(_01845_),
    .B(_01839_),
    .Y(_01846_));
 sky130_fd_sc_hd__xnor2_1 _08715_ (.A(_01839_),
    .B(_01845_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2b_1 _08716_ (.A_N(_01838_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__xnor2_1 _08717_ (.A(_01838_),
    .B(_01847_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_01837_),
    .B(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__o21ai_1 _08719_ (.A1(_01133_),
    .A2(_01140_),
    .B1(_01142_),
    .Y(_01851_));
 sky130_fd_sc_hd__xnor2_1 _08720_ (.A(_01837_),
    .B(_01849_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2b_1 _08721_ (.A_N(_01852_),
    .B(_01851_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _08722_ (.A(_01846_),
    .B(_01848_),
    .Y(_01854_));
 sky130_fd_sc_hd__o22a_1 _08723_ (.A1(net144),
    .A2(net51),
    .B1(net123),
    .B2(net53),
    .X(_01855_));
 sky130_fd_sc_hd__xnor2_1 _08724_ (.A(net90),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__o22a_1 _08725_ (.A1(net138),
    .A2(net47),
    .B1(net12),
    .B2(net146),
    .X(_01857_));
 sky130_fd_sc_hd__xnor2_1 _08726_ (.A(net111),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_1 _08727_ (.A(_01856_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__xor2_1 _08728_ (.A(_01856_),
    .B(_01858_),
    .X(_01860_));
 sky130_fd_sc_hd__o22a_1 _08729_ (.A1(net143),
    .A2(net49),
    .B1(net14),
    .B2(net140),
    .X(_01861_));
 sky130_fd_sc_hd__xnor2_1 _08730_ (.A(net86),
    .B(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__xor2_1 _08731_ (.A(_01860_),
    .B(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__o22a_1 _08732_ (.A1(_00306_),
    .A2(net92),
    .B1(net84),
    .B2(_00313_),
    .X(_01864_));
 sky130_fd_sc_hd__xnor2_1 _08733_ (.A(net130),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__o22a_1 _08734_ (.A1(_00163_),
    .A2(_00311_),
    .B1(net94),
    .B2(net102),
    .X(_01866_));
 sky130_fd_sc_hd__xnor2_1 _08735_ (.A(net172),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__o22a_1 _08736_ (.A1(net96),
    .A2(net82),
    .B1(net125),
    .B2(net55),
    .X(_01868_));
 sky130_fd_sc_hd__xnor2_1 _08737_ (.A(net127),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__or2_1 _08738_ (.A(_01867_),
    .B(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__xnor2_1 _08739_ (.A(_01867_),
    .B(_01869_),
    .Y(_01871_));
 sky130_fd_sc_hd__or2_1 _08740_ (.A(_01865_),
    .B(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__xor2_1 _08741_ (.A(_01865_),
    .B(_01871_),
    .X(_01873_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(_06491_),
    .B(_06508_),
    .Y(_01874_));
 sky130_fd_sc_hd__a21o_1 _08743_ (.A1(_06514_),
    .A2(_06515_),
    .B1(_00411_),
    .X(_01875_));
 sky130_fd_sc_hd__nand3_1 _08744_ (.A(net115),
    .B(_01874_),
    .C(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a21o_1 _08745_ (.A1(_01874_),
    .A2(_01875_),
    .B1(net115),
    .X(_01877_));
 sky130_fd_sc_hd__a211o_1 _08746_ (.A1(_01876_),
    .A2(_01877_),
    .B1(_01825_),
    .C1(_01827_),
    .X(_01878_));
 sky130_fd_sc_hd__o211ai_2 _08747_ (.A1(_01825_),
    .A2(_01827_),
    .B1(_01876_),
    .C1(_01877_),
    .Y(_01879_));
 sky130_fd_sc_hd__o22a_1 _08748_ (.A1(net215),
    .A2(net30),
    .B1(net169),
    .B2(net31),
    .X(_01880_));
 sky130_fd_sc_hd__xnor2_1 _08749_ (.A(net118),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand3_2 _08750_ (.A(_01878_),
    .B(_01879_),
    .C(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21o_1 _08751_ (.A1(_01878_),
    .A2(_01879_),
    .B1(_01881_),
    .X(_01883_));
 sky130_fd_sc_hd__nand3_1 _08752_ (.A(_01873_),
    .B(_01882_),
    .C(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__a21o_1 _08753_ (.A1(_01882_),
    .A2(_01883_),
    .B1(_01873_),
    .X(_01885_));
 sky130_fd_sc_hd__and3_1 _08754_ (.A(_01863_),
    .B(_01884_),
    .C(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__a21oi_1 _08755_ (.A1(_01884_),
    .A2(_01885_),
    .B1(_01863_),
    .Y(_01887_));
 sky130_fd_sc_hd__o22a_1 _08756_ (.A1(net62),
    .A2(net162),
    .B1(net160),
    .B2(net78),
    .X(_01888_));
 sky130_fd_sc_hd__xnor2_2 _08757_ (.A(net204),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__o22a_1 _08758_ (.A1(net65),
    .A2(net247),
    .B1(net58),
    .B2(net300),
    .X(_01890_));
 sky130_fd_sc_hd__xnor2_2 _08759_ (.A(net249),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__nor2_1 _08760_ (.A(_01889_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__xnor2_1 _08761_ (.A(_01889_),
    .B(_01891_),
    .Y(_01893_));
 sky130_fd_sc_hd__a21bo_1 _08762_ (.A1(_01801_),
    .A2(_01809_),
    .B1_N(_01808_),
    .X(_01894_));
 sky130_fd_sc_hd__and2b_1 _08763_ (.A_N(_01893_),
    .B(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__xnor2_1 _08764_ (.A(_01893_),
    .B(_01894_),
    .Y(_01896_));
 sky130_fd_sc_hd__o21a_1 _08765_ (.A1(_01781_),
    .A2(_01785_),
    .B1(_01896_),
    .X(_01897_));
 sky130_fd_sc_hd__nor3_1 _08766_ (.A(_01781_),
    .B(_01785_),
    .C(_01896_),
    .Y(_01898_));
 sky130_fd_sc_hd__or2_1 _08767_ (.A(_01897_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__nor3_1 _08768_ (.A(_01886_),
    .B(_01887_),
    .C(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__o21ai_1 _08769_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01899_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2b_1 _08770_ (.A_N(_01900_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__o21bai_2 _08771_ (.A1(net118),
    .A2(_01812_),
    .B1_N(_01817_),
    .Y(_01903_));
 sky130_fd_sc_hd__o22a_1 _08772_ (.A1(_00155_),
    .A2(net137),
    .B1(net69),
    .B2(net171),
    .X(_01904_));
 sky130_fd_sc_hd__xnor2_2 _08773_ (.A(net185),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__o22a_1 _08774_ (.A1(net76),
    .A2(net167),
    .B1(net165),
    .B2(net73),
    .X(_01906_));
 sky130_fd_sc_hd__xnor2_2 _08775_ (.A(net208),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__o22a_1 _08776_ (.A1(net105),
    .A2(net134),
    .B1(net132),
    .B2(net101),
    .X(_01908_));
 sky130_fd_sc_hd__xnor2_2 _08777_ (.A(net187),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__or2_1 _08778_ (.A(_01907_),
    .B(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__xnor2_2 _08779_ (.A(_01907_),
    .B(_01909_),
    .Y(_01911_));
 sky130_fd_sc_hd__xor2_2 _08780_ (.A(_01905_),
    .B(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__a21o_1 _08781_ (.A1(_01796_),
    .A2(_01798_),
    .B1(_01795_),
    .X(_01913_));
 sky130_fd_sc_hd__xor2_2 _08782_ (.A(_01912_),
    .B(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__and2b_1 _08783_ (.A_N(_01903_),
    .B(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__xnor2_2 _08784_ (.A(_01903_),
    .B(_01914_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_2 _08785_ (.A(_01902_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a21bo_1 _08786_ (.A1(_01790_),
    .A2(_01834_),
    .B1_N(_01833_),
    .X(_01918_));
 sky130_fd_sc_hd__a21o_1 _08787_ (.A1(_01108_),
    .A2(_01789_),
    .B1(_01788_),
    .X(_01919_));
 sky130_fd_sc_hd__a21boi_2 _08788_ (.A1(_01799_),
    .A2(_01820_),
    .B1_N(_01819_),
    .Y(_01920_));
 sky130_fd_sc_hd__a21oi_2 _08789_ (.A1(_01823_),
    .A2(_01831_),
    .B1(_01830_),
    .Y(_01921_));
 sky130_fd_sc_hd__nor2_1 _08790_ (.A(_01920_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__xor2_2 _08791_ (.A(_01920_),
    .B(_01921_),
    .X(_01923_));
 sky130_fd_sc_hd__xnor2_2 _08792_ (.A(_01919_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__a21oi_2 _08793_ (.A1(_01840_),
    .A2(_01844_),
    .B1(_01843_),
    .Y(_01925_));
 sky130_fd_sc_hd__xnor2_2 _08794_ (.A(_01924_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2b_1 _08795_ (.A_N(_01926_),
    .B(_01918_),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_2 _08796_ (.A(_01918_),
    .B(_01926_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_01917_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_2 _08798_ (.A(_01917_),
    .B(_01928_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2b_1 _08799_ (.A_N(_01930_),
    .B(_01854_),
    .Y(_01931_));
 sky130_fd_sc_hd__xor2_1 _08800_ (.A(_01854_),
    .B(_01930_),
    .X(_01932_));
 sky130_fd_sc_hd__and3_1 _08801_ (.A(_01850_),
    .B(_01853_),
    .C(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__a21o_1 _08802_ (.A1(_01850_),
    .A2(_01853_),
    .B1(_01932_),
    .X(_01934_));
 sky130_fd_sc_hd__inv_2 _08803_ (.A(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2b_2 _08804_ (.A_N(_01933_),
    .B(_01934_),
    .Y(_01936_));
 sky130_fd_sc_hd__xor2_1 _08805_ (.A(_01851_),
    .B(_01852_),
    .X(_01937_));
 sky130_fd_sc_hd__and3_1 _08806_ (.A(_01144_),
    .B(_01147_),
    .C(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__a21o_1 _08807_ (.A1(_01144_),
    .A2(_01147_),
    .B1(_01937_),
    .X(_01939_));
 sky130_fd_sc_hd__nand2b_2 _08808_ (.A_N(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__or2_1 _08809_ (.A(_01936_),
    .B(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__o21ai_2 _08810_ (.A1(_01924_),
    .A2(_01925_),
    .B1(_01927_),
    .Y(_01942_));
 sky130_fd_sc_hd__o21a_1 _08811_ (.A1(_01905_),
    .A2(_01911_),
    .B1(_01910_),
    .X(_01943_));
 sky130_fd_sc_hd__and2_1 _08812_ (.A(_00812_),
    .B(_00814_),
    .X(_01944_));
 sky130_fd_sc_hd__or2_1 _08813_ (.A(_00815_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__a21oi_1 _08814_ (.A1(_01870_),
    .A2(_01872_),
    .B1(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__and3_1 _08815_ (.A(_01870_),
    .B(_01872_),
    .C(_01945_),
    .X(_01947_));
 sky130_fd_sc_hd__nor2_1 _08816_ (.A(_01946_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__and2b_1 _08817_ (.A_N(_01943_),
    .B(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__xnor2_2 _08818_ (.A(_01943_),
    .B(_01948_),
    .Y(_01950_));
 sky130_fd_sc_hd__o22a_1 _08819_ (.A1(net147),
    .A2(net80),
    .B1(net34),
    .B2(net175),
    .X(_01951_));
 sky130_fd_sc_hd__xnor2_1 _08820_ (.A(net115),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _08821_ (.A(net215),
    .B(net38),
    .Y(_01953_));
 sky130_fd_sc_hd__xnor2_2 _08822_ (.A(_06472_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__and2_1 _08823_ (.A(_01952_),
    .B(_01954_),
    .X(_01955_));
 sky130_fd_sc_hd__xnor2_1 _08824_ (.A(_01952_),
    .B(_01954_),
    .Y(_01956_));
 sky130_fd_sc_hd__o22a_1 _08825_ (.A1(net30),
    .A2(net168),
    .B1(net158),
    .B2(_06527_),
    .X(_01957_));
 sky130_fd_sc_hd__xnor2_1 _08826_ (.A(net118),
    .B(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__and2b_1 _08827_ (.A_N(_01956_),
    .B(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__and2b_1 _08828_ (.A_N(_01958_),
    .B(_01956_),
    .X(_01960_));
 sky130_fd_sc_hd__or2_2 _08829_ (.A(_01959_),
    .B(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__inv_2 _08830_ (.A(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__xnor2_2 _08831_ (.A(_00806_),
    .B(_00808_),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(net121),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__xnor2_2 _08833_ (.A(net121),
    .B(_01963_),
    .Y(_01965_));
 sky130_fd_sc_hd__xor2_2 _08834_ (.A(_01892_),
    .B(_01965_),
    .X(_01966_));
 sky130_fd_sc_hd__o22a_1 _08835_ (.A1(net53),
    .A2(net125),
    .B1(net123),
    .B2(net51),
    .X(_01967_));
 sky130_fd_sc_hd__xnor2_1 _08836_ (.A(net90),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__o32a_1 _08837_ (.A1(net138),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net47),
    .B2(net140),
    .X(_01969_));
 sky130_fd_sc_hd__xnor2_1 _08838_ (.A(net111),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(_01968_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xor2_1 _08840_ (.A(_01968_),
    .B(_01970_),
    .X(_01972_));
 sky130_fd_sc_hd__o22a_1 _08841_ (.A1(net144),
    .A2(_00433_),
    .B1(net14),
    .B2(net142),
    .X(_01973_));
 sky130_fd_sc_hd__xnor2_1 _08842_ (.A(_00431_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _08843_ (.A(_01972_),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__or2_1 _08844_ (.A(_01972_),
    .B(_01974_),
    .X(_01976_));
 sky130_fd_sc_hd__and2_1 _08845_ (.A(_01975_),
    .B(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__and2b_1 _08846_ (.A_N(_01966_),
    .B(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__xnor2_2 _08847_ (.A(_01966_),
    .B(_01977_),
    .Y(_01979_));
 sky130_fd_sc_hd__xnor2_2 _08848_ (.A(_01961_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__and2_1 _08849_ (.A(_01950_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__xor2_2 _08850_ (.A(_01950_),
    .B(_01980_),
    .X(_01982_));
 sky130_fd_sc_hd__a21bo_1 _08851_ (.A1(_01860_),
    .A2(_01862_),
    .B1_N(_01859_),
    .X(_01983_));
 sky130_fd_sc_hd__o22a_1 _08852_ (.A1(_00306_),
    .A2(net94),
    .B1(_00329_),
    .B2(_00313_),
    .X(_01984_));
 sky130_fd_sc_hd__xnor2_1 _08853_ (.A(net131),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__o22a_1 _08854_ (.A1(_00163_),
    .A2(net101),
    .B1(_00311_),
    .B2(net102),
    .X(_01986_));
 sky130_fd_sc_hd__xnor2_1 _08855_ (.A(net172),
    .B(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__o22a_1 _08856_ (.A1(net96),
    .A2(net84),
    .B1(net82),
    .B2(net55),
    .X(_01988_));
 sky130_fd_sc_hd__xnor2_1 _08857_ (.A(net127),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__or2_1 _08858_ (.A(_01987_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__nand2_1 _08859_ (.A(_01987_),
    .B(_01989_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _08860_ (.A(_01990_),
    .B(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__xor2_1 _08861_ (.A(_01985_),
    .B(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__xnor2_1 _08862_ (.A(_01983_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__a21oi_1 _08863_ (.A1(_01878_),
    .A2(_01882_),
    .B1(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__and3_1 _08864_ (.A(_01878_),
    .B(_01882_),
    .C(_01994_),
    .X(_01996_));
 sky130_fd_sc_hd__nor2_1 _08865_ (.A(_01995_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__xor2_2 _08866_ (.A(_01982_),
    .B(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__a21oi_2 _08867_ (.A1(_01901_),
    .A2(_01916_),
    .B1(_01900_),
    .Y(_01999_));
 sky130_fd_sc_hd__a21o_1 _08868_ (.A1(_01912_),
    .A2(_01913_),
    .B1(_01915_),
    .X(_02000_));
 sky130_fd_sc_hd__a21bo_2 _08869_ (.A1(_01863_),
    .A2(_01885_),
    .B1_N(_01884_),
    .X(_02001_));
 sky130_fd_sc_hd__nor2_2 _08870_ (.A(_01895_),
    .B(_01897_),
    .Y(_02002_));
 sky130_fd_sc_hd__o21a_1 _08871_ (.A1(_01895_),
    .A2(_01897_),
    .B1(_02001_),
    .X(_02003_));
 sky130_fd_sc_hd__xnor2_4 _08872_ (.A(_02001_),
    .B(_02002_),
    .Y(_02004_));
 sky130_fd_sc_hd__xnor2_2 _08873_ (.A(_02000_),
    .B(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__a21o_1 _08874_ (.A1(_01919_),
    .A2(_01923_),
    .B1(_01922_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2b_1 _08875_ (.A_N(_02005_),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__xnor2_2 _08876_ (.A(_02005_),
    .B(_02006_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2b_1 _08877_ (.A_N(_01999_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__xnor2_2 _08878_ (.A(_01999_),
    .B(_02008_),
    .Y(_02010_));
 sky130_fd_sc_hd__and2_1 _08879_ (.A(_01998_),
    .B(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__xor2_2 _08880_ (.A(_01998_),
    .B(_02010_),
    .X(_02012_));
 sky130_fd_sc_hd__xnor2_2 _08881_ (.A(_01942_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__a21oi_2 _08882_ (.A1(_01929_),
    .A2(_01931_),
    .B1(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__and3_1 _08883_ (.A(_01929_),
    .B(_01931_),
    .C(_02013_),
    .X(_02015_));
 sky130_fd_sc_hd__or2_4 _08884_ (.A(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__a21o_2 _08885_ (.A1(_01942_),
    .A2(_02012_),
    .B1(_02011_),
    .X(_02017_));
 sky130_fd_sc_hd__nand2_4 _08886_ (.A(_02007_),
    .B(_02009_),
    .Y(_02018_));
 sky130_fd_sc_hd__o31a_1 _08887_ (.A1(_01889_),
    .A2(_01891_),
    .A3(_01965_),
    .B1(_01964_),
    .X(_02019_));
 sky130_fd_sc_hd__nand2_1 _08888_ (.A(_00779_),
    .B(_00780_),
    .Y(_02020_));
 sky130_fd_sc_hd__and2_1 _08889_ (.A(_00781_),
    .B(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__o21ai_1 _08890_ (.A1(_01955_),
    .A2(_01959_),
    .B1(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__or3_1 _08891_ (.A(_01955_),
    .B(_01959_),
    .C(_02021_),
    .X(_02023_));
 sky130_fd_sc_hd__and2_1 _08892_ (.A(_02022_),
    .B(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__nand2b_1 _08893_ (.A_N(_02019_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__xnor2_1 _08894_ (.A(_02019_),
    .B(_02024_),
    .Y(_02026_));
 sky130_fd_sc_hd__o21ai_1 _08895_ (.A1(_01985_),
    .A2(_01992_),
    .B1(_01990_),
    .Y(_02027_));
 sky130_fd_sc_hd__nand2_1 _08896_ (.A(_00537_),
    .B(_00539_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand2_1 _08897_ (.A(_00540_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__a21oi_1 _08898_ (.A1(_01971_),
    .A2(_01975_),
    .B1(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__and3_1 _08899_ (.A(_01971_),
    .B(_01975_),
    .C(_02029_),
    .X(_02031_));
 sky130_fd_sc_hd__or2_1 _08900_ (.A(_02030_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__and2b_1 _08901_ (.A_N(_02032_),
    .B(_02027_),
    .X(_02033_));
 sky130_fd_sc_hd__xor2_1 _08902_ (.A(_02027_),
    .B(_02032_),
    .X(_02034_));
 sky130_fd_sc_hd__nor2_1 _08903_ (.A(_00794_),
    .B(_00796_),
    .Y(_02035_));
 sky130_fd_sc_hd__nor2_1 _08904_ (.A(_00797_),
    .B(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__a21o_1 _08905_ (.A1(_00810_),
    .A2(_00816_),
    .B1(_00815_),
    .X(_02037_));
 sky130_fd_sc_hd__or2_1 _08906_ (.A(_00769_),
    .B(_00771_),
    .X(_02038_));
 sky130_fd_sc_hd__and2_1 _08907_ (.A(_00772_),
    .B(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__nand3_1 _08908_ (.A(_00817_),
    .B(_02037_),
    .C(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__a21o_1 _08909_ (.A1(_00817_),
    .A2(_02037_),
    .B1(_02039_),
    .X(_02041_));
 sky130_fd_sc_hd__and3_1 _08910_ (.A(_02036_),
    .B(_02040_),
    .C(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__a21oi_1 _08911_ (.A1(_02040_),
    .A2(_02041_),
    .B1(_02036_),
    .Y(_02043_));
 sky130_fd_sc_hd__or3_1 _08912_ (.A(_02034_),
    .B(_02042_),
    .C(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__o21ai_1 _08913_ (.A1(_02042_),
    .A2(_02043_),
    .B1(_02034_),
    .Y(_02045_));
 sky130_fd_sc_hd__and3_1 _08914_ (.A(_02026_),
    .B(_02044_),
    .C(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__a21oi_1 _08915_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_02026_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_2 _08916_ (.A(_02046_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__a21o_1 _08917_ (.A1(_01982_),
    .A2(_01997_),
    .B1(_01981_),
    .X(_02049_));
 sky130_fd_sc_hd__a21o_2 _08918_ (.A1(_01983_),
    .A2(_01993_),
    .B1(_01995_),
    .X(_02050_));
 sky130_fd_sc_hd__or2_2 _08919_ (.A(_01946_),
    .B(_01949_),
    .X(_02051_));
 sky130_fd_sc_hd__a21oi_2 _08920_ (.A1(_01962_),
    .A2(_01979_),
    .B1(_01978_),
    .Y(_02052_));
 sky130_fd_sc_hd__o21ba_1 _08921_ (.A1(_01946_),
    .A2(_01949_),
    .B1_N(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__xnor2_4 _08922_ (.A(_02051_),
    .B(_02052_),
    .Y(_02054_));
 sky130_fd_sc_hd__xnor2_4 _08923_ (.A(_02050_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__a21oi_4 _08924_ (.A1(_02000_),
    .A2(_02004_),
    .B1(_02003_),
    .Y(_02056_));
 sky130_fd_sc_hd__xnor2_2 _08925_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2b_1 _08926_ (.A_N(_02057_),
    .B(_02049_),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_2 _08927_ (.A(_02049_),
    .B(_02057_),
    .Y(_02059_));
 sky130_fd_sc_hd__and2_1 _08928_ (.A(_02048_),
    .B(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__xor2_4 _08929_ (.A(_02048_),
    .B(_02059_),
    .X(_02061_));
 sky130_fd_sc_hd__xor2_4 _08930_ (.A(_02018_),
    .B(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__nor2_1 _08931_ (.A(_02017_),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__xnor2_4 _08932_ (.A(_02017_),
    .B(_02062_),
    .Y(_02064_));
 sky130_fd_sc_hd__or4_2 _08933_ (.A(_01776_),
    .B(_01941_),
    .C(_02016_),
    .D(_02064_),
    .X(_02065_));
 sky130_fd_sc_hd__a21oi_1 _08934_ (.A1(_02017_),
    .A2(_02062_),
    .B1(_02014_),
    .Y(_02066_));
 sky130_fd_sc_hd__or2_1 _08935_ (.A(_02063_),
    .B(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__a21oi_1 _08936_ (.A1(_01934_),
    .A2(_01939_),
    .B1(_01933_),
    .Y(_02068_));
 sky130_fd_sc_hd__inv_2 _08937_ (.A(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__o32a_1 _08938_ (.A1(_02016_),
    .A2(_02064_),
    .A3(_02069_),
    .B1(_02066_),
    .B2(_02063_),
    .X(_02070_));
 sky130_fd_sc_hd__o21ai_4 _08939_ (.A1(_02055_),
    .A2(_02056_),
    .B1(_02058_),
    .Y(_02071_));
 sky130_fd_sc_hd__xnor2_4 _08940_ (.A(_00818_),
    .B(_00820_),
    .Y(_02072_));
 sky130_fd_sc_hd__xor2_1 _08941_ (.A(_00760_),
    .B(_00761_),
    .X(_02073_));
 sky130_fd_sc_hd__xnor2_1 _08942_ (.A(_00782_),
    .B(_00783_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_02073_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__or2_1 _08944_ (.A(_02073_),
    .B(_02074_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_2 _08945_ (.A(_02075_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__xor2_4 _08946_ (.A(_02072_),
    .B(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__a21bo_1 _08947_ (.A1(_02026_),
    .A2(_02045_),
    .B1_N(_02044_),
    .X(_02079_));
 sky130_fd_sc_hd__a21o_1 _08948_ (.A1(_02050_),
    .A2(_02054_),
    .B1(_02053_),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_1 _08949_ (.A(_02022_),
    .B(_02025_),
    .Y(_02081_));
 sky130_fd_sc_hd__or2_1 _08950_ (.A(_02030_),
    .B(_02033_),
    .X(_02082_));
 sky130_fd_sc_hd__a21boi_2 _08951_ (.A1(_02036_),
    .A2(_02041_),
    .B1_N(_02040_),
    .Y(_02083_));
 sky130_fd_sc_hd__o21ba_1 _08952_ (.A1(_02030_),
    .A2(_02033_),
    .B1_N(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__xnor2_2 _08953_ (.A(_02082_),
    .B(_02083_),
    .Y(_02085_));
 sky130_fd_sc_hd__xor2_2 _08954_ (.A(_02081_),
    .B(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__xnor2_2 _08955_ (.A(_02080_),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__nand2b_1 _08956_ (.A_N(_02087_),
    .B(_02079_),
    .Y(_02088_));
 sky130_fd_sc_hd__xnor2_2 _08957_ (.A(_02079_),
    .B(_02087_),
    .Y(_02089_));
 sky130_fd_sc_hd__and2_1 _08958_ (.A(_02078_),
    .B(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__xor2_4 _08959_ (.A(_02078_),
    .B(_02089_),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_4 _08960_ (.A(_02071_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__a21oi_4 _08961_ (.A1(_02018_),
    .A2(_02061_),
    .B1(_02060_),
    .Y(_02093_));
 sky130_fd_sc_hd__or2_1 _08962_ (.A(_02092_),
    .B(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__xnor2_4 _08963_ (.A(_02092_),
    .B(_02093_),
    .Y(_02095_));
 sky130_fd_sc_hd__a21o_2 _08964_ (.A1(_02071_),
    .A2(_02091_),
    .B1(_02090_),
    .X(_02096_));
 sky130_fd_sc_hd__a21bo_2 _08965_ (.A1(_02080_),
    .A2(_02086_),
    .B1_N(_02088_),
    .X(_02097_));
 sky130_fd_sc_hd__xor2_4 _08966_ (.A(_00828_),
    .B(_00830_),
    .X(_02098_));
 sky130_fd_sc_hd__o21ai_2 _08967_ (.A1(_02072_),
    .A2(_02077_),
    .B1(_02075_),
    .Y(_02099_));
 sky130_fd_sc_hd__a21o_1 _08968_ (.A1(_02081_),
    .A2(_02085_),
    .B1(_02084_),
    .X(_02100_));
 sky130_fd_sc_hd__xor2_1 _08969_ (.A(_00821_),
    .B(_00822_),
    .X(_02101_));
 sky130_fd_sc_hd__xnor2_1 _08970_ (.A(_02100_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2b_1 _08971_ (.A_N(_02102_),
    .B(_02099_),
    .Y(_02103_));
 sky130_fd_sc_hd__xnor2_2 _08972_ (.A(_02099_),
    .B(_02102_),
    .Y(_02104_));
 sky130_fd_sc_hd__and2_1 _08973_ (.A(_02098_),
    .B(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__xor2_4 _08974_ (.A(_02098_),
    .B(_02104_),
    .X(_02106_));
 sky130_fd_sc_hd__xnor2_4 _08975_ (.A(_02097_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__and2b_1 _08976_ (.A_N(_02096_),
    .B(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__nand2b_1 _08977_ (.A_N(_02107_),
    .B(_02096_),
    .Y(_02109_));
 sky130_fd_sc_hd__xnor2_4 _08978_ (.A(_02096_),
    .B(_02107_),
    .Y(_02110_));
 sky130_fd_sc_hd__nand2b_1 _08979_ (.A_N(_02095_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__a21oi_2 _08980_ (.A1(_02097_),
    .A2(_02106_),
    .B1(_02105_),
    .Y(_02112_));
 sky130_fd_sc_hd__a21bo_1 _08981_ (.A1(_02100_),
    .A2(_02101_),
    .B1_N(_02103_),
    .X(_02113_));
 sky130_fd_sc_hd__xor2_1 _08982_ (.A(_00555_),
    .B(_00556_),
    .X(_02114_));
 sky130_fd_sc_hd__xnor2_1 _08983_ (.A(_00831_),
    .B(_00832_),
    .Y(_02115_));
 sky130_fd_sc_hd__xnor2_1 _08984_ (.A(_02114_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2b_1 _08985_ (.A_N(_02116_),
    .B(_02113_),
    .Y(_02117_));
 sky130_fd_sc_hd__xor2_2 _08986_ (.A(_02113_),
    .B(_02116_),
    .X(_02118_));
 sky130_fd_sc_hd__or2_1 _08987_ (.A(_02112_),
    .B(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_02112_),
    .B(_02118_),
    .Y(_02120_));
 sky130_fd_sc_hd__xor2_1 _08989_ (.A(_02112_),
    .B(_02118_),
    .X(_02121_));
 sky130_fd_sc_hd__nand2_2 _08990_ (.A(_02119_),
    .B(_02120_),
    .Y(_02122_));
 sky130_fd_sc_hd__a21bo_2 _08991_ (.A1(_02114_),
    .A2(_02115_),
    .B1_N(_02117_),
    .X(_02123_));
 sky130_fd_sc_hd__xor2_4 _08992_ (.A(_00834_),
    .B(_00835_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_1 _08993_ (.A(_02123_),
    .B(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand2_1 _08994_ (.A(_02123_),
    .B(_02124_),
    .Y(_02126_));
 sky130_fd_sc_hd__xnor2_4 _08995_ (.A(_02123_),
    .B(_02124_),
    .Y(_02127_));
 sky130_fd_sc_hd__a2111o_1 _08996_ (.A1(_02065_),
    .A2(_02070_),
    .B1(_02111_),
    .C1(_02122_),
    .D1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__a21boi_1 _08997_ (.A1(_02123_),
    .A2(_02124_),
    .B1_N(_02119_),
    .Y(_02129_));
 sky130_fd_sc_hd__a21o_1 _08998_ (.A1(_02094_),
    .A2(_02109_),
    .B1(_02108_),
    .X(_02130_));
 sky130_fd_sc_hd__o32a_1 _08999_ (.A1(_02122_),
    .A2(_02127_),
    .A3(_02130_),
    .B1(_02129_),
    .B2(_02125_),
    .X(_02131_));
 sky130_fd_sc_hd__nand2_2 _09000_ (.A(_02128_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__xor2_4 _09001_ (.A(_00839_),
    .B(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__and2_1 _09002_ (.A(net303),
    .B(_05403_),
    .X(_02134_));
 sky130_fd_sc_hd__nand2_4 _09003_ (.A(net303),
    .B(_05403_),
    .Y(_02135_));
 sky130_fd_sc_hd__a21o_1 _09004_ (.A1(_01150_),
    .A2(_01939_),
    .B1(_01938_),
    .X(_02136_));
 sky130_fd_sc_hd__a21o_1 _09005_ (.A1(_01390_),
    .A2(_01755_),
    .B1(_01388_),
    .X(_02137_));
 sky130_fd_sc_hd__o2bb2a_1 _09006_ (.A1_N(_01501_),
    .A2_N(_01473_),
    .B1(_01469_),
    .B2(_01428_),
    .X(_02138_));
 sky130_fd_sc_hd__and2b_1 _09007_ (.A_N(_01536_),
    .B(_01749_),
    .X(_02139_));
 sky130_fd_sc_hd__xnor2_2 _09008_ (.A(_01561_),
    .B(_01562_),
    .Y(_02140_));
 sky130_fd_sc_hd__and2_1 _09009_ (.A(_01590_),
    .B(_01744_),
    .X(_02141_));
 sky130_fd_sc_hd__nand2_1 _09010_ (.A(_01636_),
    .B(_01658_),
    .Y(_02142_));
 sky130_fd_sc_hd__xnor2_1 _09011_ (.A(_01655_),
    .B(_01656_),
    .Y(_02143_));
 sky130_fd_sc_hd__a21oi_2 _09012_ (.A1(_01671_),
    .A2(_01739_),
    .B1(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__o21a_1 _09013_ (.A1(_02142_),
    .A2(_02144_),
    .B1(_01635_),
    .X(_02145_));
 sky130_fd_sc_hd__o211ai_2 _09014_ (.A1(_02142_),
    .A2(_02144_),
    .B1(_01635_),
    .C1(_01746_),
    .Y(_02146_));
 sky130_fd_sc_hd__a21o_1 _09015_ (.A1(_02141_),
    .A2(_02146_),
    .B1(_01589_),
    .X(_02147_));
 sky130_fd_sc_hd__a211o_1 _09016_ (.A1(_02141_),
    .A2(_02146_),
    .B1(_01589_),
    .C1(_02140_),
    .X(_02148_));
 sky130_fd_sc_hd__a21o_1 _09017_ (.A1(_02139_),
    .A2(_02148_),
    .B1(_01752_),
    .X(_02149_));
 sky130_fd_sc_hd__a21o_1 _09018_ (.A1(_01428_),
    .A2(_01469_),
    .B1(_02138_),
    .X(_02150_));
 sky130_fd_sc_hd__a2111o_1 _09019_ (.A1(_02139_),
    .A2(_02148_),
    .B1(_01471_),
    .C1(_01751_),
    .D1(_01752_),
    .X(_02151_));
 sky130_fd_sc_hd__and2_2 _09020_ (.A(_02150_),
    .B(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__a2111o_1 _09021_ (.A1(_02150_),
    .A2(_02151_),
    .B1(_01388_),
    .C1(_01389_),
    .D1(_01758_),
    .X(_02153_));
 sky130_fd_sc_hd__nand2_2 _09022_ (.A(_02137_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__nand2_1 _09023_ (.A(_01762_),
    .B(_01767_),
    .Y(_02155_));
 sky130_fd_sc_hd__a2111o_2 _09024_ (.A1(_02137_),
    .A2(_02153_),
    .B1(_02155_),
    .C1(_01773_),
    .D1(_01765_),
    .X(_02156_));
 sky130_fd_sc_hd__a21o_1 _09025_ (.A1(_01295_),
    .A2(_01760_),
    .B1(_01766_),
    .X(_02157_));
 sky130_fd_sc_hd__a22oi_1 _09026_ (.A1(_01151_),
    .A2(_01195_),
    .B1(_01198_),
    .B2(_01248_),
    .Y(_02158_));
 sky130_fd_sc_hd__o32a_2 _09027_ (.A1(_01765_),
    .A2(_01773_),
    .A3(_02157_),
    .B1(_02158_),
    .B2(_01771_),
    .X(_02159_));
 sky130_fd_sc_hd__nand2_2 _09028_ (.A(_02156_),
    .B(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand3b_1 _09029_ (.A_N(_01938_),
    .B(_01939_),
    .C(_01770_),
    .Y(_02161_));
 sky130_fd_sc_hd__a21o_1 _09030_ (.A1(_02156_),
    .A2(_02159_),
    .B1(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__nand2_2 _09031_ (.A(_02136_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_4 _09032_ (.A(_01936_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__o21ai_1 _09033_ (.A1(net248),
    .A2(_01726_),
    .B1(_01724_),
    .Y(_02165_));
 sky130_fd_sc_hd__and2_1 _09034_ (.A(_01727_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__nor2_1 _09035_ (.A(_01726_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__o31ai_1 _09036_ (.A1(net203),
    .A2(_01722_),
    .A3(_01723_),
    .B1(_01727_),
    .Y(_02168_));
 sky130_fd_sc_hd__xor2_1 _09037_ (.A(_01729_),
    .B(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_1 _09038_ (.A(_02167_),
    .B(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__xor2_2 _09039_ (.A(_01717_),
    .B(_01732_),
    .X(_02171_));
 sky130_fd_sc_hd__nor2_1 _09040_ (.A(_02170_),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__xnor2_2 _09041_ (.A(_01733_),
    .B(_01734_),
    .Y(_02173_));
 sky130_fd_sc_hd__and2_1 _09042_ (.A(_02172_),
    .B(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__xor2_2 _09043_ (.A(_01735_),
    .B(_01737_),
    .X(_02175_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_02174_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__xnor2_2 _09045_ (.A(_01736_),
    .B(_01740_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _09046_ (.A(_02176_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__xnor2_2 _09047_ (.A(_01738_),
    .B(_01741_),
    .Y(_02179_));
 sky130_fd_sc_hd__and2_1 _09048_ (.A(_02178_),
    .B(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__and3_1 _09049_ (.A(_01671_),
    .B(_01739_),
    .C(_02143_),
    .X(_02181_));
 sky130_fd_sc_hd__or2_1 _09050_ (.A(_02144_),
    .B(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__o211a_1 _09051_ (.A1(_02144_),
    .A2(_02181_),
    .B1(_02179_),
    .C1(_02178_),
    .X(_02183_));
 sky130_fd_sc_hd__xnor2_2 _09052_ (.A(_01637_),
    .B(_01742_),
    .Y(_02184_));
 sky130_fd_sc_hd__and2_1 _09053_ (.A(_02183_),
    .B(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__xnor2_2 _09054_ (.A(_01746_),
    .B(_02145_),
    .Y(_02186_));
 sky130_fd_sc_hd__xnor2_2 _09055_ (.A(_01591_),
    .B(_01747_),
    .Y(_02187_));
 sky130_fd_sc_hd__and3_1 _09056_ (.A(_02185_),
    .B(_02186_),
    .C(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__xnor2_2 _09057_ (.A(_02140_),
    .B(_02147_),
    .Y(_02189_));
 sky130_fd_sc_hd__xnor2_2 _09058_ (.A(_01750_),
    .B(_01753_),
    .Y(_02190_));
 sky130_fd_sc_hd__and3_1 _09059_ (.A(_02188_),
    .B(_02189_),
    .C(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__xnor2_4 _09060_ (.A(_01751_),
    .B(_02149_),
    .Y(_02192_));
 sky130_fd_sc_hd__xnor2_4 _09061_ (.A(_01472_),
    .B(_01754_),
    .Y(_02193_));
 sky130_fd_sc_hd__and3_1 _09062_ (.A(_02191_),
    .B(_02192_),
    .C(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__xnor2_4 _09063_ (.A(_01758_),
    .B(_02152_),
    .Y(_02195_));
 sky130_fd_sc_hd__xnor2_4 _09064_ (.A(_01391_),
    .B(_01759_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand3_2 _09065_ (.A(_02194_),
    .B(_02195_),
    .C(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__xor2_4 _09066_ (.A(_01762_),
    .B(_02154_),
    .X(_02198_));
 sky130_fd_sc_hd__or2_1 _09067_ (.A(_02197_),
    .B(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__xor2_4 _09068_ (.A(_01763_),
    .B(_01767_),
    .X(_02200_));
 sky130_fd_sc_hd__or2_1 _09069_ (.A(_02199_),
    .B(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__nand4_1 _09070_ (.A(_01391_),
    .B(_01757_),
    .C(_01762_),
    .D(_01767_),
    .Y(_02202_));
 sky130_fd_sc_hd__o221a_2 _09071_ (.A1(_02137_),
    .A2(_02155_),
    .B1(_02202_),
    .B2(_02152_),
    .C1(_02157_),
    .X(_02203_));
 sky130_fd_sc_hd__xnor2_4 _09072_ (.A(_01764_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__or4_2 _09073_ (.A(_02197_),
    .B(_02198_),
    .C(_02200_),
    .D(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__xnor2_4 _09074_ (.A(_01769_),
    .B(_01772_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _09075_ (.A(_02205_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__xnor2_4 _09076_ (.A(_01770_),
    .B(_02160_),
    .Y(_02208_));
 sky130_fd_sc_hd__xnor2_4 _09077_ (.A(_01776_),
    .B(_01940_),
    .Y(_02209_));
 sky130_fd_sc_hd__or4bb_4 _09078_ (.A(_02205_),
    .B(_02206_),
    .C_N(_02208_),
    .D_N(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__nor2_1 _09079_ (.A(_02164_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__o21a_2 _09080_ (.A1(_01776_),
    .A2(_01941_),
    .B1(_02069_),
    .X(_02212_));
 sky130_fd_sc_hd__xnor2_4 _09081_ (.A(_02016_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__xor2_1 _09082_ (.A(_02016_),
    .B(_02212_),
    .X(_02214_));
 sky130_fd_sc_hd__o21bai_1 _09083_ (.A1(_01935_),
    .A2(_02014_),
    .B1_N(_02015_),
    .Y(_02215_));
 sky130_fd_sc_hd__a211o_1 _09084_ (.A1(_02136_),
    .A2(_02162_),
    .B1(_01936_),
    .C1(_02016_),
    .X(_02216_));
 sky130_fd_sc_hd__and2_1 _09085_ (.A(_02215_),
    .B(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__nand3_1 _09086_ (.A(_02064_),
    .B(_02215_),
    .C(_02216_),
    .Y(_02218_));
 sky130_fd_sc_hd__a21o_1 _09087_ (.A1(_02215_),
    .A2(_02216_),
    .B1(_02064_),
    .X(_02219_));
 sky130_fd_sc_hd__and2_2 _09088_ (.A(_02218_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__a2111o_1 _09089_ (.A1(_02218_),
    .A2(_02219_),
    .B1(_02164_),
    .C1(_02210_),
    .D1(_02214_),
    .X(_02221_));
 sky130_fd_sc_hd__and3_1 _09090_ (.A(_02065_),
    .B(_02070_),
    .C(_02095_),
    .X(_02222_));
 sky130_fd_sc_hd__a21oi_2 _09091_ (.A1(_02065_),
    .A2(_02070_),
    .B1(_02095_),
    .Y(_02223_));
 sky130_fd_sc_hd__or2_1 _09092_ (.A(_02222_),
    .B(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__o21bai_2 _09093_ (.A1(_02222_),
    .A2(_02223_),
    .B1_N(_02221_),
    .Y(_02225_));
 sky130_fd_sc_hd__o2bb2a_1 _09094_ (.A1_N(_02017_),
    .A2_N(_02062_),
    .B1(_02092_),
    .B2(_02093_),
    .X(_02226_));
 sky130_fd_sc_hd__a21o_1 _09095_ (.A1(_02092_),
    .A2(_02093_),
    .B1(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__o31ai_4 _09096_ (.A1(_02064_),
    .A2(_02095_),
    .A3(_02217_),
    .B1(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__xor2_4 _09097_ (.A(_02110_),
    .B(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__or4b_2 _09098_ (.A(_02016_),
    .B(_02064_),
    .C(_02095_),
    .D_N(_02110_),
    .X(_02230_));
 sky130_fd_sc_hd__o221ai_4 _09099_ (.A1(_02067_),
    .A2(_02111_),
    .B1(_02212_),
    .B2(_02230_),
    .C1(_02130_),
    .Y(_02231_));
 sky130_fd_sc_hd__xnor2_4 _09100_ (.A(_02122_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21bo_1 _09101_ (.A1(_02109_),
    .A2(_02119_),
    .B1_N(_02120_),
    .X(_02233_));
 sky130_fd_sc_hd__nand2_1 _09102_ (.A(_02110_),
    .B(_02121_),
    .Y(_02234_));
 sky130_fd_sc_hd__or4bb_1 _09103_ (.A(_02064_),
    .B(_02095_),
    .C_N(_02110_),
    .D_N(_02121_),
    .X(_02235_));
 sky130_fd_sc_hd__o221a_2 _09104_ (.A1(_02227_),
    .A2(_02234_),
    .B1(_02235_),
    .B2(_02217_),
    .C1(_02233_),
    .X(_02236_));
 sky130_fd_sc_hd__xor2_2 _09105_ (.A(_02127_),
    .B(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__nor4_1 _09106_ (.A(_02225_),
    .B(_02229_),
    .C(_02232_),
    .D(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__or2_1 _09107_ (.A(net150),
    .B(net3),
    .X(_02239_));
 sky130_fd_sc_hd__nand2_1 _09108_ (.A(_02133_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_1 _09109_ (.A(_06425_),
    .B(_06431_),
    .Y(_02241_));
 sky130_fd_sc_hd__or2_4 _09110_ (.A(_06425_),
    .B(_06431_),
    .X(_02242_));
 sky130_fd_sc_hd__o211a_1 _09111_ (.A1(_02133_),
    .A2(_02239_),
    .B1(_02240_),
    .C1(net202),
    .X(_02243_));
 sky130_fd_sc_hd__or4b_1 _09112_ (.A(net305),
    .B(_04487_),
    .C(_06409_),
    .D_N(_06407_),
    .X(_02244_));
 sky130_fd_sc_hd__or3b_1 _09113_ (.A(_06423_),
    .B(instruction[5]),
    .C_N(_06397_),
    .X(_02245_));
 sky130_fd_sc_hd__nor2_1 _09114_ (.A(net297),
    .B(_06449_),
    .Y(_02246_));
 sky130_fd_sc_hd__or2_4 _09115_ (.A(net297),
    .B(_06449_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(net301),
    .A1(reg1_val[30]),
    .S(net245),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _09117_ (.A0(net302),
    .A1(reg1_val[31]),
    .S(net245),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(_02248_),
    .A1(_02249_),
    .S(net216),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net245),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net245),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _09121_ (.A0(_02251_),
    .A1(_02252_),
    .S(net212),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(_02250_),
    .A1(_02253_),
    .S(net218),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _09123_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net244),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net244),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _09125_ (.A0(_02255_),
    .A1(_02256_),
    .S(net211),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _09126_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net243),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net243),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _09128_ (.A0(_02258_),
    .A1(_02259_),
    .S(net211),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _09129_ (.A0(_02257_),
    .A1(_02260_),
    .S(net218),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(_02254_),
    .A1(_02261_),
    .S(net220),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _09131_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net243),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net243),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _09133_ (.A0(_02263_),
    .A1(_02264_),
    .S(net211),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net243),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _09135_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net243),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(_02266_),
    .A1(_02267_),
    .S(net211),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _09137_ (.A0(_02265_),
    .A1(_02268_),
    .S(net217),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _09138_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net243),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _09139_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net243),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(_02270_),
    .A1(_02271_),
    .S(net212),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _09141_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(net243),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _09142_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(net243),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(_02273_),
    .A1(_02274_),
    .S(net211),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _09144_ (.A0(_02272_),
    .A1(_02275_),
    .S(net217),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _09145_ (.A0(_02269_),
    .A1(_02276_),
    .S(net220),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(_02262_),
    .A1(_02277_),
    .S(net222),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(reg1_val[24]),
    .A1(reg1_val[7]),
    .S(net244),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _09148_ (.A0(reg1_val[25]),
    .A1(reg1_val[6]),
    .S(net243),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _09149_ (.A0(_02279_),
    .A1(_02280_),
    .S(net212),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(reg1_val[26]),
    .A1(reg1_val[5]),
    .S(net245),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _09151_ (.A0(reg1_val[27]),
    .A1(reg1_val[4]),
    .S(net245),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _09152_ (.A0(_02282_),
    .A1(_02283_),
    .S(net212),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _09153_ (.A0(_02281_),
    .A1(_02284_),
    .S(net218),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(reg1_val[28]),
    .A1(reg1_val[3]),
    .S(net245),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(reg1_val[29]),
    .A1(reg1_val[2]),
    .S(net245),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(_02286_),
    .A1(_02287_),
    .S(net212),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(reg1_val[30]),
    .A1(net301),
    .S(net245),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(reg1_val[31]),
    .A1(net302),
    .S(net245),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(_02289_),
    .A1(_02290_),
    .S(net212),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(_02288_),
    .A1(_02291_),
    .S(net219),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(_02285_),
    .A1(_02292_),
    .S(net220),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(reg1_val[16]),
    .A1(reg1_val[15]),
    .S(net243),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(reg1_val[17]),
    .A1(reg1_val[14]),
    .S(net244),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(_02294_),
    .A1(_02295_),
    .S(net211),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _09165_ (.A0(reg1_val[18]),
    .A1(reg1_val[13]),
    .S(net244),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(reg1_val[19]),
    .A1(reg1_val[12]),
    .S(net243),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(_02297_),
    .A1(_02298_),
    .S(net211),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(_02296_),
    .A1(_02299_),
    .S(net217),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(reg1_val[20]),
    .A1(reg1_val[11]),
    .S(net243),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(reg1_val[21]),
    .A1(reg1_val[10]),
    .S(net243),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _09171_ (.A0(_02301_),
    .A1(_02302_),
    .S(net211),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(reg1_val[22]),
    .A1(reg1_val[9]),
    .S(net243),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _09173_ (.A0(reg1_val[23]),
    .A1(reg1_val[8]),
    .S(net244),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(_02304_),
    .A1(_02305_),
    .S(net211),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _09175_ (.A0(_02303_),
    .A1(_02306_),
    .S(net218),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(_02300_),
    .A1(_02307_),
    .S(net220),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _09177_ (.A0(_02293_),
    .A1(_02308_),
    .S(net224),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(_02278_),
    .A1(_02309_),
    .S(net226),
    .X(_02310_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(net302),
    .B(curr_PC[0]),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_1 _09180_ (.A(net302),
    .B(curr_PC[0]),
    .X(_02312_));
 sky130_fd_sc_hd__a21o_1 _09181_ (.A1(_02311_),
    .A2(_02312_),
    .B1(net229),
    .X(_02313_));
 sky130_fd_sc_hd__o211a_1 _09182_ (.A1(net260),
    .A2(_02310_),
    .B1(_02313_),
    .C1(net210),
    .X(_02314_));
 sky130_fd_sc_hd__nor2_4 _09183_ (.A(net304),
    .B(_06449_),
    .Y(_02315_));
 sky130_fd_sc_hd__or2_4 _09184_ (.A(net304),
    .B(_06449_),
    .X(_02316_));
 sky130_fd_sc_hd__nor2_8 _09185_ (.A(_06409_),
    .B(_06431_),
    .Y(_02317_));
 sky130_fd_sc_hd__or2_4 _09186_ (.A(_06409_),
    .B(_06431_),
    .X(_02318_));
 sky130_fd_sc_hd__nor3_1 _09187_ (.A(net306),
    .B(_04487_),
    .C(_06425_),
    .Y(_02319_));
 sky130_fd_sc_hd__or3_4 _09188_ (.A(net305),
    .B(_04487_),
    .C(_06425_),
    .X(_02320_));
 sky130_fd_sc_hd__a21oi_1 _09189_ (.A1(_02318_),
    .A2(net200),
    .B1(_06411_),
    .Y(_02321_));
 sky130_fd_sc_hd__and4bb_2 _09190_ (.A_N(instruction[3]),
    .B_N(net305),
    .C(instruction[5]),
    .D(instruction[4]),
    .X(_02322_));
 sky130_fd_sc_hd__or4b_4 _09191_ (.A(instruction[3]),
    .B(net305),
    .C(_04487_),
    .D_N(instruction[4]),
    .X(_02323_));
 sky130_fd_sc_hd__nor3_2 _09192_ (.A(net305),
    .B(instruction[5]),
    .C(_06409_),
    .Y(_02324_));
 sky130_fd_sc_hd__or3_2 _09193_ (.A(net305),
    .B(instruction[5]),
    .C(_06409_),
    .X(_02325_));
 sky130_fd_sc_hd__nor3_4 _09194_ (.A(net305),
    .B(_04487_),
    .C(_06423_),
    .Y(_02326_));
 sky130_fd_sc_hd__or3_4 _09195_ (.A(net305),
    .B(_04487_),
    .C(_06423_),
    .X(_02327_));
 sky130_fd_sc_hd__o21a_1 _09196_ (.A1(net242),
    .A2(net240),
    .B1(_06411_),
    .X(_02328_));
 sky130_fd_sc_hd__or3_1 _09197_ (.A(_02321_),
    .B(_02322_),
    .C(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__and4_2 _09198_ (.A(instruction[4]),
    .B(_04476_),
    .C(net306),
    .D(_04487_),
    .X(_02330_));
 sky130_fd_sc_hd__or3b_1 _09199_ (.A(instruction[3]),
    .B(_06431_),
    .C_N(instruction[4]),
    .X(_02331_));
 sky130_fd_sc_hd__and3_2 _09200_ (.A(net305),
    .B(_04487_),
    .C(_06424_),
    .X(_02332_));
 sky130_fd_sc_hd__or3b_4 _09201_ (.A(instruction[5]),
    .B(_06423_),
    .C_N(net305),
    .X(_02333_));
 sky130_fd_sc_hd__or2_1 _09202_ (.A(_06409_),
    .B(_06432_),
    .X(_02334_));
 sky130_fd_sc_hd__a2bb2o_1 _09203_ (.A1_N(net302),
    .A2_N(net237),
    .B1(_02330_),
    .B2(\div_res[0] ),
    .X(_02335_));
 sky130_fd_sc_hd__a221o_1 _09204_ (.A1(_06412_),
    .A2(_02329_),
    .B1(_02332_),
    .B2(\div_shifter[32] ),
    .C1(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__nor2_2 _09205_ (.A(_04552_),
    .B(net209),
    .Y(_02337_));
 sky130_fd_sc_hd__or2_4 _09206_ (.A(net225),
    .B(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(_02290_),
    .A1(_02337_),
    .S(net212),
    .X(_02339_));
 sky130_fd_sc_hd__o21ai_1 _09208_ (.A1(_06327_),
    .A2(_02337_),
    .B1(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__inv_2 _09209_ (.A(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__or2_1 _09210_ (.A(_06321_),
    .B(_02337_),
    .X(_02342_));
 sky130_fd_sc_hd__and2_1 _09211_ (.A(_02341_),
    .B(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__nor2_1 _09212_ (.A(net224),
    .B(_02337_),
    .Y(_02344_));
 sky130_fd_sc_hd__or2_2 _09213_ (.A(net224),
    .B(_02337_),
    .X(_02345_));
 sky130_fd_sc_hd__nand3_2 _09214_ (.A(_02338_),
    .B(_02343_),
    .C(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__inv_2 _09215_ (.A(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__a221o_1 _09216_ (.A1(_02310_),
    .A2(_02315_),
    .B1(_02347_),
    .B2(net245),
    .C1(_02336_),
    .X(_02348_));
 sky130_fd_sc_hd__nor2_1 _09217_ (.A(_02314_),
    .B(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__and4b_1 _09218_ (.A_N(_02243_),
    .B(_02244_),
    .C(_02245_),
    .D(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__o22a_2 _09219_ (.A1(net216),
    .A2(net251),
    .B1(_06457_),
    .B2(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__or2_1 _09220_ (.A(curr_PC[0]),
    .B(net253),
    .X(_02352_));
 sky130_fd_sc_hd__o21ai_4 _09221_ (.A1(net258),
    .A2(_02351_),
    .B1(_02352_),
    .Y(dest_val[0]));
 sky130_fd_sc_hd__or2_1 _09222_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .X(_02353_));
 sky130_fd_sc_hd__nand2_1 _09223_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .Y(_02354_));
 sky130_fd_sc_hd__a21o_1 _09224_ (.A1(_02133_),
    .A2(net3),
    .B1(net150),
    .X(_02355_));
 sky130_fd_sc_hd__a21oi_4 _09225_ (.A1(_00560_),
    .A2(_00751_),
    .B1(_00750_),
    .Y(_02356_));
 sky130_fd_sc_hd__nand2_2 _09226_ (.A(_00746_),
    .B(_00748_),
    .Y(_02357_));
 sky130_fd_sc_hd__a32o_1 _09227_ (.A1(_00647_),
    .A2(_00648_),
    .A3(_00657_),
    .B1(_00658_),
    .B2(_00638_),
    .X(_02358_));
 sky130_fd_sc_hd__o22a_1 _09228_ (.A1(net139),
    .A2(net28),
    .B1(net26),
    .B2(net147),
    .X(_02359_));
 sky130_fd_sc_hd__xnor2_2 _09229_ (.A(net68),
    .B(_02359_),
    .Y(_02360_));
 sky130_fd_sc_hd__o22a_1 _09230_ (.A1(net145),
    .A2(net30),
    .B1(net122),
    .B2(net31),
    .X(_02361_));
 sky130_fd_sc_hd__xor2_2 _09231_ (.A(net118),
    .B(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__xnor2_1 _09232_ (.A(_02360_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__o22a_1 _09233_ (.A1(net38),
    .A2(net143),
    .B1(net141),
    .B2(net36),
    .X(_02364_));
 sky130_fd_sc_hd__xnor2_1 _09234_ (.A(net119),
    .B(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__or2_1 _09235_ (.A(_02363_),
    .B(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(_02363_),
    .B(_02365_),
    .Y(_02367_));
 sky130_fd_sc_hd__nand2_1 _09237_ (.A(_02366_),
    .B(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__a21o_1 _09238_ (.A1(_00618_),
    .A2(_00627_),
    .B1(_00625_),
    .X(_02369_));
 sky130_fd_sc_hd__xor2_1 _09239_ (.A(_02368_),
    .B(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__and2b_1 _09240_ (.A_N(_02370_),
    .B(_02358_),
    .X(_02371_));
 sky130_fd_sc_hd__and2b_1 _09241_ (.A_N(_02358_),
    .B(_02370_),
    .X(_02372_));
 sky130_fd_sc_hd__nor2_2 _09242_ (.A(_02371_),
    .B(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__and2_1 _09243_ (.A(_00643_),
    .B(_00647_),
    .X(_02374_));
 sky130_fd_sc_hd__a21oi_2 _09244_ (.A1(_00694_),
    .A2(_00697_),
    .B1(_00693_),
    .Y(_02375_));
 sky130_fd_sc_hd__a21oi_2 _09245_ (.A1(_00634_),
    .A2(_00637_),
    .B1(_00633_),
    .Y(_02376_));
 sky130_fd_sc_hd__or2_1 _09246_ (.A(_02375_),
    .B(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__xor2_2 _09247_ (.A(_02375_),
    .B(_02376_),
    .X(_02378_));
 sky130_fd_sc_hd__nand2b_1 _09248_ (.A_N(_02374_),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__xnor2_2 _09249_ (.A(_02374_),
    .B(_02378_),
    .Y(_02380_));
 sky130_fd_sc_hd__o22a_1 _09250_ (.A1(net103),
    .A2(net78),
    .B1(net62),
    .B2(net107),
    .X(_02381_));
 sky130_fd_sc_hd__xnor2_1 _09251_ (.A(_00146_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand2_1 _09252_ (.A(_00180_),
    .B(_00271_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(_00190_),
    .B(_00284_),
    .Y(_02384_));
 sky130_fd_sc_hd__a21o_1 _09254_ (.A1(_02383_),
    .A2(_02384_),
    .B1(net184),
    .X(_02385_));
 sky130_fd_sc_hd__nand3_1 _09255_ (.A(net184),
    .B(_02383_),
    .C(_02384_),
    .Y(_02386_));
 sky130_fd_sc_hd__and3_1 _09256_ (.A(_02382_),
    .B(_02385_),
    .C(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__a21oi_2 _09257_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_02382_),
    .Y(_02388_));
 sky130_fd_sc_hd__nor2_1 _09258_ (.A(_02387_),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__o22a_1 _09259_ (.A1(net133),
    .A2(net65),
    .B1(net58),
    .B2(net135),
    .X(_02390_));
 sky130_fd_sc_hd__xnor2_2 _09260_ (.A(net186),
    .B(_02390_),
    .Y(_02391_));
 sky130_fd_sc_hd__xnor2_2 _09261_ (.A(_02389_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__o22a_1 _09262_ (.A1(net75),
    .A2(net98),
    .B1(net56),
    .B2(net72),
    .X(_02393_));
 sky130_fd_sc_hd__xnor2_1 _09263_ (.A(net129),
    .B(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__o22a_1 _09264_ (.A1(net104),
    .A2(net52),
    .B1(net50),
    .B2(net100),
    .X(_02395_));
 sky130_fd_sc_hd__xnor2_1 _09265_ (.A(net89),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2b_1 _09266_ (.A_N(_02394_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__xor2_1 _09267_ (.A(_02394_),
    .B(_02396_),
    .X(_02398_));
 sky130_fd_sc_hd__o22a_1 _09268_ (.A1(net69),
    .A2(net95),
    .B1(net54),
    .B2(net109),
    .X(_02399_));
 sky130_fd_sc_hd__xnor2_1 _09269_ (.A(net128),
    .B(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__or2_1 _09270_ (.A(_02398_),
    .B(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__nand2_1 _09271_ (.A(_02398_),
    .B(_02400_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(_02401_),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__o22a_2 _09273_ (.A1(net160),
    .A2(net18),
    .B1(net9),
    .B2(net162),
    .X(_02404_));
 sky130_fd_sc_hd__xnor2_4 _09274_ (.A(net204),
    .B(_02404_),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _09275_ (.A(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__o22a_2 _09276_ (.A1(net164),
    .A2(net24),
    .B1(net20),
    .B2(net166),
    .X(_02407_));
 sky130_fd_sc_hd__xnor2_4 _09277_ (.A(net207),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_1 _09278_ (.A(net249),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__xnor2_4 _09279_ (.A(_00255_),
    .B(_02408_),
    .Y(_02410_));
 sky130_fd_sc_hd__xnor2_4 _09280_ (.A(_02405_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__xnor2_2 _09281_ (.A(_02403_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__xor2_2 _09282_ (.A(_02392_),
    .B(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(_00224_),
    .B(net44),
    .Y(_02414_));
 sky130_fd_sc_hd__a21bo_1 _09284_ (.A1(_00651_),
    .A2(_00656_),
    .B1_N(_00655_),
    .X(_02415_));
 sky130_fd_sc_hd__o22a_1 _09285_ (.A1(net174),
    .A2(net16),
    .B1(net159),
    .B2(net7),
    .X(_02416_));
 sky130_fd_sc_hd__xnor2_2 _09286_ (.A(net40),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__and2b_1 _09287_ (.A_N(_02417_),
    .B(_02415_),
    .X(_02418_));
 sky130_fd_sc_hd__xnor2_2 _09288_ (.A(_02415_),
    .B(_02417_),
    .Y(_02419_));
 sky130_fd_sc_hd__xnor2_2 _09289_ (.A(_02414_),
    .B(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__and2_1 _09290_ (.A(_02413_),
    .B(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__xor2_2 _09291_ (.A(_02413_),
    .B(_02420_),
    .X(_02422_));
 sky130_fd_sc_hd__xnor2_1 _09292_ (.A(_02380_),
    .B(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__o21ai_2 _09293_ (.A1(_00604_),
    .A2(_00606_),
    .B1(_00602_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_1 _09294_ (.A(_06508_),
    .B(_00445_),
    .Y(_02425_));
 sky130_fd_sc_hd__or2_1 _09295_ (.A(net34),
    .B(net124),
    .X(_02426_));
 sky130_fd_sc_hd__and3_1 _09296_ (.A(net114),
    .B(_02425_),
    .C(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__a21oi_1 _09297_ (.A1(_02425_),
    .A2(_02426_),
    .B1(net114),
    .Y(_02428_));
 sky130_fd_sc_hd__o22a_1 _09298_ (.A1(net57),
    .A2(net49),
    .B1(net13),
    .B2(net93),
    .X(_02429_));
 sky130_fd_sc_hd__and2_1 _09299_ (.A(net85),
    .B(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__nor2_1 _09300_ (.A(net85),
    .B(_02429_),
    .Y(_02431_));
 sky130_fd_sc_hd__o22a_1 _09301_ (.A1(_02427_),
    .A2(_02428_),
    .B1(_02430_),
    .B2(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__or4_1 _09302_ (.A(_02427_),
    .B(_02428_),
    .C(_02430_),
    .D(_02431_),
    .X(_02433_));
 sky130_fd_sc_hd__and2b_1 _09303_ (.A_N(_02432_),
    .B(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__o22a_1 _09304_ (.A1(net91),
    .A2(net46),
    .B1(net12),
    .B2(net83),
    .X(_02435_));
 sky130_fd_sc_hd__xnor2_2 _09305_ (.A(net111),
    .B(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__xor2_2 _09306_ (.A(_02434_),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__a31o_2 _09307_ (.A1(net213),
    .A2(net44),
    .A3(_00670_),
    .B1(_00669_),
    .X(_02438_));
 sky130_fd_sc_hd__nand2_1 _09308_ (.A(_02437_),
    .B(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__xor2_2 _09309_ (.A(_02437_),
    .B(_02438_),
    .X(_02440_));
 sky130_fd_sc_hd__xnor2_1 _09310_ (.A(_02424_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__nor2_1 _09311_ (.A(_02423_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__nand2_1 _09312_ (.A(_02423_),
    .B(_02441_),
    .Y(_02443_));
 sky130_fd_sc_hd__and2b_1 _09313_ (.A_N(_02442_),
    .B(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__xor2_4 _09314_ (.A(_02373_),
    .B(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__a21o_1 _09315_ (.A1(_00617_),
    .A2(_00711_),
    .B1(_00710_),
    .X(_02446_));
 sky130_fd_sc_hd__nand2_2 _09316_ (.A(_00613_),
    .B(_00616_),
    .Y(_02447_));
 sky130_fd_sc_hd__a21o_2 _09317_ (.A1(_00628_),
    .A2(_00673_),
    .B1(_00672_),
    .X(_02448_));
 sky130_fd_sc_hd__a21o_1 _09318_ (.A1(_00684_),
    .A2(_00708_),
    .B1(_00707_),
    .X(_02449_));
 sky130_fd_sc_hd__nand2_1 _09319_ (.A(_02448_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__xor2_4 _09320_ (.A(_02448_),
    .B(_02449_),
    .X(_02451_));
 sky130_fd_sc_hd__xnor2_4 _09321_ (.A(_02447_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21oi_4 _09322_ (.A1(_00739_),
    .A2(_00743_),
    .B1(_00742_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_2 _09323_ (.A(_02452_),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__nand2b_1 _09324_ (.A_N(_02454_),
    .B(_02446_),
    .Y(_02455_));
 sky130_fd_sc_hd__xnor2_2 _09325_ (.A(_02446_),
    .B(_02454_),
    .Y(_02456_));
 sky130_fd_sc_hd__and2_1 _09326_ (.A(_02445_),
    .B(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__xor2_4 _09327_ (.A(_02445_),
    .B(_02456_),
    .X(_02458_));
 sky130_fd_sc_hd__xnor2_4 _09328_ (.A(_02357_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__or2_1 _09329_ (.A(_02356_),
    .B(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__and2_1 _09330_ (.A(_02356_),
    .B(_02459_),
    .X(_02461_));
 sky130_fd_sc_hd__xnor2_4 _09331_ (.A(_02356_),
    .B(_02459_),
    .Y(_02462_));
 sky130_fd_sc_hd__a21o_1 _09332_ (.A1(_00837_),
    .A2(_02126_),
    .B1(_00838_),
    .X(_02463_));
 sky130_fd_sc_hd__o31a_1 _09333_ (.A1(_00839_),
    .A2(_02127_),
    .A3(_02236_),
    .B1(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__xnor2_2 _09334_ (.A(_02462_),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__o21ai_1 _09335_ (.A1(_02355_),
    .A2(_02465_),
    .B1(net202),
    .Y(_02466_));
 sky130_fd_sc_hd__a21oi_1 _09336_ (.A1(_02355_),
    .A2(_02465_),
    .B1(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__o21ba_1 _09337_ (.A1(_06411_),
    .A2(net248),
    .B1_N(_01725_),
    .X(_02468_));
 sky130_fd_sc_hd__a41o_1 _09338_ (.A1(reg1_val[0]),
    .A2(net213),
    .A3(_00224_),
    .A4(_00255_),
    .B1(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__o21ai_1 _09339_ (.A1(_06411_),
    .A2(net150),
    .B1(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__o311a_1 _09340_ (.A1(_06411_),
    .A2(net150),
    .A3(_02469_),
    .B1(_02470_),
    .C1(_02317_),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(_02248_),
    .A1(_02251_),
    .S(net212),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(_02252_),
    .A1(_02255_),
    .S(net211),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(_02472_),
    .A1(_02473_),
    .S(net218),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(_02256_),
    .A1(_02258_),
    .S(net211),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(_02259_),
    .A1(_02263_),
    .S(net211),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(_02475_),
    .A1(_02476_),
    .S(net217),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _09347_ (.A0(_02474_),
    .A1(_02477_),
    .S(net220),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(_02264_),
    .A1(_02266_),
    .S(net211),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _09349_ (.A0(_02267_),
    .A1(_02270_),
    .S(net212),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(_02479_),
    .A1(_02480_),
    .S(net217),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(_02271_),
    .A1(_02273_),
    .S(net212),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(_02274_),
    .A1(_02294_),
    .S(net211),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _09353_ (.A0(_02482_),
    .A1(_02483_),
    .S(net217),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(_02481_),
    .A1(_02484_),
    .S(net221),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(_02478_),
    .A1(_02485_),
    .S(net222),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(_02280_),
    .A1(_02282_),
    .S(net212),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(_02283_),
    .A1(_02286_),
    .S(net212),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _09358_ (.A0(_02487_),
    .A1(_02488_),
    .S(net218),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(_02287_),
    .A1(_02289_),
    .S(net212),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(_02339_),
    .A1(_02490_),
    .S(_06327_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(_02489_),
    .A1(_02491_),
    .S(net220),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _09362_ (.A0(_02295_),
    .A1(_02297_),
    .S(net213),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _09363_ (.A0(_02298_),
    .A1(_02301_),
    .S(net211),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(_02493_),
    .A1(_02494_),
    .S(net217),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _09365_ (.A0(_02302_),
    .A1(_02304_),
    .S(net211),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _09366_ (.A0(_02279_),
    .A1(_02305_),
    .S(net216),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _09367_ (.A0(_02496_),
    .A1(_02497_),
    .S(net218),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _09368_ (.A0(_02495_),
    .A1(_02498_),
    .S(net220),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _09369_ (.A0(_02492_),
    .A1(_02499_),
    .S(net224),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(_02486_),
    .A1(_02500_),
    .S(net227),
    .X(_02501_));
 sky130_fd_sc_hd__nor2_1 _09371_ (.A(net301),
    .B(curr_PC[1]),
    .Y(_02502_));
 sky130_fd_sc_hd__and2_1 _09372_ (.A(net301),
    .B(curr_PC[1]),
    .X(_02503_));
 sky130_fd_sc_hd__nor2_1 _09373_ (.A(_02502_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__xnor2_1 _09374_ (.A(_02311_),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__or2_1 _09375_ (.A(net229),
    .B(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__o211a_1 _09376_ (.A1(net260),
    .A2(_02501_),
    .B1(_02506_),
    .C1(net210),
    .X(_02507_));
 sky130_fd_sc_hd__a21oi_1 _09377_ (.A1(\div_res[0] ),
    .A2(net153),
    .B1(\div_res[1] ),
    .Y(_02508_));
 sky130_fd_sc_hd__a31o_1 _09378_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .A3(net153),
    .B1(net198),
    .X(_02509_));
 sky130_fd_sc_hd__nor2_1 _09379_ (.A(_02508_),
    .B(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__xnor2_1 _09380_ (.A(_06330_),
    .B(_06334_),
    .Y(_02511_));
 sky130_fd_sc_hd__o21ai_1 _09381_ (.A1(net304),
    .A2(net216),
    .B1(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__or3_1 _09382_ (.A(net304),
    .B(net216),
    .C(_02511_),
    .X(_02513_));
 sky130_fd_sc_hd__nor2_1 _09383_ (.A(_06330_),
    .B(_02327_),
    .Y(_02514_));
 sky130_fd_sc_hd__and2_2 _09384_ (.A(divi1_sign),
    .B(net304),
    .X(_02515_));
 sky130_fd_sc_hd__and3_1 _09385_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .C(net235),
    .X(_02516_));
 sky130_fd_sc_hd__a21oi_1 _09386_ (.A1(\div_shifter[32] ),
    .A2(net235),
    .B1(\div_shifter[33] ),
    .Y(_02517_));
 sky130_fd_sc_hd__o32a_1 _09387_ (.A1(net238),
    .A2(_02516_),
    .A3(_02517_),
    .B1(net236),
    .B2(reg1_val[1]),
    .X(_02518_));
 sky130_fd_sc_hd__o21ai_1 _09388_ (.A1(_06327_),
    .A2(net251),
    .B1(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__a31o_1 _09389_ (.A1(net301),
    .A2(net219),
    .A3(net201),
    .B1(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__a211o_1 _09390_ (.A1(_06329_),
    .A2(net273),
    .B1(_02514_),
    .C1(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__a311o_1 _09391_ (.A1(_02324_),
    .A2(_02512_),
    .A3(_02513_),
    .B1(_02521_),
    .C1(_02510_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(_02291_),
    .A1(_02337_),
    .S(net219),
    .X(_02523_));
 sky130_fd_sc_hd__o21ai_1 _09393_ (.A1(net221),
    .A2(_02523_),
    .B1(_02342_),
    .Y(_02524_));
 sky130_fd_sc_hd__inv_2 _09394_ (.A(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__a21oi_1 _09395_ (.A1(net224),
    .A2(_02524_),
    .B1(_02344_),
    .Y(_02526_));
 sky130_fd_sc_hd__o21a_1 _09396_ (.A1(net227),
    .A2(_02526_),
    .B1(_02338_),
    .X(_02527_));
 sky130_fd_sc_hd__a221o_1 _09397_ (.A1(_02315_),
    .A2(_02501_),
    .B1(_02527_),
    .B2(net246),
    .C1(_02522_),
    .X(_02528_));
 sky130_fd_sc_hd__o41a_1 _09398_ (.A1(_02467_),
    .A2(_02471_),
    .A3(_02507_),
    .A4(_02528_),
    .B1(net255),
    .X(_02529_));
 sky130_fd_sc_hd__a31o_4 _09399_ (.A1(net258),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_02529_),
    .X(dest_val[1]));
 sky130_fd_sc_hd__and3_1 _09400_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .X(_02530_));
 sky130_fd_sc_hd__a21oi_1 _09401_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .B1(curr_PC[2]),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _09402_ (.A(_02530_),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__a31o_1 _09403_ (.A1(_02133_),
    .A2(net3),
    .A3(_02465_),
    .B1(net148),
    .X(_02533_));
 sky130_fd_sc_hd__a21oi_4 _09404_ (.A1(_02357_),
    .A2(_02458_),
    .B1(_02457_),
    .Y(_02534_));
 sky130_fd_sc_hd__o21ai_4 _09405_ (.A1(_02452_),
    .A2(_02453_),
    .B1(_02455_),
    .Y(_02535_));
 sky130_fd_sc_hd__a32o_2 _09406_ (.A1(_02401_),
    .A2(_02402_),
    .A3(_02411_),
    .B1(_02412_),
    .B2(_02392_),
    .X(_02536_));
 sky130_fd_sc_hd__o22a_1 _09407_ (.A1(net141),
    .A2(net28),
    .B1(net26),
    .B2(net139),
    .X(_02537_));
 sky130_fd_sc_hd__xnor2_1 _09408_ (.A(net68),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__o22a_1 _09409_ (.A1(net31),
    .A2(net124),
    .B1(net122),
    .B2(net30),
    .X(_02539_));
 sky130_fd_sc_hd__xor2_1 _09410_ (.A(net118),
    .B(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__or2_1 _09411_ (.A(_02538_),
    .B(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(_02538_),
    .B(_02540_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _09413_ (.A(_02541_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__o22a_1 _09414_ (.A1(net38),
    .A2(net145),
    .B1(net143),
    .B2(net36),
    .X(_02544_));
 sky130_fd_sc_hd__xnor2_1 _09415_ (.A(net119),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__xnor2_1 _09416_ (.A(_02543_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__a21o_1 _09417_ (.A1(_02377_),
    .A2(_02379_),
    .B1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__nand3_1 _09418_ (.A(_02377_),
    .B(_02379_),
    .C(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_2 _09419_ (.A(_02547_),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2b_1 _09420_ (.A_N(_02549_),
    .B(_02536_),
    .Y(_02550_));
 sky130_fd_sc_hd__xnor2_4 _09421_ (.A(_02536_),
    .B(_02549_),
    .Y(_02551_));
 sky130_fd_sc_hd__o21ai_2 _09422_ (.A1(_02360_),
    .A2(_02362_),
    .B1(_02366_),
    .Y(_02552_));
 sky130_fd_sc_hd__o22ai_1 _09423_ (.A1(net100),
    .A2(net49),
    .B1(net13),
    .B2(net57),
    .Y(_02553_));
 sky130_fd_sc_hd__xor2_1 _09424_ (.A(net86),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__o22a_1 _09425_ (.A1(net80),
    .A2(net83),
    .B1(net81),
    .B2(net34),
    .X(_02555_));
 sky130_fd_sc_hd__xnor2_1 _09426_ (.A(net114),
    .B(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__and2_1 _09427_ (.A(_02554_),
    .B(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__xor2_1 _09428_ (.A(_02554_),
    .B(_02556_),
    .X(_02558_));
 sky130_fd_sc_hd__o22a_1 _09429_ (.A1(net93),
    .A2(net46),
    .B1(net12),
    .B2(net91),
    .X(_02559_));
 sky130_fd_sc_hd__xnor2_1 _09430_ (.A(net111),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__and2_1 _09431_ (.A(_02558_),
    .B(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__nor2_1 _09432_ (.A(_02558_),
    .B(_02560_),
    .Y(_02562_));
 sky130_fd_sc_hd__nor2_1 _09433_ (.A(_02561_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__a31o_1 _09434_ (.A1(_00224_),
    .A2(net44),
    .A3(_02419_),
    .B1(_02418_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _09435_ (.A(_02563_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__xor2_1 _09436_ (.A(_02563_),
    .B(_02564_),
    .X(_02566_));
 sky130_fd_sc_hd__xnor2_1 _09437_ (.A(_02552_),
    .B(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__and2_1 _09438_ (.A(_02397_),
    .B(_02401_),
    .X(_02568_));
 sky130_fd_sc_hd__a21oi_1 _09439_ (.A1(_02433_),
    .A2(_02436_),
    .B1(_02432_),
    .Y(_02569_));
 sky130_fd_sc_hd__o21bai_2 _09440_ (.A1(_02388_),
    .A2(_02391_),
    .B1_N(_02387_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2b_1 _09441_ (.A_N(_02569_),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__xnor2_1 _09442_ (.A(_02569_),
    .B(_02570_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2b_1 _09443_ (.A_N(_02568_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_1 _09444_ (.A(_02568_),
    .B(_02572_),
    .Y(_02574_));
 sky130_fd_sc_hd__o22a_1 _09445_ (.A1(net107),
    .A2(net65),
    .B1(net62),
    .B2(net103),
    .X(_02575_));
 sky130_fd_sc_hd__xnor2_1 _09446_ (.A(net173),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__o22a_1 _09447_ (.A1(net170),
    .A2(_00264_),
    .B1(net22),
    .B2(net136),
    .X(_02577_));
 sky130_fd_sc_hd__xnor2_1 _09448_ (.A(net184),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__nor2_1 _09449_ (.A(_02576_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__xor2_1 _09450_ (.A(_02576_),
    .B(_02578_),
    .X(_02580_));
 sky130_fd_sc_hd__o22a_1 _09451_ (.A1(net135),
    .A2(net61),
    .B1(net58),
    .B2(net133),
    .X(_02581_));
 sky130_fd_sc_hd__xnor2_1 _09452_ (.A(net188),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__and2b_1 _09453_ (.A_N(_02582_),
    .B(_02580_),
    .X(_02583_));
 sky130_fd_sc_hd__and2b_1 _09454_ (.A_N(_02580_),
    .B(_02582_),
    .X(_02584_));
 sky130_fd_sc_hd__nor2_1 _09455_ (.A(_02583_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__o22a_1 _09456_ (.A1(net77),
    .A2(net98),
    .B1(net56),
    .B2(net75),
    .X(_02586_));
 sky130_fd_sc_hd__xnor2_1 _09457_ (.A(net129),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__o22a_1 _09458_ (.A1(net109),
    .A2(net52),
    .B1(net50),
    .B2(net105),
    .X(_02588_));
 sky130_fd_sc_hd__xnor2_1 _09459_ (.A(_00388_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__or2_1 _09460_ (.A(_02587_),
    .B(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__nand2_1 _09461_ (.A(_02587_),
    .B(_02589_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _09462_ (.A(_02590_),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__o22a_1 _09463_ (.A1(net72),
    .A2(net95),
    .B1(net54),
    .B2(net69),
    .X(_02593_));
 sky130_fd_sc_hd__xnor2_1 _09464_ (.A(net126),
    .B(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__xnor2_1 _09465_ (.A(_02592_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__o22a_1 _09466_ (.A1(net164),
    .A2(net20),
    .B1(net18),
    .B2(net166),
    .X(_02596_));
 sky130_fd_sc_hd__xnor2_2 _09467_ (.A(net207),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__nor2_1 _09468_ (.A(net249),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__xnor2_2 _09469_ (.A(_00255_),
    .B(_02597_),
    .Y(_02599_));
 sky130_fd_sc_hd__a21oi_1 _09470_ (.A1(_00287_),
    .A2(_00567_),
    .B1(net205),
    .Y(_02600_));
 sky130_fd_sc_hd__a31o_2 _09471_ (.A1(_00236_),
    .A2(_00279_),
    .A3(_00567_),
    .B1(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__xor2_2 _09472_ (.A(_02599_),
    .B(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__nand2b_1 _09473_ (.A_N(_02595_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__xnor2_1 _09474_ (.A(_02595_),
    .B(_02602_),
    .Y(_02604_));
 sky130_fd_sc_hd__xor2_1 _09475_ (.A(_02585_),
    .B(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__nor2_1 _09476_ (.A(net159),
    .B(net40),
    .Y(_02606_));
 sky130_fd_sc_hd__a21oi_2 _09477_ (.A1(_02406_),
    .A2(_02410_),
    .B1(_02409_),
    .Y(_02607_));
 sky130_fd_sc_hd__o22a_1 _09478_ (.A1(net147),
    .A2(net16),
    .B1(net7),
    .B2(net174),
    .X(_02608_));
 sky130_fd_sc_hd__xnor2_2 _09479_ (.A(net44),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__and2b_1 _09480_ (.A_N(_02607_),
    .B(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__xnor2_2 _09481_ (.A(_02607_),
    .B(_02609_),
    .Y(_02611_));
 sky130_fd_sc_hd__xor2_2 _09482_ (.A(_02606_),
    .B(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__and2_1 _09483_ (.A(_02605_),
    .B(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__xor2_1 _09484_ (.A(_02605_),
    .B(_02612_),
    .X(_02614_));
 sky130_fd_sc_hd__xnor2_1 _09485_ (.A(_02574_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__nor2_1 _09486_ (.A(_02567_),
    .B(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _09487_ (.A(_02567_),
    .B(_02615_),
    .Y(_02617_));
 sky130_fd_sc_hd__and2b_1 _09488_ (.A_N(_02616_),
    .B(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__xor2_4 _09489_ (.A(_02551_),
    .B(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__a21o_1 _09490_ (.A1(_02373_),
    .A2(_02443_),
    .B1(_02442_),
    .X(_02620_));
 sky130_fd_sc_hd__a31o_2 _09491_ (.A1(_02366_),
    .A2(_02367_),
    .A3(_02369_),
    .B1(_02371_),
    .X(_02621_));
 sky130_fd_sc_hd__a21oi_4 _09492_ (.A1(_02380_),
    .A2(_02422_),
    .B1(_02421_),
    .Y(_02622_));
 sky130_fd_sc_hd__a21boi_4 _09493_ (.A1(_02424_),
    .A2(_02440_),
    .B1_N(_02439_),
    .Y(_02623_));
 sky130_fd_sc_hd__nor2_1 _09494_ (.A(_02622_),
    .B(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__xor2_4 _09495_ (.A(_02622_),
    .B(_02623_),
    .X(_02625_));
 sky130_fd_sc_hd__xnor2_4 _09496_ (.A(_02621_),
    .B(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__a21boi_4 _09497_ (.A1(_02447_),
    .A2(_02451_),
    .B1_N(_02450_),
    .Y(_02627_));
 sky130_fd_sc_hd__xnor2_2 _09498_ (.A(_02626_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2b_1 _09499_ (.A_N(_02628_),
    .B(_02620_),
    .Y(_02629_));
 sky130_fd_sc_hd__xnor2_2 _09500_ (.A(_02620_),
    .B(_02628_),
    .Y(_02630_));
 sky130_fd_sc_hd__and2_1 _09501_ (.A(_02619_),
    .B(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__xor2_4 _09502_ (.A(_02619_),
    .B(_02630_),
    .X(_02632_));
 sky130_fd_sc_hd__xnor2_4 _09503_ (.A(_02535_),
    .B(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__or2_1 _09504_ (.A(_02534_),
    .B(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__and2_1 _09505_ (.A(_02534_),
    .B(_02633_),
    .X(_02635_));
 sky130_fd_sc_hd__xnor2_4 _09506_ (.A(_02534_),
    .B(_02633_),
    .Y(_02636_));
 sky130_fd_sc_hd__nor4_1 _09507_ (.A(_00839_),
    .B(_02122_),
    .C(_02127_),
    .D(_02462_),
    .Y(_02637_));
 sky130_fd_sc_hd__a21oi_2 _09508_ (.A1(_00837_),
    .A2(_02460_),
    .B1(_02461_),
    .Y(_02638_));
 sky130_fd_sc_hd__nor4_1 _09509_ (.A(_00839_),
    .B(_02125_),
    .C(_02129_),
    .D(_02462_),
    .Y(_02639_));
 sky130_fd_sc_hd__a211oi_4 _09510_ (.A1(_02231_),
    .A2(net5),
    .B1(_02638_),
    .C1(net4),
    .Y(_02640_));
 sky130_fd_sc_hd__xnor2_2 _09511_ (.A(_02636_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21ai_1 _09512_ (.A1(_02533_),
    .A2(_02641_),
    .B1(net202),
    .Y(_02642_));
 sky130_fd_sc_hd__a21oi_1 _09513_ (.A1(_02533_),
    .A2(_02641_),
    .B1(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(_01726_),
    .B(net157),
    .Y(_02644_));
 sky130_fd_sc_hd__mux2_1 _09515_ (.A0(_01724_),
    .A1(_02166_),
    .S(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__o21ai_1 _09516_ (.A1(net221),
    .A2(_02491_),
    .B1(_02342_),
    .Y(_02646_));
 sky130_fd_sc_hd__inv_2 _09517_ (.A(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__a21oi_1 _09518_ (.A1(net224),
    .A2(_02646_),
    .B1(_02344_),
    .Y(_02648_));
 sky130_fd_sc_hd__o21a_1 _09519_ (.A1(net227),
    .A2(_02648_),
    .B1(_02338_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _09520_ (.A0(_02253_),
    .A1(_02257_),
    .S(net218),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _09521_ (.A0(_02260_),
    .A1(_02265_),
    .S(net217),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _09522_ (.A0(_02650_),
    .A1(_02651_),
    .S(net220),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _09523_ (.A0(_02268_),
    .A1(_02272_),
    .S(net217),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _09524_ (.A0(_02275_),
    .A1(_02296_),
    .S(net217),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _09525_ (.A0(_02653_),
    .A1(_02654_),
    .S(net220),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _09526_ (.A0(_02652_),
    .A1(_02655_),
    .S(net222),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _09527_ (.A0(_02284_),
    .A1(_02288_),
    .S(net218),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _09528_ (.A0(_02523_),
    .A1(_02657_),
    .S(_06321_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(_02299_),
    .A1(_02303_),
    .S(net217),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _09530_ (.A0(_02281_),
    .A1(_02306_),
    .S(_06327_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _09531_ (.A0(_02659_),
    .A1(_02660_),
    .S(net221),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _09532_ (.A0(_02658_),
    .A1(_02661_),
    .S(net224),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _09533_ (.A0(_02656_),
    .A1(_02662_),
    .S(net227),
    .X(_02663_));
 sky130_fd_sc_hd__o21ba_1 _09534_ (.A1(_02311_),
    .A2(_02502_),
    .B1_N(_02503_),
    .X(_02664_));
 sky130_fd_sc_hd__nor2_1 _09535_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _09536_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02666_));
 sky130_fd_sc_hd__and2b_1 _09537_ (.A_N(_02665_),
    .B(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__xnor2_1 _09538_ (.A(_02664_),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__or2_1 _09539_ (.A(net229),
    .B(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__or2_1 _09540_ (.A(\div_res[1] ),
    .B(\div_res[0] ),
    .X(_02670_));
 sky130_fd_sc_hd__a21oi_1 _09541_ (.A1(net153),
    .A2(_02670_),
    .B1(\div_res[2] ),
    .Y(_02671_));
 sky130_fd_sc_hd__a31o_1 _09542_ (.A1(\div_res[2] ),
    .A2(net153),
    .A3(_02670_),
    .B1(net198),
    .X(_02672_));
 sky130_fd_sc_hd__a22o_1 _09543_ (.A1(net301),
    .A2(net219),
    .B1(net213),
    .B2(net302),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_1 _09544_ (.A(_06329_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__mux2_1 _09545_ (.A0(_06336_),
    .A1(_02674_),
    .S(net298),
    .X(_02675_));
 sky130_fd_sc_hd__a21oi_1 _09546_ (.A1(_06325_),
    .A2(_02675_),
    .B1(net241),
    .Y(_02676_));
 sky130_fd_sc_hd__o21ai_1 _09547_ (.A1(_06325_),
    .A2(_02675_),
    .B1(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__o21a_1 _09548_ (.A1(\div_shifter[33] ),
    .A2(\div_shifter[32] ),
    .B1(net235),
    .X(_02678_));
 sky130_fd_sc_hd__xnor2_1 _09549_ (.A(\div_shifter[34] ),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__o22a_1 _09550_ (.A1(reg1_val[2]),
    .A2(net237),
    .B1(_02679_),
    .B2(_02333_),
    .X(_02680_));
 sky130_fd_sc_hd__mux2_1 _09551_ (.A0(_02649_),
    .A1(_02663_),
    .S(net298),
    .X(_02681_));
 sky130_fd_sc_hd__o211a_1 _09552_ (.A1(net260),
    .A2(_02663_),
    .B1(_02669_),
    .C1(net210),
    .X(_02682_));
 sky130_fd_sc_hd__o221a_1 _09553_ (.A1(_06321_),
    .A2(net251),
    .B1(_02323_),
    .B2(_06323_),
    .C1(_02680_),
    .X(_02683_));
 sky130_fd_sc_hd__o221a_1 _09554_ (.A1(_06324_),
    .A2(net200),
    .B1(_02327_),
    .B2(_06325_),
    .C1(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__o211ai_1 _09555_ (.A1(_02671_),
    .A2(_02672_),
    .B1(_02677_),
    .C1(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__a211o_1 _09556_ (.A1(_06448_),
    .A2(_02681_),
    .B1(_02682_),
    .C1(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__a211o_1 _09557_ (.A1(_02317_),
    .A2(_02645_),
    .B1(_02686_),
    .C1(_02643_),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_8 _09558_ (.A0(_02532_),
    .A1(_02687_),
    .S(net253),
    .X(dest_val[2]));
 sky130_fd_sc_hd__and4_1 _09559_ (.A(_02133_),
    .B(net3),
    .C(_02465_),
    .D(_02641_),
    .X(_02688_));
 sky130_fd_sc_hd__or2_1 _09560_ (.A(net148),
    .B(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__a21oi_4 _09561_ (.A1(_02535_),
    .A2(_02632_),
    .B1(_02631_),
    .Y(_02690_));
 sky130_fd_sc_hd__o21ai_4 _09562_ (.A1(_02626_),
    .A2(_02627_),
    .B1(_02629_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21bo_2 _09563_ (.A1(_02585_),
    .A2(_02604_),
    .B1_N(_02603_),
    .X(_02692_));
 sky130_fd_sc_hd__o22a_1 _09564_ (.A1(net143),
    .A2(net28),
    .B1(net26),
    .B2(net141),
    .X(_02693_));
 sky130_fd_sc_hd__xnor2_1 _09565_ (.A(net68),
    .B(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__o22a_1 _09566_ (.A1(net31),
    .A2(net81),
    .B1(net124),
    .B2(net30),
    .X(_02695_));
 sky130_fd_sc_hd__xor2_1 _09567_ (.A(net118),
    .B(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__or2_1 _09568_ (.A(_02694_),
    .B(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__nand2_1 _09569_ (.A(_02694_),
    .B(_02696_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _09570_ (.A(_02697_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__o22a_1 _09571_ (.A1(net36),
    .A2(net145),
    .B1(net122),
    .B2(net38),
    .X(_02700_));
 sky130_fd_sc_hd__xnor2_1 _09572_ (.A(net119),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__xnor2_1 _09573_ (.A(_02699_),
    .B(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__a21oi_1 _09574_ (.A1(_02571_),
    .A2(_02573_),
    .B1(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__and3_1 _09575_ (.A(_02571_),
    .B(_02573_),
    .C(_02702_),
    .X(_02704_));
 sky130_fd_sc_hd__nor2_2 _09576_ (.A(_02703_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__xor2_4 _09577_ (.A(_02692_),
    .B(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__o21ai_2 _09578_ (.A1(_02543_),
    .A2(_02545_),
    .B1(_02541_),
    .Y(_02707_));
 sky130_fd_sc_hd__o22a_1 _09579_ (.A1(net105),
    .A2(net49),
    .B1(net14),
    .B2(net100),
    .X(_02708_));
 sky130_fd_sc_hd__xnor2_1 _09580_ (.A(net86),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__o22a_1 _09581_ (.A1(net80),
    .A2(net91),
    .B1(net83),
    .B2(net34),
    .X(_02710_));
 sky130_fd_sc_hd__xnor2_1 _09582_ (.A(net114),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__and2_1 _09583_ (.A(_02709_),
    .B(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__xnor2_1 _09584_ (.A(_02709_),
    .B(_02711_),
    .Y(_02713_));
 sky130_fd_sc_hd__o22a_1 _09585_ (.A1(net57),
    .A2(net46),
    .B1(net12),
    .B2(net93),
    .X(_02714_));
 sky130_fd_sc_hd__xnor2_1 _09586_ (.A(net110),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__nor2_1 _09587_ (.A(_02713_),
    .B(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__and2_1 _09588_ (.A(_02713_),
    .B(_02715_),
    .X(_02717_));
 sky130_fd_sc_hd__nor2_1 _09589_ (.A(_02716_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21o_1 _09590_ (.A1(_02606_),
    .A2(_02611_),
    .B1(_02610_),
    .X(_02719_));
 sky130_fd_sc_hd__nand2_1 _09591_ (.A(_02718_),
    .B(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__xor2_2 _09592_ (.A(_02718_),
    .B(_02719_),
    .X(_02721_));
 sky130_fd_sc_hd__xor2_1 _09593_ (.A(_02707_),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__o21ai_2 _09594_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02590_),
    .Y(_02723_));
 sky130_fd_sc_hd__o22ai_2 _09595_ (.A1(_02557_),
    .A2(_02561_),
    .B1(_02579_),
    .B2(_02583_),
    .Y(_02724_));
 sky130_fd_sc_hd__or4_2 _09596_ (.A(_02557_),
    .B(_02561_),
    .C(_02579_),
    .D(_02583_),
    .X(_02725_));
 sky130_fd_sc_hd__and3_1 _09597_ (.A(_02723_),
    .B(_02724_),
    .C(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__a21oi_1 _09598_ (.A1(_02724_),
    .A2(_02725_),
    .B1(_02723_),
    .Y(_02727_));
 sky130_fd_sc_hd__or2_1 _09599_ (.A(_02726_),
    .B(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_06491_),
    .B(net44),
    .Y(_02729_));
 sky130_fd_sc_hd__a21oi_2 _09601_ (.A1(_02599_),
    .A2(_02601_),
    .B1(_02598_),
    .Y(_02730_));
 sky130_fd_sc_hd__o22a_1 _09602_ (.A1(net139),
    .A2(net16),
    .B1(net7),
    .B2(net147),
    .X(_02731_));
 sky130_fd_sc_hd__xnor2_2 _09603_ (.A(net43),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__and2b_1 _09604_ (.A_N(_02730_),
    .B(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__xnor2_2 _09605_ (.A(_02730_),
    .B(_02732_),
    .Y(_02734_));
 sky130_fd_sc_hd__xnor2_2 _09606_ (.A(_02729_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__o22a_1 _09607_ (.A1(net103),
    .A2(net65),
    .B1(net58),
    .B2(net107),
    .X(_02736_));
 sky130_fd_sc_hd__xnor2_1 _09608_ (.A(net173),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__o22a_1 _09609_ (.A1(net136),
    .A2(_00264_),
    .B1(net20),
    .B2(net170),
    .X(_02738_));
 sky130_fd_sc_hd__xnor2_1 _09610_ (.A(net184),
    .B(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__nor2_1 _09611_ (.A(_02737_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__xor2_1 _09612_ (.A(_02737_),
    .B(_02739_),
    .X(_02741_));
 sky130_fd_sc_hd__o22a_1 _09613_ (.A1(net135),
    .A2(net22),
    .B1(net61),
    .B2(net133),
    .X(_02742_));
 sky130_fd_sc_hd__xnor2_1 _09614_ (.A(net186),
    .B(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__and2b_1 _09615_ (.A_N(_02743_),
    .B(_02741_),
    .X(_02744_));
 sky130_fd_sc_hd__and2b_1 _09616_ (.A_N(_02741_),
    .B(_02743_),
    .X(_02745_));
 sky130_fd_sc_hd__nor2_1 _09617_ (.A(_02744_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__o22a_1 _09618_ (.A1(net164),
    .A2(net18),
    .B1(net9),
    .B2(net166),
    .X(_02747_));
 sky130_fd_sc_hd__xnor2_2 _09619_ (.A(net206),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__nor2_1 _09620_ (.A(_00255_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__xnor2_2 _09621_ (.A(net249),
    .B(_02748_),
    .Y(_02750_));
 sky130_fd_sc_hd__xnor2_2 _09622_ (.A(net204),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__o22a_1 _09623_ (.A1(net62),
    .A2(net98),
    .B1(net56),
    .B2(net77),
    .X(_02752_));
 sky130_fd_sc_hd__xnor2_1 _09624_ (.A(net129),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__o22a_1 _09625_ (.A1(net69),
    .A2(net53),
    .B1(net51),
    .B2(net109),
    .X(_02754_));
 sky130_fd_sc_hd__xnor2_1 _09626_ (.A(_00388_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__or2_1 _09627_ (.A(_02753_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(_02753_),
    .B(_02755_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_2 _09629_ (.A(_02756_),
    .B(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__o22a_1 _09630_ (.A1(net75),
    .A2(net96),
    .B1(net55),
    .B2(net72),
    .X(_02759_));
 sky130_fd_sc_hd__xnor2_2 _09631_ (.A(net126),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__xnor2_1 _09632_ (.A(_02758_),
    .B(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__nor2_1 _09633_ (.A(_02751_),
    .B(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__xor2_1 _09634_ (.A(_02751_),
    .B(_02761_),
    .X(_02763_));
 sky130_fd_sc_hd__xor2_1 _09635_ (.A(_02746_),
    .B(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__nand2_1 _09636_ (.A(_02735_),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__xnor2_1 _09637_ (.A(_02735_),
    .B(_02764_),
    .Y(_02766_));
 sky130_fd_sc_hd__xor2_1 _09638_ (.A(_02728_),
    .B(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_02722_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__or2_1 _09640_ (.A(_02722_),
    .B(_02767_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_2 _09641_ (.A(_02768_),
    .B(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__xor2_4 _09642_ (.A(_02706_),
    .B(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__a21o_1 _09643_ (.A1(_02551_),
    .A2(_02617_),
    .B1(_02616_),
    .X(_02772_));
 sky130_fd_sc_hd__a21o_1 _09644_ (.A1(_02621_),
    .A2(_02625_),
    .B1(_02624_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_2 _09645_ (.A(_02547_),
    .B(_02550_),
    .Y(_02774_));
 sky130_fd_sc_hd__a21bo_2 _09646_ (.A1(_02552_),
    .A2(_02566_),
    .B1_N(_02565_),
    .X(_02775_));
 sky130_fd_sc_hd__a21o_2 _09647_ (.A1(_02574_),
    .A2(_02614_),
    .B1(_02613_),
    .X(_02776_));
 sky130_fd_sc_hd__nand2_1 _09648_ (.A(_02775_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__xor2_4 _09649_ (.A(_02775_),
    .B(_02776_),
    .X(_02778_));
 sky130_fd_sc_hd__xor2_2 _09650_ (.A(_02774_),
    .B(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__xnor2_2 _09651_ (.A(_02773_),
    .B(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2b_1 _09652_ (.A_N(_02780_),
    .B(_02772_),
    .Y(_02781_));
 sky130_fd_sc_hd__xnor2_2 _09653_ (.A(_02772_),
    .B(_02780_),
    .Y(_02782_));
 sky130_fd_sc_hd__and2_1 _09654_ (.A(_02771_),
    .B(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__xor2_4 _09655_ (.A(_02771_),
    .B(_02782_),
    .X(_02784_));
 sky130_fd_sc_hd__xnor2_4 _09656_ (.A(_02691_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__or2_1 _09657_ (.A(_02690_),
    .B(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__and2_1 _09658_ (.A(_02690_),
    .B(_02785_),
    .X(_02787_));
 sky130_fd_sc_hd__xnor2_4 _09659_ (.A(_02690_),
    .B(_02785_),
    .Y(_02788_));
 sky130_fd_sc_hd__or4_2 _09660_ (.A(_00839_),
    .B(_02127_),
    .C(_02462_),
    .D(_02636_),
    .X(_02789_));
 sky130_fd_sc_hd__a21o_1 _09661_ (.A1(_02460_),
    .A2(_02634_),
    .B1(_02635_),
    .X(_02790_));
 sky130_fd_sc_hd__a2111o_1 _09662_ (.A1(_00837_),
    .A2(_02126_),
    .B1(_02462_),
    .C1(_02636_),
    .D1(_00838_),
    .X(_02791_));
 sky130_fd_sc_hd__o211a_2 _09663_ (.A1(_02236_),
    .A2(_02789_),
    .B1(_02790_),
    .C1(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__xnor2_4 _09664_ (.A(_02788_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__or2_1 _09665_ (.A(_02689_),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_1 _09666_ (.A(_02689_),
    .B(_02793_),
    .Y(_02795_));
 sky130_fd_sc_hd__o21ai_1 _09667_ (.A1(net148),
    .A2(_02167_),
    .B1(_02169_),
    .Y(_02796_));
 sky130_fd_sc_hd__or3_1 _09668_ (.A(net148),
    .B(_02167_),
    .C(_02169_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(_02473_),
    .A1(_02475_),
    .S(net217),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(_02476_),
    .A1(_02479_),
    .S(net217),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(_02798_),
    .A1(_02799_),
    .S(net220),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _09672_ (.A0(_02480_),
    .A1(_02482_),
    .S(net217),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _09673_ (.A0(_02483_),
    .A1(_02493_),
    .S(net217),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _09674_ (.A0(_02801_),
    .A1(_02802_),
    .S(net220),
    .X(_02803_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(_02800_),
    .A1(_02803_),
    .S(net222),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _09676_ (.A0(_02488_),
    .A1(_02490_),
    .S(net218),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(_02341_),
    .A1(_02805_),
    .S(_06321_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _09678_ (.A0(_02494_),
    .A1(_02496_),
    .S(net217),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(_02487_),
    .A1(_02497_),
    .S(_06327_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _09680_ (.A0(_02807_),
    .A1(_02808_),
    .S(net220),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(_02806_),
    .A1(_02809_),
    .S(net224),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_2 _09682_ (.A0(_02804_),
    .A1(_02810_),
    .S(net226),
    .X(_02811_));
 sky130_fd_sc_hd__o21a_1 _09683_ (.A1(_02664_),
    .A2(_02665_),
    .B1(_02666_),
    .X(_02812_));
 sky130_fd_sc_hd__nor2_1 _09684_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_1 _09685_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02814_));
 sky130_fd_sc_hd__and2b_1 _09686_ (.A_N(_02813_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__o21ai_1 _09687_ (.A1(_02812_),
    .A2(_02815_),
    .B1(net260),
    .Y(_02816_));
 sky130_fd_sc_hd__a21o_1 _09688_ (.A1(_02812_),
    .A2(_02815_),
    .B1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__o211a_1 _09689_ (.A1(net260),
    .A2(_02811_),
    .B1(_02817_),
    .C1(net210),
    .X(_02818_));
 sky130_fd_sc_hd__o21a_1 _09690_ (.A1(net221),
    .A2(_02292_),
    .B1(_02342_),
    .X(_02819_));
 sky130_fd_sc_hd__o21a_1 _09691_ (.A1(net223),
    .A2(_02819_),
    .B1(_02345_),
    .X(_02820_));
 sky130_fd_sc_hd__o21a_1 _09692_ (.A1(net227),
    .A2(_02820_),
    .B1(_02338_),
    .X(_02821_));
 sky130_fd_sc_hd__a21boi_1 _09693_ (.A1(_06329_),
    .A2(_02673_),
    .B1_N(_06324_),
    .Y(_02822_));
 sky130_fd_sc_hd__nor2_1 _09694_ (.A(_06323_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__mux2_1 _09695_ (.A0(_06338_),
    .A1(_02823_),
    .S(net298),
    .X(_02824_));
 sky130_fd_sc_hd__o21ai_1 _09696_ (.A1(_06318_),
    .A2(_02824_),
    .B1(_02324_),
    .Y(_02825_));
 sky130_fd_sc_hd__a21oi_1 _09697_ (.A1(_06318_),
    .A2(_02824_),
    .B1(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__o31a_1 _09698_ (.A1(\div_res[2] ),
    .A2(\div_res[1] ),
    .A3(\div_res[0] ),
    .B1(net152),
    .X(_02827_));
 sky130_fd_sc_hd__a21oi_1 _09699_ (.A1(\div_res[3] ),
    .A2(_02827_),
    .B1(net198),
    .Y(_02828_));
 sky130_fd_sc_hd__o21a_1 _09700_ (.A1(\div_res[3] ),
    .A2(_02827_),
    .B1(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__or3_1 _09701_ (.A(\div_shifter[34] ),
    .B(\div_shifter[33] ),
    .C(\div_shifter[32] ),
    .X(_02830_));
 sky130_fd_sc_hd__a21oi_1 _09702_ (.A1(net234),
    .A2(_02830_),
    .B1(\div_shifter[35] ),
    .Y(_02831_));
 sky130_fd_sc_hd__and3_1 _09703_ (.A(\div_shifter[35] ),
    .B(net234),
    .C(_02830_),
    .X(_02832_));
 sky130_fd_sc_hd__o32a_1 _09704_ (.A1(net238),
    .A2(_02831_),
    .A3(_02832_),
    .B1(net236),
    .B2(reg1_val[3]),
    .X(_02833_));
 sky130_fd_sc_hd__o221a_1 _09705_ (.A1(_06314_),
    .A2(net251),
    .B1(net200),
    .B2(_06317_),
    .C1(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__o221a_1 _09706_ (.A1(_06316_),
    .A2(_02323_),
    .B1(_02327_),
    .B2(_06319_),
    .C1(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__or4b_1 _09707_ (.A(_02818_),
    .B(_02826_),
    .C(_02829_),
    .D_N(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__a221o_1 _09708_ (.A1(_02315_),
    .A2(_02811_),
    .B1(_02821_),
    .B2(net245),
    .C1(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__a31o_1 _09709_ (.A1(_02317_),
    .A2(_02796_),
    .A3(_02797_),
    .B1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__a31o_1 _09710_ (.A1(net202),
    .A2(_02794_),
    .A3(_02795_),
    .B1(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__or2_1 _09711_ (.A(curr_PC[3]),
    .B(_02530_),
    .X(_02840_));
 sky130_fd_sc_hd__and2_1 _09712_ (.A(curr_PC[3]),
    .B(_02530_),
    .X(_02841_));
 sky130_fd_sc_hd__nor2_1 _09713_ (.A(net253),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__a22o_4 _09714_ (.A1(net253),
    .A2(_02839_),
    .B1(_02840_),
    .B2(_02842_),
    .X(dest_val[3]));
 sky130_fd_sc_hd__and2_1 _09715_ (.A(_02688_),
    .B(_02793_),
    .X(_02843_));
 sky130_fd_sc_hd__or2_1 _09716_ (.A(net148),
    .B(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__a21oi_4 _09717_ (.A1(_02691_),
    .A2(_02784_),
    .B1(_02783_),
    .Y(_02845_));
 sky130_fd_sc_hd__a21bo_2 _09718_ (.A1(_02773_),
    .A2(_02779_),
    .B1_N(_02781_),
    .X(_02846_));
 sky130_fd_sc_hd__a21o_2 _09719_ (.A1(_02746_),
    .A2(_02763_),
    .B1(_02762_),
    .X(_02847_));
 sky130_fd_sc_hd__o22a_1 _09720_ (.A1(net145),
    .A2(net28),
    .B1(net26),
    .B2(net143),
    .X(_02848_));
 sky130_fd_sc_hd__xnor2_1 _09721_ (.A(net68),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__o22a_1 _09722_ (.A1(net31),
    .A2(net83),
    .B1(net81),
    .B2(net30),
    .X(_02850_));
 sky130_fd_sc_hd__xor2_1 _09723_ (.A(net118),
    .B(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__or2_1 _09724_ (.A(_02849_),
    .B(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__nand2_1 _09725_ (.A(_02849_),
    .B(_02851_),
    .Y(_02853_));
 sky130_fd_sc_hd__nand2_2 _09726_ (.A(_02852_),
    .B(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__o22a_2 _09727_ (.A1(net38),
    .A2(net124),
    .B1(net122),
    .B2(net36),
    .X(_02855_));
 sky130_fd_sc_hd__xnor2_4 _09728_ (.A(net119),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__xnor2_4 _09729_ (.A(_02854_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__a21boi_4 _09730_ (.A1(_02723_),
    .A2(_02725_),
    .B1_N(_02724_),
    .Y(_02858_));
 sky130_fd_sc_hd__xnor2_4 _09731_ (.A(_02857_),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2b_1 _09732_ (.A_N(_02859_),
    .B(_02847_),
    .Y(_02860_));
 sky130_fd_sc_hd__xnor2_4 _09733_ (.A(_02847_),
    .B(_02859_),
    .Y(_02861_));
 sky130_fd_sc_hd__o21ai_4 _09734_ (.A1(_02758_),
    .A2(_02760_),
    .B1(_02756_),
    .Y(_02862_));
 sky130_fd_sc_hd__o22a_1 _09735_ (.A1(_02712_),
    .A2(_02716_),
    .B1(_02740_),
    .B2(_02744_),
    .X(_02863_));
 sky130_fd_sc_hd__or4_2 _09736_ (.A(_02712_),
    .B(_02716_),
    .C(_02740_),
    .D(_02744_),
    .X(_02864_));
 sky130_fd_sc_hd__and2b_1 _09737_ (.A_N(_02863_),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__xnor2_2 _09738_ (.A(_02862_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__o22a_1 _09739_ (.A1(net107),
    .A2(net61),
    .B1(net58),
    .B2(net103),
    .X(_02867_));
 sky130_fd_sc_hd__xnor2_1 _09740_ (.A(net173),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__o22a_1 _09741_ (.A1(net65),
    .A2(net98),
    .B1(net56),
    .B2(net62),
    .X(_02869_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(_00298_),
    .B(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__o22a_1 _09743_ (.A1(net135),
    .A2(_00264_),
    .B1(net22),
    .B2(net133),
    .X(_02871_));
 sky130_fd_sc_hd__xnor2_1 _09744_ (.A(net186),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__nor2_1 _09745_ (.A(_02870_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__xnor2_1 _09746_ (.A(_02870_),
    .B(_02872_),
    .Y(_02874_));
 sky130_fd_sc_hd__nor2_2 _09747_ (.A(_02868_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__and2_1 _09748_ (.A(_02868_),
    .B(_02874_),
    .X(_02876_));
 sky130_fd_sc_hd__nor2_1 _09749_ (.A(_02875_),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__o22a_1 _09750_ (.A1(net77),
    .A2(net95),
    .B1(net54),
    .B2(net75),
    .X(_02878_));
 sky130_fd_sc_hd__xnor2_1 _09751_ (.A(net126),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__or2_1 _09752_ (.A(net109),
    .B(net49),
    .X(_02880_));
 sky130_fd_sc_hd__a21o_1 _09753_ (.A1(_00438_),
    .A2(_00439_),
    .B1(net105),
    .X(_02881_));
 sky130_fd_sc_hd__nand3_1 _09754_ (.A(net85),
    .B(_02880_),
    .C(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__a21o_1 _09755_ (.A1(_02880_),
    .A2(_02881_),
    .B1(net85),
    .X(_02883_));
 sky130_fd_sc_hd__a21oi_1 _09756_ (.A1(_02882_),
    .A2(_02883_),
    .B1(_02879_),
    .Y(_02884_));
 sky130_fd_sc_hd__and3_1 _09757_ (.A(_02879_),
    .B(_02882_),
    .C(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__or2_1 _09758_ (.A(_02884_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__o22a_1 _09759_ (.A1(net72),
    .A2(net53),
    .B1(net51),
    .B2(net69),
    .X(_02887_));
 sky130_fd_sc_hd__xnor2_2 _09760_ (.A(_00388_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__xor2_2 _09761_ (.A(_02886_),
    .B(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__o22a_1 _09762_ (.A1(net136),
    .A2(_00349_),
    .B1(net18),
    .B2(net170),
    .X(_02890_));
 sky130_fd_sc_hd__xnor2_1 _09763_ (.A(net183),
    .B(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__nor2_1 _09764_ (.A(_00239_),
    .B(net9),
    .Y(_02892_));
 sky130_fd_sc_hd__o22ai_2 _09765_ (.A1(_00247_),
    .A2(net9),
    .B1(_02892_),
    .B2(net206),
    .Y(_02893_));
 sky130_fd_sc_hd__and2b_1 _09766_ (.A_N(_02893_),
    .B(_02891_),
    .X(_02894_));
 sky130_fd_sc_hd__and2b_1 _09767_ (.A_N(_02891_),
    .B(_02893_),
    .X(_02895_));
 sky130_fd_sc_hd__or2_1 _09768_ (.A(_02894_),
    .B(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__nand2_1 _09769_ (.A(_02889_),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__xnor2_2 _09770_ (.A(_02889_),
    .B(_02896_),
    .Y(_02898_));
 sky130_fd_sc_hd__xnor2_2 _09771_ (.A(_02877_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__or2_1 _09772_ (.A(net147),
    .B(net40),
    .X(_02900_));
 sky130_fd_sc_hd__a21oi_2 _09773_ (.A1(net203),
    .A2(_02750_),
    .B1(_02749_),
    .Y(_02901_));
 sky130_fd_sc_hd__o22a_1 _09774_ (.A1(net141),
    .A2(net16),
    .B1(net7),
    .B2(net139),
    .X(_02902_));
 sky130_fd_sc_hd__xnor2_2 _09775_ (.A(net44),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__and2b_1 _09776_ (.A_N(_02901_),
    .B(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__xnor2_2 _09777_ (.A(_02901_),
    .B(_02903_),
    .Y(_02905_));
 sky130_fd_sc_hd__xnor2_2 _09778_ (.A(_02900_),
    .B(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__nand2_1 _09779_ (.A(_02899_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__xnor2_2 _09780_ (.A(_02899_),
    .B(_02906_),
    .Y(_02908_));
 sky130_fd_sc_hd__xnor2_1 _09781_ (.A(_02866_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__o21ai_2 _09782_ (.A1(_02699_),
    .A2(_02701_),
    .B1(_02697_),
    .Y(_02910_));
 sky130_fd_sc_hd__o22a_1 _09783_ (.A1(net80),
    .A2(net93),
    .B1(net91),
    .B2(net34),
    .X(_02911_));
 sky130_fd_sc_hd__xnor2_1 _09784_ (.A(net114),
    .B(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__o22a_1 _09785_ (.A1(net100),
    .A2(net46),
    .B1(net12),
    .B2(_00311_),
    .X(_02913_));
 sky130_fd_sc_hd__xnor2_1 _09786_ (.A(net111),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__and2_1 _09787_ (.A(_02912_),
    .B(_02914_),
    .X(_02915_));
 sky130_fd_sc_hd__nor2_1 _09788_ (.A(_02912_),
    .B(_02914_),
    .Y(_02916_));
 sky130_fd_sc_hd__nor2_2 _09789_ (.A(_02915_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a31o_1 _09790_ (.A1(_06491_),
    .A2(net44),
    .A3(_02734_),
    .B1(_02733_),
    .X(_02918_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__xor2_2 _09792_ (.A(_02917_),
    .B(_02918_),
    .X(_02920_));
 sky130_fd_sc_hd__xnor2_1 _09793_ (.A(_02910_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__nor2_1 _09794_ (.A(_02909_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_1 _09795_ (.A(_02909_),
    .B(_02921_),
    .Y(_02923_));
 sky130_fd_sc_hd__and2b_1 _09796_ (.A_N(_02922_),
    .B(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__xor2_4 _09797_ (.A(_02861_),
    .B(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__a21bo_2 _09798_ (.A1(_02706_),
    .A2(_02770_),
    .B1_N(_02768_),
    .X(_02926_));
 sky130_fd_sc_hd__a21o_2 _09799_ (.A1(_02692_),
    .A2(_02705_),
    .B1(_02703_),
    .X(_02927_));
 sky130_fd_sc_hd__a21boi_4 _09800_ (.A1(_02707_),
    .A2(_02721_),
    .B1_N(_02720_),
    .Y(_02928_));
 sky130_fd_sc_hd__o21a_2 _09801_ (.A1(_02728_),
    .A2(_02766_),
    .B1(_02765_),
    .X(_02929_));
 sky130_fd_sc_hd__nor2_1 _09802_ (.A(_02928_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__xor2_4 _09803_ (.A(_02928_),
    .B(_02929_),
    .X(_02931_));
 sky130_fd_sc_hd__xnor2_4 _09804_ (.A(_02927_),
    .B(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__a21boi_4 _09805_ (.A1(_02774_),
    .A2(_02778_),
    .B1_N(_02777_),
    .Y(_02933_));
 sky130_fd_sc_hd__xnor2_2 _09806_ (.A(_02932_),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2b_1 _09807_ (.A_N(_02934_),
    .B(_02926_),
    .Y(_02935_));
 sky130_fd_sc_hd__xnor2_4 _09808_ (.A(_02926_),
    .B(_02934_),
    .Y(_02936_));
 sky130_fd_sc_hd__and2_1 _09809_ (.A(_02925_),
    .B(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__xor2_4 _09810_ (.A(_02925_),
    .B(_02936_),
    .X(_02938_));
 sky130_fd_sc_hd__xnor2_4 _09811_ (.A(_02846_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__or2_1 _09812_ (.A(_02845_),
    .B(_02939_),
    .X(_02940_));
 sky130_fd_sc_hd__and2_1 _09813_ (.A(_02845_),
    .B(_02939_),
    .X(_02941_));
 sky130_fd_sc_hd__xnor2_4 _09814_ (.A(_02845_),
    .B(_02939_),
    .Y(_02942_));
 sky130_fd_sc_hd__a21o_1 _09815_ (.A1(_02634_),
    .A2(_02786_),
    .B1(_02787_),
    .X(_02943_));
 sky130_fd_sc_hd__or2_1 _09816_ (.A(_02636_),
    .B(_02788_),
    .X(_02944_));
 sky130_fd_sc_hd__o21a_2 _09817_ (.A1(_02640_),
    .A2(_02944_),
    .B1(_02943_),
    .X(_02945_));
 sky130_fd_sc_hd__xnor2_4 _09818_ (.A(_02942_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__a21oi_1 _09819_ (.A1(_02844_),
    .A2(_02946_),
    .B1(_02242_),
    .Y(_02947_));
 sky130_fd_sc_hd__o21a_1 _09820_ (.A1(_02844_),
    .A2(_02946_),
    .B1(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__and2_1 _09821_ (.A(net151),
    .B(_02170_),
    .X(_02949_));
 sky130_fd_sc_hd__a21oi_1 _09822_ (.A1(_02171_),
    .A2(_02949_),
    .B1(_02318_),
    .Y(_02950_));
 sky130_fd_sc_hd__o21a_1 _09823_ (.A1(_02171_),
    .A2(_02949_),
    .B1(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__o31a_1 _09824_ (.A1(_06316_),
    .A2(_06323_),
    .A3(_02822_),
    .B1(_06317_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(_06340_),
    .A1(_02952_),
    .S(net298),
    .X(_02953_));
 sky130_fd_sc_hd__a21oi_1 _09826_ (.A1(_06312_),
    .A2(_02953_),
    .B1(net241),
    .Y(_02954_));
 sky130_fd_sc_hd__o21a_1 _09827_ (.A1(_06312_),
    .A2(_02953_),
    .B1(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__o21ai_1 _09828_ (.A1(net222),
    .A2(_02806_),
    .B1(_02345_),
    .Y(_02956_));
 sky130_fd_sc_hd__a21boi_1 _09829_ (.A1(net225),
    .A2(_02956_),
    .B1_N(_02338_),
    .Y(_02957_));
 sky130_fd_sc_hd__mux2_1 _09830_ (.A0(_02261_),
    .A1(_02269_),
    .S(net220),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(_02276_),
    .A1(_02300_),
    .S(net220),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _09832_ (.A0(_02958_),
    .A1(_02959_),
    .S(net222),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(_02285_),
    .A1(_02307_),
    .S(_06321_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _09834_ (.A0(_02819_),
    .A1(_02961_),
    .S(net224),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(_02960_),
    .A1(_02962_),
    .S(net226),
    .X(_02963_));
 sky130_fd_sc_hd__a21o_1 _09836_ (.A1(net229),
    .A2(net210),
    .B1(_02315_),
    .X(_02964_));
 sky130_fd_sc_hd__inv_2 _09837_ (.A(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__or4_2 _09838_ (.A(\div_res[3] ),
    .B(\div_res[2] ),
    .C(\div_res[1] ),
    .D(\div_res[0] ),
    .X(_02966_));
 sky130_fd_sc_hd__a21oi_1 _09839_ (.A1(net152),
    .A2(_02966_),
    .B1(\div_res[4] ),
    .Y(_02967_));
 sky130_fd_sc_hd__a311o_1 _09840_ (.A1(\div_res[4] ),
    .A2(net153),
    .A3(_02966_),
    .B1(_02967_),
    .C1(net198),
    .X(_02968_));
 sky130_fd_sc_hd__or2_1 _09841_ (.A(\div_shifter[35] ),
    .B(_02830_),
    .X(_02969_));
 sky130_fd_sc_hd__and3_1 _09842_ (.A(\div_shifter[36] ),
    .B(net234),
    .C(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__a21oi_1 _09843_ (.A1(net234),
    .A2(_02969_),
    .B1(\div_shifter[36] ),
    .Y(_02971_));
 sky130_fd_sc_hd__o32a_1 _09844_ (.A1(net238),
    .A2(_02970_),
    .A3(_02971_),
    .B1(net236),
    .B2(reg1_val[4]),
    .X(_02972_));
 sky130_fd_sc_hd__o221a_1 _09845_ (.A1(net225),
    .A2(net252),
    .B1(net200),
    .B2(_06311_),
    .C1(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__o21a_1 _09846_ (.A1(_02812_),
    .A2(_02813_),
    .B1(_02814_),
    .X(_02974_));
 sky130_fd_sc_hd__nor2_1 _09847_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _09848_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2b_1 _09849_ (.A_N(_02975_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__xnor2_1 _09850_ (.A(_02974_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(_06299_),
    .B(net210),
    .Y(_02979_));
 sky130_fd_sc_hd__o221a_1 _09852_ (.A1(_06310_),
    .A2(_02323_),
    .B1(_02978_),
    .B2(_02979_),
    .C1(_02973_),
    .X(_02980_));
 sky130_fd_sc_hd__o211ai_1 _09853_ (.A1(_06312_),
    .A2(_02327_),
    .B1(_02968_),
    .C1(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__a221o_1 _09854_ (.A1(net245),
    .A2(_02957_),
    .B1(_02963_),
    .B2(_02964_),
    .C1(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__o41a_1 _09855_ (.A1(_02948_),
    .A2(_02951_),
    .A3(_02955_),
    .A4(_02982_),
    .B1(net255),
    .X(_02983_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(curr_PC[4]),
    .B(_02841_),
    .Y(_02984_));
 sky130_fd_sc_hd__or2_1 _09857_ (.A(curr_PC[4]),
    .B(_02841_),
    .X(_02985_));
 sky130_fd_sc_hd__a31o_4 _09858_ (.A1(net258),
    .A2(_02984_),
    .A3(_02985_),
    .B1(_02983_),
    .X(dest_val[4]));
 sky130_fd_sc_hd__a31o_1 _09859_ (.A1(_02688_),
    .A2(_02793_),
    .A3(_02946_),
    .B1(net148),
    .X(_02986_));
 sky130_fd_sc_hd__a21oi_4 _09860_ (.A1(_02846_),
    .A2(_02938_),
    .B1(_02937_),
    .Y(_02987_));
 sky130_fd_sc_hd__o21ai_4 _09861_ (.A1(_02932_),
    .A2(_02933_),
    .B1(_02935_),
    .Y(_02988_));
 sky130_fd_sc_hd__o31ai_4 _09862_ (.A1(_02875_),
    .A2(_02876_),
    .A3(_02898_),
    .B1(_02897_),
    .Y(_02989_));
 sky130_fd_sc_hd__a21oi_4 _09863_ (.A1(_02862_),
    .A2(_02864_),
    .B1(_02863_),
    .Y(_02990_));
 sky130_fd_sc_hd__o22a_1 _09864_ (.A1(net38),
    .A2(net81),
    .B1(net124),
    .B2(net36),
    .X(_02991_));
 sky130_fd_sc_hd__xnor2_1 _09865_ (.A(net121),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__o22a_1 _09866_ (.A1(net80),
    .A2(net57),
    .B1(net94),
    .B2(net34),
    .X(_02993_));
 sky130_fd_sc_hd__xnor2_1 _09867_ (.A(net114),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__and2_1 _09868_ (.A(_02992_),
    .B(_02994_),
    .X(_02995_));
 sky130_fd_sc_hd__nor2_1 _09869_ (.A(_02992_),
    .B(_02994_),
    .Y(_02996_));
 sky130_fd_sc_hd__nor2_2 _09870_ (.A(_02995_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__o22a_1 _09871_ (.A1(net31),
    .A2(_00329_),
    .B1(net83),
    .B2(net30),
    .X(_02998_));
 sky130_fd_sc_hd__xor2_4 _09872_ (.A(net118),
    .B(_02998_),
    .X(_02999_));
 sky130_fd_sc_hd__xnor2_4 _09873_ (.A(_02997_),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2b_1 _09874_ (.A_N(_02990_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__xnor2_4 _09875_ (.A(_02990_),
    .B(_03000_),
    .Y(_03002_));
 sky130_fd_sc_hd__xnor2_4 _09876_ (.A(_02989_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__o21ba_1 _09877_ (.A1(_02885_),
    .A2(_02888_),
    .B1_N(_02884_),
    .X(_03004_));
 sky130_fd_sc_hd__nor2_1 _09878_ (.A(_02894_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_1 _09879_ (.A(_02894_),
    .B(_03004_),
    .Y(_03006_));
 sky130_fd_sc_hd__o21ba_1 _09880_ (.A1(_02873_),
    .A2(_02875_),
    .B1_N(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__or3b_1 _09881_ (.A(_02873_),
    .B(_02875_),
    .C_N(_03006_),
    .X(_03008_));
 sky130_fd_sc_hd__and2b_1 _09882_ (.A_N(_03007_),
    .B(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__o22a_1 _09883_ (.A1(net145),
    .A2(net26),
    .B1(net122),
    .B2(_00230_),
    .X(_03010_));
 sky130_fd_sc_hd__xnor2_1 _09884_ (.A(net68),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__or2_1 _09885_ (.A(net139),
    .B(net40),
    .X(_03012_));
 sky130_fd_sc_hd__nor2_1 _09886_ (.A(_03011_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__xor2_1 _09887_ (.A(_03011_),
    .B(_03012_),
    .X(_03014_));
 sky130_fd_sc_hd__o22a_1 _09888_ (.A1(net143),
    .A2(net16),
    .B1(net7),
    .B2(net141),
    .X(_03015_));
 sky130_fd_sc_hd__xnor2_1 _09889_ (.A(net43),
    .B(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__and2_1 _09890_ (.A(_03014_),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__nor2_1 _09891_ (.A(_03014_),
    .B(_03016_),
    .Y(_03018_));
 sky130_fd_sc_hd__or2_1 _09892_ (.A(_03017_),
    .B(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__o22a_1 _09893_ (.A1(net136),
    .A2(net18),
    .B1(net9),
    .B2(net170),
    .X(_03020_));
 sky130_fd_sc_hd__xnor2_1 _09894_ (.A(net183),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__o22a_1 _09895_ (.A1(net133),
    .A2(net24),
    .B1(net20),
    .B2(net135),
    .X(_03022_));
 sky130_fd_sc_hd__xnor2_2 _09896_ (.A(net186),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__inv_2 _09897_ (.A(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__xnor2_1 _09898_ (.A(net206),
    .B(_03023_),
    .Y(_03025_));
 sky130_fd_sc_hd__nand2b_1 _09899_ (.A_N(_03021_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__xnor2_1 _09900_ (.A(_03021_),
    .B(_03025_),
    .Y(_03027_));
 sky130_fd_sc_hd__o22a_1 _09901_ (.A1(net58),
    .A2(net98),
    .B1(net56),
    .B2(net65),
    .X(_03028_));
 sky130_fd_sc_hd__xor2_1 _09902_ (.A(net129),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__a21o_1 _09903_ (.A1(_00267_),
    .A2(_00269_),
    .B1(net107),
    .X(_03030_));
 sky130_fd_sc_hd__or2_1 _09904_ (.A(net103),
    .B(net61),
    .X(_03031_));
 sky130_fd_sc_hd__a21o_1 _09905_ (.A1(_03030_),
    .A2(_03031_),
    .B1(net173),
    .X(_03032_));
 sky130_fd_sc_hd__nand3_1 _09906_ (.A(net173),
    .B(_03030_),
    .C(_03031_),
    .Y(_03033_));
 sky130_fd_sc_hd__o22a_1 _09907_ (.A1(net62),
    .A2(net95),
    .B1(net54),
    .B2(net77),
    .X(_03034_));
 sky130_fd_sc_hd__xnor2_1 _09908_ (.A(_00319_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__nand3_1 _09909_ (.A(_03032_),
    .B(_03033_),
    .C(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__a21o_1 _09910_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_03035_),
    .X(_03037_));
 sky130_fd_sc_hd__nand3_1 _09911_ (.A(_03029_),
    .B(_03036_),
    .C(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__a21o_1 _09912_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_03029_),
    .X(_03039_));
 sky130_fd_sc_hd__and3_1 _09913_ (.A(_02915_),
    .B(_03038_),
    .C(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__a21oi_1 _09914_ (.A1(_03038_),
    .A2(_03039_),
    .B1(_02915_),
    .Y(_03041_));
 sky130_fd_sc_hd__nor3b_2 _09915_ (.A(_03040_),
    .B(_03041_),
    .C_N(_03027_),
    .Y(_03042_));
 sky130_fd_sc_hd__o21ba_1 _09916_ (.A1(_03040_),
    .A2(_03041_),
    .B1_N(_03027_),
    .X(_03043_));
 sky130_fd_sc_hd__or3_1 _09917_ (.A(_03019_),
    .B(_03042_),
    .C(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__o21ai_2 _09918_ (.A1(_03042_),
    .A2(_03043_),
    .B1(_03019_),
    .Y(_03045_));
 sky130_fd_sc_hd__and3_1 _09919_ (.A(_03009_),
    .B(_03044_),
    .C(_03045_),
    .X(_03046_));
 sky130_fd_sc_hd__a21oi_1 _09920_ (.A1(_03044_),
    .A2(_03045_),
    .B1(_03009_),
    .Y(_03047_));
 sky130_fd_sc_hd__nor2_1 _09921_ (.A(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__o21ai_2 _09922_ (.A1(_02854_),
    .A2(_02856_),
    .B1(_02852_),
    .Y(_03049_));
 sky130_fd_sc_hd__o22a_1 _09923_ (.A1(net75),
    .A2(net53),
    .B1(net51),
    .B2(net72),
    .X(_03050_));
 sky130_fd_sc_hd__xnor2_1 _09924_ (.A(net89),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__o32a_1 _09925_ (.A1(net101),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net46),
    .B2(net105),
    .X(_03052_));
 sky130_fd_sc_hd__xnor2_1 _09926_ (.A(_06504_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__and2_1 _09927_ (.A(_03051_),
    .B(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__nor2_1 _09928_ (.A(_03051_),
    .B(_03053_),
    .Y(_03055_));
 sky130_fd_sc_hd__nor2_1 _09929_ (.A(_03054_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__o22a_1 _09930_ (.A1(net69),
    .A2(net48),
    .B1(net13),
    .B2(net109),
    .X(_03057_));
 sky130_fd_sc_hd__xnor2_2 _09931_ (.A(net85),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__xor2_2 _09932_ (.A(_03056_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__a41o_1 _09933_ (.A1(_06477_),
    .A2(_06478_),
    .A3(net43),
    .A4(_02905_),
    .B1(_02904_),
    .X(_03060_));
 sky130_fd_sc_hd__nand2_1 _09934_ (.A(_03059_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__xor2_2 _09935_ (.A(_03059_),
    .B(_03060_),
    .X(_03062_));
 sky130_fd_sc_hd__xor2_1 _09936_ (.A(_03049_),
    .B(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__nand2_1 _09937_ (.A(_03048_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__or2_1 _09938_ (.A(_03048_),
    .B(_03063_),
    .X(_03065_));
 sky130_fd_sc_hd__nand2_2 _09939_ (.A(_03064_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__xor2_4 _09940_ (.A(_03003_),
    .B(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__a21o_2 _09941_ (.A1(_02861_),
    .A2(_02923_),
    .B1(_02922_),
    .X(_03068_));
 sky130_fd_sc_hd__o21ai_4 _09942_ (.A1(_02857_),
    .A2(_02858_),
    .B1(_02860_),
    .Y(_03069_));
 sky130_fd_sc_hd__o21a_1 _09943_ (.A1(_02866_),
    .A2(_02908_),
    .B1(_02907_),
    .X(_03070_));
 sky130_fd_sc_hd__o21ai_2 _09944_ (.A1(_02866_),
    .A2(_02908_),
    .B1(_02907_),
    .Y(_03071_));
 sky130_fd_sc_hd__a21boi_4 _09945_ (.A1(_02910_),
    .A2(_02920_),
    .B1_N(_02919_),
    .Y(_03072_));
 sky130_fd_sc_hd__nor2_1 _09946_ (.A(_03070_),
    .B(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__xnor2_4 _09947_ (.A(_03071_),
    .B(_03072_),
    .Y(_03074_));
 sky130_fd_sc_hd__xnor2_4 _09948_ (.A(_03069_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__a21oi_4 _09949_ (.A1(_02927_),
    .A2(_02931_),
    .B1(_02930_),
    .Y(_03076_));
 sky130_fd_sc_hd__xnor2_2 _09950_ (.A(_03075_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand2b_1 _09951_ (.A_N(_03077_),
    .B(_03068_),
    .Y(_03078_));
 sky130_fd_sc_hd__xnor2_4 _09952_ (.A(_03068_),
    .B(_03077_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_1 _09953_ (.A(_03067_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__xor2_4 _09954_ (.A(_03067_),
    .B(_03079_),
    .X(_03081_));
 sky130_fd_sc_hd__xnor2_4 _09955_ (.A(_02988_),
    .B(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__or2_1 _09956_ (.A(_02987_),
    .B(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__and2_1 _09957_ (.A(_02987_),
    .B(_03082_),
    .X(_03084_));
 sky130_fd_sc_hd__xnor2_4 _09958_ (.A(_02987_),
    .B(_03082_),
    .Y(_03085_));
 sky130_fd_sc_hd__a21oi_1 _09959_ (.A1(_02786_),
    .A2(_02940_),
    .B1(_02941_),
    .Y(_03086_));
 sky130_fd_sc_hd__or2_1 _09960_ (.A(_02788_),
    .B(_02942_),
    .X(_03087_));
 sky130_fd_sc_hd__o21ba_1 _09961_ (.A1(_02792_),
    .A2(_03087_),
    .B1_N(_03086_),
    .X(_03088_));
 sky130_fd_sc_hd__xnor2_2 _09962_ (.A(_03085_),
    .B(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__a21oi_1 _09963_ (.A1(_02986_),
    .A2(_03089_),
    .B1(_02242_),
    .Y(_03090_));
 sky130_fd_sc_hd__o21a_1 _09964_ (.A1(_02986_),
    .A2(_03089_),
    .B1(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__o21ai_1 _09965_ (.A1(net148),
    .A2(_02172_),
    .B1(_02173_),
    .Y(_03092_));
 sky130_fd_sc_hd__or3_1 _09966_ (.A(net148),
    .B(_02172_),
    .C(_02173_),
    .X(_03093_));
 sky130_fd_sc_hd__o21a_1 _09967_ (.A1(_06310_),
    .A2(_02952_),
    .B1(_06311_),
    .X(_03094_));
 sky130_fd_sc_hd__nor2_1 _09968_ (.A(net303),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a21oi_1 _09969_ (.A1(net303),
    .A2(_06342_),
    .B1(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__xnor2_1 _09970_ (.A(_06306_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__o21ai_1 _09971_ (.A1(net222),
    .A2(_02658_),
    .B1(_02345_),
    .Y(_03098_));
 sky130_fd_sc_hd__a21boi_2 _09972_ (.A1(net225),
    .A2(_03098_),
    .B1_N(_02338_),
    .Y(_03099_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(_02477_),
    .A1(_02481_),
    .S(net220),
    .X(_03100_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(_02484_),
    .A1(_02495_),
    .S(net221),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _09975_ (.A0(_03100_),
    .A1(_03101_),
    .S(net222),
    .X(_03102_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(_02489_),
    .A1(_02498_),
    .S(_06321_),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _09977_ (.A0(_02647_),
    .A1(_03103_),
    .S(net224),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(_03102_),
    .A1(_03104_),
    .S(net226),
    .X(_03105_));
 sky130_fd_sc_hd__o21a_1 _09979_ (.A1(\div_res[4] ),
    .A2(_02966_),
    .B1(net152),
    .X(_03106_));
 sky130_fd_sc_hd__nand2_1 _09980_ (.A(\div_res[5] ),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__o21a_1 _09981_ (.A1(\div_res[5] ),
    .A2(_03106_),
    .B1(_02330_),
    .X(_03108_));
 sky130_fd_sc_hd__or2_1 _09982_ (.A(\div_shifter[36] ),
    .B(_02969_),
    .X(_03109_));
 sky130_fd_sc_hd__a21oi_1 _09983_ (.A1(net234),
    .A2(_03109_),
    .B1(\div_shifter[37] ),
    .Y(_03110_));
 sky130_fd_sc_hd__a31o_1 _09984_ (.A1(\div_shifter[37] ),
    .A2(net235),
    .A3(_03109_),
    .B1(net238),
    .X(_03111_));
 sky130_fd_sc_hd__o22a_1 _09985_ (.A1(reg1_val[5]),
    .A2(net236),
    .B1(_03110_),
    .B2(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__o221ai_1 _09986_ (.A1(_06301_),
    .A2(net252),
    .B1(net200),
    .B2(_06305_),
    .C1(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__a221o_1 _09987_ (.A1(_06304_),
    .A2(net273),
    .B1(net240),
    .B2(_06306_),
    .C1(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__o21a_1 _09988_ (.A1(_02974_),
    .A2(_02975_),
    .B1(_02976_),
    .X(_03115_));
 sky130_fd_sc_hd__nor2_1 _09989_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2_1 _09990_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03117_));
 sky130_fd_sc_hd__and2b_1 _09991_ (.A_N(_03116_),
    .B(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__xnor2_1 _09992_ (.A(_03115_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__a31o_1 _09993_ (.A1(net260),
    .A2(net210),
    .A3(_03119_),
    .B1(_03114_),
    .X(_03120_));
 sky130_fd_sc_hd__a221o_1 _09994_ (.A1(_02964_),
    .A2(_03105_),
    .B1(_03107_),
    .B2(_03108_),
    .C1(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__a221o_1 _09995_ (.A1(_02324_),
    .A2(_03097_),
    .B1(_03099_),
    .B2(net246),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__a311o_1 _09996_ (.A1(_02317_),
    .A2(_03092_),
    .A3(_03093_),
    .B1(_03122_),
    .C1(_03091_),
    .X(_03123_));
 sky130_fd_sc_hd__a31o_1 _09997_ (.A1(curr_PC[3]),
    .A2(curr_PC[4]),
    .A3(_02530_),
    .B1(curr_PC[5]),
    .X(_03124_));
 sky130_fd_sc_hd__and3_1 _09998_ (.A(curr_PC[4]),
    .B(curr_PC[5]),
    .C(_02841_),
    .X(_03125_));
 sky130_fd_sc_hd__nor2_1 _09999_ (.A(net253),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__a22o_4 _10000_ (.A1(net253),
    .A2(_03123_),
    .B1(_03124_),
    .B2(_03126_),
    .X(dest_val[5]));
 sky130_fd_sc_hd__nand2_1 _10001_ (.A(_02946_),
    .B(_03089_),
    .Y(_03127_));
 sky130_fd_sc_hd__and3_1 _10002_ (.A(_02843_),
    .B(_02946_),
    .C(_03089_),
    .X(_03128_));
 sky130_fd_sc_hd__or2_1 _10003_ (.A(net148),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__a21boi_4 _10004_ (.A1(_02988_),
    .A2(_03081_),
    .B1_N(_03080_),
    .Y(_03130_));
 sky130_fd_sc_hd__o21ai_4 _10005_ (.A1(_03075_),
    .A2(_03076_),
    .B1(_03078_),
    .Y(_03131_));
 sky130_fd_sc_hd__nor2_2 _10006_ (.A(_03040_),
    .B(_03042_),
    .Y(_03132_));
 sky130_fd_sc_hd__o22a_1 _10007_ (.A1(net31),
    .A2(net93),
    .B1(net91),
    .B2(net30),
    .X(_03133_));
 sky130_fd_sc_hd__xnor2_1 _10008_ (.A(net118),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__o22a_1 _10009_ (.A1(net109),
    .A2(net46),
    .B1(net12),
    .B2(net105),
    .X(_03135_));
 sky130_fd_sc_hd__xnor2_1 _10010_ (.A(net111),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__and2_1 _10011_ (.A(_03134_),
    .B(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(_03134_),
    .B(_03136_),
    .Y(_03138_));
 sky130_fd_sc_hd__nor2_1 _10013_ (.A(_03137_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__a2bb2o_1 _10014_ (.A1_N(net34),
    .A2_N(net57),
    .B1(net99),
    .B2(_06508_),
    .X(_03140_));
 sky130_fd_sc_hd__xnor2_1 _10015_ (.A(net115),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__xnor2_1 _10016_ (.A(_03139_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__o21ai_1 _10017_ (.A1(_03005_),
    .A2(_03007_),
    .B1(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__or3_1 _10018_ (.A(_03005_),
    .B(_03007_),
    .C(_03142_),
    .X(_03144_));
 sky130_fd_sc_hd__nand2_2 _10019_ (.A(_03143_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__xor2_4 _10020_ (.A(_03132_),
    .B(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__o21bai_1 _10021_ (.A1(_02996_),
    .A2(_02999_),
    .B1_N(_02995_),
    .Y(_03147_));
 sky130_fd_sc_hd__o22a_1 _10022_ (.A1(net77),
    .A2(net52),
    .B1(net50),
    .B2(net75),
    .X(_03148_));
 sky130_fd_sc_hd__xnor2_1 _10023_ (.A(net89),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__o22a_1 _10024_ (.A1(net72),
    .A2(net49),
    .B1(net14),
    .B2(net69),
    .X(_03150_));
 sky130_fd_sc_hd__xnor2_1 _10025_ (.A(net85),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_1 _10026_ (.A(_03149_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__or2_1 _10027_ (.A(_03149_),
    .B(_03151_),
    .X(_03153_));
 sky130_fd_sc_hd__and2_1 _10028_ (.A(_03152_),
    .B(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__o21ai_1 _10029_ (.A1(_03013_),
    .A2(_03017_),
    .B1(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__or3_1 _10030_ (.A(_03013_),
    .B(_03017_),
    .C(_03154_),
    .X(_03156_));
 sky130_fd_sc_hd__and2_1 _10031_ (.A(_03155_),
    .B(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__nand2_1 _10032_ (.A(_03147_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__xnor2_1 _10033_ (.A(_03147_),
    .B(_03157_),
    .Y(_03159_));
 sky130_fd_sc_hd__a21bo_1 _10034_ (.A1(net206),
    .A2(_03024_),
    .B1_N(_03026_),
    .X(_03160_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_06522_),
    .B(net45),
    .Y(_03161_));
 sky130_fd_sc_hd__a21oi_1 _10036_ (.A1(_03036_),
    .A2(_03038_),
    .B1(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__and3_1 _10037_ (.A(_03036_),
    .B(_03038_),
    .C(_03161_),
    .X(_03163_));
 sky130_fd_sc_hd__nor2_1 _10038_ (.A(_03162_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__and2_1 _10039_ (.A(_03160_),
    .B(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__xor2_2 _10040_ (.A(_03160_),
    .B(_03164_),
    .X(_03166_));
 sky130_fd_sc_hd__a21o_1 _10041_ (.A1(_03056_),
    .A2(_03058_),
    .B1(_03054_),
    .X(_03167_));
 sky130_fd_sc_hd__o22a_1 _10042_ (.A1(net61),
    .A2(net98),
    .B1(net56),
    .B2(net58),
    .X(_03168_));
 sky130_fd_sc_hd__xnor2_1 _10043_ (.A(net129),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__o22a_1 _10044_ (.A1(net107),
    .A2(net24),
    .B1(net22),
    .B2(net103),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_1 _10045_ (.A(net173),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__o22a_1 _10046_ (.A1(net65),
    .A2(net95),
    .B1(net54),
    .B2(net62),
    .X(_03172_));
 sky130_fd_sc_hd__xnor2_1 _10047_ (.A(net126),
    .B(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__or2_1 _10048_ (.A(_03171_),
    .B(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__xnor2_1 _10049_ (.A(_03171_),
    .B(_03173_),
    .Y(_03175_));
 sky130_fd_sc_hd__xnor2_1 _10050_ (.A(_03169_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand2b_1 _10051_ (.A_N(_03176_),
    .B(_03167_),
    .Y(_03177_));
 sky130_fd_sc_hd__xnor2_1 _10052_ (.A(_03167_),
    .B(_03176_),
    .Y(_03178_));
 sky130_fd_sc_hd__o22a_1 _10053_ (.A1(net133),
    .A2(net20),
    .B1(net18),
    .B2(net135),
    .X(_03179_));
 sky130_fd_sc_hd__xnor2_2 _10054_ (.A(net186),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__inv_2 _10055_ (.A(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__a21oi_1 _10056_ (.A1(_00176_),
    .A2(net10),
    .B1(net183),
    .Y(_03182_));
 sky130_fd_sc_hd__a31o_2 _10057_ (.A1(net183),
    .A2(_00178_),
    .A3(net10),
    .B1(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__xor2_2 _10058_ (.A(_03180_),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__nand2_1 _10059_ (.A(_03178_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__or2_1 _10060_ (.A(_03178_),
    .B(_03184_),
    .X(_03186_));
 sky130_fd_sc_hd__xnor2_1 _10061_ (.A(_03178_),
    .B(_03184_),
    .Y(_03187_));
 sky130_fd_sc_hd__o22a_2 _10062_ (.A1(_00230_),
    .A2(net124),
    .B1(net122),
    .B2(net26),
    .X(_03188_));
 sky130_fd_sc_hd__xnor2_4 _10063_ (.A(net68),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__o22a_2 _10064_ (.A1(net145),
    .A2(net16),
    .B1(net7),
    .B2(net143),
    .X(_03190_));
 sky130_fd_sc_hd__xnor2_4 _10065_ (.A(net43),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__o22a_2 _10066_ (.A1(net38),
    .A2(net83),
    .B1(net81),
    .B2(net36),
    .X(_03192_));
 sky130_fd_sc_hd__xnor2_4 _10067_ (.A(net121),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _10068_ (.A(_03191_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__xor2_4 _10069_ (.A(_03191_),
    .B(_03193_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2b_1 _10070_ (.A_N(_03189_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__xnor2_4 _10071_ (.A(_03189_),
    .B(_03195_),
    .Y(_03197_));
 sky130_fd_sc_hd__xnor2_2 _10072_ (.A(_03187_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__xnor2_1 _10073_ (.A(_03166_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__nor2_1 _10074_ (.A(_03159_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _10075_ (.A(_03159_),
    .B(_03199_),
    .Y(_03201_));
 sky130_fd_sc_hd__and2b_1 _10076_ (.A_N(_03200_),
    .B(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__xor2_4 _10077_ (.A(_03146_),
    .B(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__o21ai_2 _10078_ (.A1(_03003_),
    .A2(_03066_),
    .B1(_03064_),
    .Y(_03204_));
 sky130_fd_sc_hd__a21o_1 _10079_ (.A1(_03069_),
    .A2(_03074_),
    .B1(_03073_),
    .X(_03205_));
 sky130_fd_sc_hd__a21bo_1 _10080_ (.A1(_02989_),
    .A2(_03002_),
    .B1_N(_03001_),
    .X(_03206_));
 sky130_fd_sc_hd__a21boi_2 _10081_ (.A1(_03009_),
    .A2(_03045_),
    .B1_N(_03044_),
    .Y(_03207_));
 sky130_fd_sc_hd__a21boi_2 _10082_ (.A1(_03049_),
    .A2(_03062_),
    .B1_N(_03061_),
    .Y(_03208_));
 sky130_fd_sc_hd__nor2_1 _10083_ (.A(_03207_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__xor2_2 _10084_ (.A(_03207_),
    .B(_03208_),
    .X(_03210_));
 sky130_fd_sc_hd__xor2_2 _10085_ (.A(_03206_),
    .B(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__xnor2_2 _10086_ (.A(_03205_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2b_1 _10087_ (.A_N(_03212_),
    .B(_03204_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_2 _10088_ (.A(_03204_),
    .B(_03212_),
    .Y(_03214_));
 sky130_fd_sc_hd__and2_1 _10089_ (.A(_03203_),
    .B(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__xor2_4 _10090_ (.A(_03203_),
    .B(_03214_),
    .X(_03216_));
 sky130_fd_sc_hd__xnor2_4 _10091_ (.A(_03131_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__or2_1 _10092_ (.A(_03130_),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__and2_1 _10093_ (.A(_03130_),
    .B(_03217_),
    .X(_03219_));
 sky130_fd_sc_hd__xnor2_4 _10094_ (.A(_03130_),
    .B(_03217_),
    .Y(_03220_));
 sky130_fd_sc_hd__nor2_1 _10095_ (.A(_02942_),
    .B(_03085_),
    .Y(_03221_));
 sky130_fd_sc_hd__or2_1 _10096_ (.A(_02942_),
    .B(_03085_),
    .X(_03222_));
 sky130_fd_sc_hd__a21oi_1 _10097_ (.A1(_02940_),
    .A2(_03083_),
    .B1(_03084_),
    .Y(_03223_));
 sky130_fd_sc_hd__o21ba_1 _10098_ (.A1(_02943_),
    .A2(_03222_),
    .B1_N(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__o41a_2 _10099_ (.A1(_02640_),
    .A2(_02942_),
    .A3(_02944_),
    .A4(_03085_),
    .B1(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__xnor2_4 _10100_ (.A(_03220_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__a21oi_1 _10101_ (.A1(_03129_),
    .A2(_03226_),
    .B1(_02242_),
    .Y(_03227_));
 sky130_fd_sc_hd__o21ai_1 _10102_ (.A1(_03129_),
    .A2(_03226_),
    .B1(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__o21a_1 _10103_ (.A1(net148),
    .A2(_02174_),
    .B1(_02175_),
    .X(_03229_));
 sky130_fd_sc_hd__or3_1 _10104_ (.A(net148),
    .B(_02174_),
    .C(_02175_),
    .X(_03230_));
 sky130_fd_sc_hd__or3b_1 _10105_ (.A(_02318_),
    .B(_03229_),
    .C_N(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__o21ai_1 _10106_ (.A1(_06303_),
    .A2(_03094_),
    .B1(_06305_),
    .Y(_03232_));
 sky130_fd_sc_hd__mux2_1 _10107_ (.A0(_06344_),
    .A1(_03232_),
    .S(net298),
    .X(_03233_));
 sky130_fd_sc_hd__nand2_1 _10108_ (.A(_06298_),
    .B(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__o21a_1 _10109_ (.A1(_06298_),
    .A2(_03233_),
    .B1(net242),
    .X(_03235_));
 sky130_fd_sc_hd__o21a_1 _10110_ (.A1(net222),
    .A2(_02492_),
    .B1(_02345_),
    .X(_03236_));
 sky130_fd_sc_hd__o21ai_2 _10111_ (.A1(net226),
    .A2(_03236_),
    .B1(_02338_),
    .Y(_03237_));
 sky130_fd_sc_hd__or2_1 _10112_ (.A(_06321_),
    .B(_02653_),
    .X(_03238_));
 sky130_fd_sc_hd__o211a_1 _10113_ (.A1(net221),
    .A2(_02651_),
    .B1(_03238_),
    .C1(net224),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(_02654_),
    .A1(_02659_),
    .S(net221),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(_02657_),
    .A1(_02660_),
    .S(_06321_),
    .X(_03241_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(_02525_),
    .A1(_03241_),
    .S(net224),
    .X(_03242_));
 sky130_fd_sc_hd__a211o_1 _10117_ (.A1(net223),
    .A2(_03240_),
    .B1(_03239_),
    .C1(net226),
    .X(_03243_));
 sky130_fd_sc_hd__o21ai_1 _10118_ (.A1(net225),
    .A2(_03242_),
    .B1(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__or3_1 _10119_ (.A(\div_res[5] ),
    .B(\div_res[4] ),
    .C(_02966_),
    .X(_03245_));
 sky130_fd_sc_hd__a21oi_1 _10120_ (.A1(net152),
    .A2(_03245_),
    .B1(\div_res[6] ),
    .Y(_03246_));
 sky130_fd_sc_hd__a31o_1 _10121_ (.A1(\div_res[6] ),
    .A2(net152),
    .A3(_03245_),
    .B1(net198),
    .X(_03247_));
 sky130_fd_sc_hd__or3_1 _10122_ (.A(\div_shifter[37] ),
    .B(\div_shifter[36] ),
    .C(_02969_),
    .X(_03248_));
 sky130_fd_sc_hd__a21oi_1 _10123_ (.A1(net235),
    .A2(_03248_),
    .B1(\div_shifter[38] ),
    .Y(_03249_));
 sky130_fd_sc_hd__a31o_1 _10124_ (.A1(\div_shifter[38] ),
    .A2(net235),
    .A3(_03248_),
    .B1(net239),
    .X(_03250_));
 sky130_fd_sc_hd__o22ai_2 _10125_ (.A1(reg1_val[6]),
    .A2(net236),
    .B1(_03249_),
    .B2(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__a221o_1 _10126_ (.A1(_06294_),
    .A2(_06455_),
    .B1(net201),
    .B2(_06296_),
    .C1(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__a221o_1 _10127_ (.A1(_06295_),
    .A2(net273),
    .B1(net240),
    .B2(_06298_),
    .C1(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__o21a_1 _10128_ (.A1(_03115_),
    .A2(_03116_),
    .B1(_03117_),
    .X(_03254_));
 sky130_fd_sc_hd__nor2_1 _10129_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03255_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03256_));
 sky130_fd_sc_hd__and2b_1 _10131_ (.A_N(_03255_),
    .B(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__xnor2_1 _10132_ (.A(_03254_),
    .B(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__a31oi_1 _10133_ (.A1(net261),
    .A2(net210),
    .A3(_03258_),
    .B1(_03253_),
    .Y(_03259_));
 sky130_fd_sc_hd__o221a_1 _10134_ (.A1(_02965_),
    .A2(_03244_),
    .B1(_03246_),
    .B2(_03247_),
    .C1(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__o21ai_2 _10135_ (.A1(_02247_),
    .A2(_03237_),
    .B1(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__a21oi_1 _10136_ (.A1(_03234_),
    .A2(_03235_),
    .B1(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__a31o_2 _10137_ (.A1(_03228_),
    .A2(_03231_),
    .A3(_03262_),
    .B1(net259),
    .X(_03263_));
 sky130_fd_sc_hd__and2_2 _10138_ (.A(curr_PC[6]),
    .B(_03125_),
    .X(_03264_));
 sky130_fd_sc_hd__o21ai_2 _10139_ (.A1(curr_PC[6]),
    .A2(_03125_),
    .B1(net258),
    .Y(_03265_));
 sky130_fd_sc_hd__o21ai_4 _10140_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_03263_),
    .Y(dest_val[6]));
 sky130_fd_sc_hd__a21oi_1 _10141_ (.A1(_03128_),
    .A2(_03226_),
    .B1(net148),
    .Y(_03266_));
 sky130_fd_sc_hd__a21oi_2 _10142_ (.A1(_03131_),
    .A2(_03216_),
    .B1(_03215_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21bo_1 _10143_ (.A1(_03205_),
    .A2(_03211_),
    .B1_N(_03213_),
    .X(_03268_));
 sky130_fd_sc_hd__o22a_1 _10144_ (.A1(net16),
    .A2(net122),
    .B1(net7),
    .B2(net145),
    .X(_03269_));
 sky130_fd_sc_hd__xnor2_1 _10145_ (.A(net43),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__o21ai_1 _10146_ (.A1(_03181_),
    .A2(_03183_),
    .B1(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__or3_1 _10147_ (.A(_03181_),
    .B(_03183_),
    .C(_03270_),
    .X(_03272_));
 sky130_fd_sc_hd__nand2_1 _10148_ (.A(_03271_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_2 _10149_ (.A(_06513_),
    .B(net45),
    .Y(_03274_));
 sky130_fd_sc_hd__xnor2_2 _10150_ (.A(_03273_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__o21a_1 _10151_ (.A1(_03169_),
    .A2(_03175_),
    .B1(_03174_),
    .X(_03276_));
 sky130_fd_sc_hd__o22a_1 _10152_ (.A1(net103),
    .A2(net24),
    .B1(net20),
    .B2(net107),
    .X(_03277_));
 sky130_fd_sc_hd__xnor2_2 _10153_ (.A(net173),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__and2b_1 _10154_ (.A_N(_03278_),
    .B(net183),
    .X(_03279_));
 sky130_fd_sc_hd__xor2_2 _10155_ (.A(net183),
    .B(_03278_),
    .X(_03280_));
 sky130_fd_sc_hd__o22a_1 _10156_ (.A1(net133),
    .A2(net18),
    .B1(net9),
    .B2(net135),
    .X(_03281_));
 sky130_fd_sc_hd__xnor2_2 _10157_ (.A(net186),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__xnor2_2 _10158_ (.A(_03280_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(_03276_),
    .B(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__xor2_2 _10160_ (.A(_03276_),
    .B(_03283_),
    .X(_03285_));
 sky130_fd_sc_hd__xor2_2 _10161_ (.A(_03152_),
    .B(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__o22a_1 _10162_ (.A1(net28),
    .A2(net81),
    .B1(net124),
    .B2(net26),
    .X(_03287_));
 sky130_fd_sc_hd__xnor2_1 _10163_ (.A(net68),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__o22ai_1 _10164_ (.A1(net31),
    .A2(net57),
    .B1(net93),
    .B2(net29),
    .Y(_03289_));
 sky130_fd_sc_hd__xor2_1 _10165_ (.A(net118),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__nand2b_1 _10166_ (.A_N(_03288_),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__xor2_1 _10167_ (.A(_03288_),
    .B(_03290_),
    .X(_03292_));
 sky130_fd_sc_hd__o22a_1 _10168_ (.A1(net38),
    .A2(net91),
    .B1(net83),
    .B2(net36),
    .X(_03293_));
 sky130_fd_sc_hd__xnor2_1 _10169_ (.A(net121),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nand2b_1 _10170_ (.A_N(_03292_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2b_1 _10171_ (.A_N(_03294_),
    .B(_03292_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_1 _10172_ (.A(_03295_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__or2_1 _10173_ (.A(_03286_),
    .B(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__xnor2_2 _10174_ (.A(_03286_),
    .B(_03297_),
    .Y(_03299_));
 sky130_fd_sc_hd__xor2_1 _10175_ (.A(_03275_),
    .B(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__o21ba_1 _10176_ (.A1(_03138_),
    .A2(_03141_),
    .B1_N(_03137_),
    .X(_03301_));
 sky130_fd_sc_hd__o22a_1 _10177_ (.A1(net22),
    .A2(net98),
    .B1(net56),
    .B2(net61),
    .X(_03302_));
 sky130_fd_sc_hd__xor2_1 _10178_ (.A(net129),
    .B(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__o22a_1 _10179_ (.A1(net62),
    .A2(net52),
    .B1(net50),
    .B2(net77),
    .X(_03304_));
 sky130_fd_sc_hd__xnor2_1 _10180_ (.A(net89),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__nand2_1 _10181_ (.A(_03303_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__xnor2_1 _10182_ (.A(_03303_),
    .B(_03305_),
    .Y(_03307_));
 sky130_fd_sc_hd__o22a_1 _10183_ (.A1(net58),
    .A2(net95),
    .B1(net54),
    .B2(net65),
    .X(_03308_));
 sky130_fd_sc_hd__xnor2_1 _10184_ (.A(net128),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__xnor2_1 _10185_ (.A(_03307_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__a21oi_1 _10186_ (.A1(_03194_),
    .A2(_03196_),
    .B1(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__and3_1 _10187_ (.A(_03194_),
    .B(_03196_),
    .C(_03310_),
    .X(_03312_));
 sky130_fd_sc_hd__nor2_1 _10188_ (.A(_03311_),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__and2b_1 _10189_ (.A_N(_03301_),
    .B(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__xnor2_1 _10190_ (.A(_03301_),
    .B(_03313_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _10191_ (.A(_03300_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__or2_1 _10192_ (.A(_03300_),
    .B(_03315_),
    .X(_03317_));
 sky130_fd_sc_hd__nand2_1 _10193_ (.A(_03316_),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2_1 _10194_ (.A(_03177_),
    .B(_03185_),
    .Y(_03319_));
 sky130_fd_sc_hd__o22a_1 _10195_ (.A1(net79),
    .A2(net105),
    .B1(net100),
    .B2(net33),
    .X(_03320_));
 sky130_fd_sc_hd__xnor2_1 _10196_ (.A(net114),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__o22a_1 _10197_ (.A1(net74),
    .A2(net48),
    .B1(net13),
    .B2(net71),
    .X(_03322_));
 sky130_fd_sc_hd__xnor2_1 _10198_ (.A(net85),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__and2_1 _10199_ (.A(_03321_),
    .B(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__nor2_1 _10200_ (.A(_03321_),
    .B(_03323_),
    .Y(_03325_));
 sky130_fd_sc_hd__nor2_1 _10201_ (.A(_03324_),
    .B(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__o22a_1 _10202_ (.A1(net69),
    .A2(net46),
    .B1(net11),
    .B2(net108),
    .X(_03327_));
 sky130_fd_sc_hd__xnor2_1 _10203_ (.A(net110),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__xnor2_1 _10204_ (.A(_03326_),
    .B(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__o21a_1 _10205_ (.A1(_03162_),
    .A2(_03165_),
    .B1(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__nor3_1 _10206_ (.A(_03162_),
    .B(_03165_),
    .C(_03329_),
    .Y(_03331_));
 sky130_fd_sc_hd__nor2_1 _10207_ (.A(_03330_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__xnor2_1 _10208_ (.A(_03319_),
    .B(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__xor2_1 _10209_ (.A(_03318_),
    .B(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__a21o_1 _10210_ (.A1(_03146_),
    .A2(_03201_),
    .B1(_03200_),
    .X(_03335_));
 sky130_fd_sc_hd__o21ai_2 _10211_ (.A1(_03132_),
    .A2(_03145_),
    .B1(_03143_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _10212_ (.A(_03155_),
    .B(_03158_),
    .Y(_03337_));
 sky130_fd_sc_hd__a32oi_4 _10213_ (.A1(_03185_),
    .A2(_03186_),
    .A3(_03197_),
    .B1(_03198_),
    .B2(_03166_),
    .Y(_03338_));
 sky130_fd_sc_hd__a21oi_1 _10214_ (.A1(_03155_),
    .A2(_03158_),
    .B1(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__xnor2_2 _10215_ (.A(_03337_),
    .B(_03338_),
    .Y(_03340_));
 sky130_fd_sc_hd__xnor2_2 _10216_ (.A(_03336_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__a21oi_2 _10217_ (.A1(_03206_),
    .A2(_03210_),
    .B1(_03209_),
    .Y(_03342_));
 sky130_fd_sc_hd__xnor2_1 _10218_ (.A(_03341_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2b_1 _10219_ (.A_N(_03343_),
    .B(_03335_),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_1 _10220_ (.A(_03335_),
    .B(_03343_),
    .Y(_03345_));
 sky130_fd_sc_hd__and2_1 _10221_ (.A(_03334_),
    .B(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__or2_1 _10222_ (.A(_03334_),
    .B(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__xor2_1 _10223_ (.A(_03334_),
    .B(_03345_),
    .X(_03348_));
 sky130_fd_sc_hd__xnor2_2 _10224_ (.A(_03268_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__or2_1 _10225_ (.A(_03267_),
    .B(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__and2_1 _10226_ (.A(_03267_),
    .B(_03349_),
    .X(_03351_));
 sky130_fd_sc_hd__xnor2_2 _10227_ (.A(_03267_),
    .B(_03349_),
    .Y(_03352_));
 sky130_fd_sc_hd__nor2_1 _10228_ (.A(_03085_),
    .B(_03220_),
    .Y(_03353_));
 sky130_fd_sc_hd__or4_1 _10229_ (.A(_02788_),
    .B(_02942_),
    .C(_03085_),
    .D(_03220_),
    .X(_03354_));
 sky130_fd_sc_hd__or3_1 _10230_ (.A(_02236_),
    .B(_02789_),
    .C(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__a21o_1 _10231_ (.A1(_02790_),
    .A2(_02791_),
    .B1(_03354_),
    .X(_03356_));
 sky130_fd_sc_hd__a21oi_1 _10232_ (.A1(_03083_),
    .A2(_03218_),
    .B1(_03219_),
    .Y(_03357_));
 sky130_fd_sc_hd__a21oi_1 _10233_ (.A1(_03086_),
    .A2(_03353_),
    .B1(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__o21ai_1 _10234_ (.A1(_02792_),
    .A2(_03354_),
    .B1(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__xnor2_2 _10235_ (.A(_03352_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__a21oi_1 _10236_ (.A1(_03266_),
    .A2(_03360_),
    .B1(_02242_),
    .Y(_03361_));
 sky130_fd_sc_hd__o21a_1 _10237_ (.A1(_03266_),
    .A2(_03360_),
    .B1(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__a21oi_1 _10238_ (.A1(net151),
    .A2(_02176_),
    .B1(_02177_),
    .Y(_03363_));
 sky130_fd_sc_hd__a311oi_1 _10239_ (.A1(net151),
    .A2(_02176_),
    .A3(_02177_),
    .B1(_02318_),
    .C1(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__a21oi_1 _10240_ (.A1(_06295_),
    .A2(_03232_),
    .B1(_06296_),
    .Y(_03365_));
 sky130_fd_sc_hd__mux2_1 _10241_ (.A0(_06346_),
    .A1(_03365_),
    .S(net298),
    .X(_03366_));
 sky130_fd_sc_hd__a21oi_1 _10242_ (.A1(_06292_),
    .A2(_03366_),
    .B1(net241),
    .Y(_03367_));
 sky130_fd_sc_hd__o21a_1 _10243_ (.A1(_06292_),
    .A2(_03366_),
    .B1(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__o21a_1 _10244_ (.A1(net222),
    .A2(_02293_),
    .B1(_02345_),
    .X(_03369_));
 sky130_fd_sc_hd__o21a_1 _10245_ (.A1(net226),
    .A2(_03369_),
    .B1(_02338_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(_02799_),
    .A1(_02801_),
    .S(net221),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _10247_ (.A0(_02802_),
    .A1(_02807_),
    .S(net220),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(_03371_),
    .A1(_03372_),
    .S(net222),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(_02805_),
    .A1(_02808_),
    .S(_06321_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(_02343_),
    .A1(_03374_),
    .S(net224),
    .X(_03375_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(_03373_),
    .A1(_03375_),
    .S(net226),
    .X(_03376_));
 sky130_fd_sc_hd__or2_1 _10252_ (.A(\div_res[6] ),
    .B(_03245_),
    .X(_03377_));
 sky130_fd_sc_hd__a21oi_1 _10253_ (.A1(net152),
    .A2(_03377_),
    .B1(\div_res[7] ),
    .Y(_03378_));
 sky130_fd_sc_hd__a31o_1 _10254_ (.A1(\div_res[7] ),
    .A2(net152),
    .A3(_03377_),
    .B1(net198),
    .X(_03379_));
 sky130_fd_sc_hd__o2bb2a_1 _10255_ (.A1_N(_06289_),
    .A2_N(_06455_),
    .B1(net237),
    .B2(reg1_val[7]),
    .X(_03380_));
 sky130_fd_sc_hd__or2_1 _10256_ (.A(\div_shifter[38] ),
    .B(_03248_),
    .X(_03381_));
 sky130_fd_sc_hd__a21oi_1 _10257_ (.A1(net235),
    .A2(_03381_),
    .B1(\div_shifter[39] ),
    .Y(_03382_));
 sky130_fd_sc_hd__a31o_1 _10258_ (.A1(\div_shifter[39] ),
    .A2(net235),
    .A3(_03381_),
    .B1(net239),
    .X(_03383_));
 sky130_fd_sc_hd__o22a_1 _10259_ (.A1(_06291_),
    .A2(net200),
    .B1(_03382_),
    .B2(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__o211a_1 _10260_ (.A1(_06290_),
    .A2(_02323_),
    .B1(_03380_),
    .C1(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__o221a_1 _10261_ (.A1(_06292_),
    .A2(_02327_),
    .B1(_03378_),
    .B2(_03379_),
    .C1(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__o21a_1 _10262_ (.A1(_03254_),
    .A2(_03255_),
    .B1(_03256_),
    .X(_03387_));
 sky130_fd_sc_hd__nor2_1 _10263_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03388_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2b_1 _10265_ (.A_N(_03388_),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__xnor2_1 _10266_ (.A(_03387_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__o31ai_1 _10267_ (.A1(net229),
    .A2(net209),
    .A3(_03391_),
    .B1(_03386_),
    .Y(_03392_));
 sky130_fd_sc_hd__a221o_1 _10268_ (.A1(net246),
    .A2(_03370_),
    .B1(_03376_),
    .B2(_02964_),
    .C1(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__or4_2 _10269_ (.A(_03362_),
    .B(_03364_),
    .C(_03368_),
    .D(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__or2_1 _10270_ (.A(curr_PC[7]),
    .B(_03264_),
    .X(_03395_));
 sky130_fd_sc_hd__a21oi_1 _10271_ (.A1(curr_PC[7]),
    .A2(_03264_),
    .B1(net253),
    .Y(_03396_));
 sky130_fd_sc_hd__a22o_4 _10272_ (.A1(net253),
    .A2(_03394_),
    .B1(_03395_),
    .B2(_03396_),
    .X(dest_val[7]));
 sky130_fd_sc_hd__nand4b_2 _10273_ (.A_N(_03360_),
    .B(_03226_),
    .C(_02793_),
    .D(_02688_),
    .Y(_03397_));
 sky130_fd_sc_hd__o21a_1 _10274_ (.A1(_03127_),
    .A2(_03397_),
    .B1(net151),
    .X(_03398_));
 sky130_fd_sc_hd__a21oi_2 _10275_ (.A1(_03268_),
    .A2(_03347_),
    .B1(_03346_),
    .Y(_03399_));
 sky130_fd_sc_hd__o21ai_4 _10276_ (.A1(_03341_),
    .A2(_03342_),
    .B1(_03344_),
    .Y(_03400_));
 sky130_fd_sc_hd__o22a_1 _10277_ (.A1(_00409_),
    .A2(net124),
    .B1(net122),
    .B2(net7),
    .X(_03401_));
 sky130_fd_sc_hd__xnor2_1 _10278_ (.A(net43),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__o22a_1 _10279_ (.A1(net28),
    .A2(net83),
    .B1(net81),
    .B2(_00231_),
    .X(_03403_));
 sky130_fd_sc_hd__xor2_1 _10280_ (.A(net68),
    .B(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__and3_1 _10281_ (.A(_06502_),
    .B(net43),
    .C(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__a21oi_1 _10282_ (.A1(_06502_),
    .A2(net43),
    .B1(_03404_),
    .Y(_03406_));
 sky130_fd_sc_hd__nor2_1 _10283_ (.A(_03405_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__xnor2_1 _10284_ (.A(_03402_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__o21ai_1 _10285_ (.A1(_03307_),
    .A2(_03309_),
    .B1(_03306_),
    .Y(_03409_));
 sky130_fd_sc_hd__o21ba_1 _10286_ (.A1(_03280_),
    .A2(_03282_),
    .B1_N(_03279_),
    .X(_03410_));
 sky130_fd_sc_hd__o22a_1 _10287_ (.A1(net103),
    .A2(net20),
    .B1(net18),
    .B2(net107),
    .X(_03411_));
 sky130_fd_sc_hd__xnor2_1 _10288_ (.A(_00146_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__a21oi_1 _10289_ (.A1(_00204_),
    .A2(net10),
    .B1(net186),
    .Y(_03413_));
 sky130_fd_sc_hd__a31o_2 _10290_ (.A1(net186),
    .A2(_00203_),
    .A3(net10),
    .B1(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__or2_1 _10291_ (.A(_03412_),
    .B(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__nand2_1 _10292_ (.A(_03412_),
    .B(_03414_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__and2b_1 _10294_ (.A_N(_03410_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__xnor2_1 _10295_ (.A(_03410_),
    .B(_03417_),
    .Y(_03419_));
 sky130_fd_sc_hd__and2_1 _10296_ (.A(_03409_),
    .B(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__xor2_1 _10297_ (.A(_03409_),
    .B(_03419_),
    .X(_03421_));
 sky130_fd_sc_hd__o22a_1 _10298_ (.A1(net79),
    .A2(net108),
    .B1(net104),
    .B2(net33),
    .X(_03422_));
 sky130_fd_sc_hd__xor2_1 _10299_ (.A(net113),
    .B(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__o22a_1 _10300_ (.A1(net37),
    .A2(net93),
    .B1(net91),
    .B2(net35),
    .X(_03424_));
 sky130_fd_sc_hd__xnor2_1 _10301_ (.A(net119),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__nor2_1 _10302_ (.A(_03423_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__and2_1 _10303_ (.A(_03423_),
    .B(_03425_),
    .X(_03427_));
 sky130_fd_sc_hd__nor2_1 _10304_ (.A(_03426_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__o22a_1 _10305_ (.A1(net31),
    .A2(net100),
    .B1(net57),
    .B2(net30),
    .X(_03429_));
 sky130_fd_sc_hd__xnor2_1 _10306_ (.A(net118),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__and2_1 _10307_ (.A(_03428_),
    .B(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__nor2_1 _10308_ (.A(_03428_),
    .B(_03430_),
    .Y(_03432_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(_03431_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _10310_ (.A(_03421_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__xnor2_1 _10311_ (.A(_03421_),
    .B(_03433_),
    .Y(_03435_));
 sky130_fd_sc_hd__xor2_1 _10312_ (.A(_03408_),
    .B(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__o21ba_1 _10313_ (.A1(_03325_),
    .A2(_03328_),
    .B1_N(_03324_),
    .X(_03437_));
 sky130_fd_sc_hd__o22a_1 _10314_ (.A1(net24),
    .A2(net98),
    .B1(net56),
    .B2(net22),
    .X(_03438_));
 sky130_fd_sc_hd__xnor2_1 _10315_ (.A(net129),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__o22a_1 _10316_ (.A1(net61),
    .A2(net95),
    .B1(net54),
    .B2(net58),
    .X(_03440_));
 sky130_fd_sc_hd__xnor2_1 _10317_ (.A(net126),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__xnor2_1 _10318_ (.A(_03439_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__a21oi_1 _10319_ (.A1(_03291_),
    .A2(_03295_),
    .B1(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__and3_1 _10320_ (.A(_03291_),
    .B(_03295_),
    .C(_03442_),
    .X(_03444_));
 sky130_fd_sc_hd__nor2_1 _10321_ (.A(_03443_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__and2b_1 _10322_ (.A_N(_03437_),
    .B(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__xnor2_1 _10323_ (.A(_03437_),
    .B(_03445_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _10324_ (.A(_03436_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__or2_1 _10325_ (.A(_03436_),
    .B(_03447_),
    .X(_03449_));
 sky130_fd_sc_hd__nand2_2 _10326_ (.A(_03448_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__a31o_1 _10327_ (.A1(_03149_),
    .A2(_03151_),
    .A3(_03285_),
    .B1(_03284_),
    .X(_03451_));
 sky130_fd_sc_hd__o22a_1 _10328_ (.A1(_00246_),
    .A2(net52),
    .B1(net50),
    .B2(net63),
    .X(_03452_));
 sky130_fd_sc_hd__xnor2_1 _10329_ (.A(net88),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__o22a_1 _10330_ (.A1(net71),
    .A2(net47),
    .B1(net11),
    .B2(net70),
    .X(_03454_));
 sky130_fd_sc_hd__xnor2_1 _10331_ (.A(net112),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__and2_1 _10332_ (.A(_03453_),
    .B(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__nor2_1 _10333_ (.A(_03453_),
    .B(_03455_),
    .Y(_03457_));
 sky130_fd_sc_hd__nor2_1 _10334_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__o22a_1 _10335_ (.A1(net77),
    .A2(net48),
    .B1(net13),
    .B2(net74),
    .X(_03459_));
 sky130_fd_sc_hd__xnor2_2 _10336_ (.A(net87),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__xnor2_2 _10337_ (.A(_03458_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__o21a_1 _10338_ (.A1(_03273_),
    .A2(_03274_),
    .B1(_03271_),
    .X(_03462_));
 sky130_fd_sc_hd__nor2_1 _10339_ (.A(_03461_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__xor2_2 _10340_ (.A(_03461_),
    .B(_03462_),
    .X(_03464_));
 sky130_fd_sc_hd__xnor2_2 _10341_ (.A(_03451_),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__xor2_2 _10342_ (.A(_03450_),
    .B(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__o21ai_1 _10343_ (.A1(_03318_),
    .A2(_03333_),
    .B1(_03316_),
    .Y(_03467_));
 sky130_fd_sc_hd__a21o_1 _10344_ (.A1(_03319_),
    .A2(_03332_),
    .B1(_03330_),
    .X(_03468_));
 sky130_fd_sc_hd__o21ai_2 _10345_ (.A1(_03275_),
    .A2(_03299_),
    .B1(_03298_),
    .Y(_03469_));
 sky130_fd_sc_hd__nor2_1 _10346_ (.A(_03311_),
    .B(_03314_),
    .Y(_03470_));
 sky130_fd_sc_hd__o21a_1 _10347_ (.A1(_03311_),
    .A2(_03314_),
    .B1(_03469_),
    .X(_03471_));
 sky130_fd_sc_hd__xnor2_2 _10348_ (.A(_03469_),
    .B(_03470_),
    .Y(_03472_));
 sky130_fd_sc_hd__xnor2_2 _10349_ (.A(_03468_),
    .B(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__a21oi_2 _10350_ (.A1(_03336_),
    .A2(_03340_),
    .B1(_03339_),
    .Y(_03474_));
 sky130_fd_sc_hd__xnor2_1 _10351_ (.A(_03473_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand2b_1 _10352_ (.A_N(_03475_),
    .B(_03467_),
    .Y(_03476_));
 sky130_fd_sc_hd__xnor2_1 _10353_ (.A(_03467_),
    .B(_03475_),
    .Y(_03477_));
 sky130_fd_sc_hd__and2_1 _10354_ (.A(_03466_),
    .B(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__or2_1 _10355_ (.A(_03466_),
    .B(_03477_),
    .X(_03479_));
 sky130_fd_sc_hd__xor2_1 _10356_ (.A(_03466_),
    .B(_03477_),
    .X(_03480_));
 sky130_fd_sc_hd__xnor2_2 _10357_ (.A(_03400_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__or2_1 _10358_ (.A(_03399_),
    .B(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__and2_1 _10359_ (.A(_03399_),
    .B(_03481_),
    .X(_03483_));
 sky130_fd_sc_hd__xnor2_2 _10360_ (.A(_03399_),
    .B(_03481_),
    .Y(_03484_));
 sky130_fd_sc_hd__nor2_1 _10361_ (.A(_03220_),
    .B(_03352_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(_03221_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__a21oi_1 _10363_ (.A1(_03218_),
    .A2(_03350_),
    .B1(_03351_),
    .Y(_03487_));
 sky130_fd_sc_hd__a21o_1 _10364_ (.A1(_03223_),
    .A2(_03485_),
    .B1(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__o21ba_1 _10365_ (.A1(_02945_),
    .A2(_03486_),
    .B1_N(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__xor2_2 _10366_ (.A(_03484_),
    .B(_03489_),
    .X(_03490_));
 sky130_fd_sc_hd__a21oi_1 _10367_ (.A1(_03398_),
    .A2(_03490_),
    .B1(_02242_),
    .Y(_03491_));
 sky130_fd_sc_hd__o21a_1 _10368_ (.A1(_03398_),
    .A2(_03490_),
    .B1(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__o21ai_1 _10369_ (.A1(net149),
    .A2(_02178_),
    .B1(_02179_),
    .Y(_03493_));
 sky130_fd_sc_hd__or3_1 _10370_ (.A(net149),
    .B(_02178_),
    .C(_02179_),
    .X(_03494_));
 sky130_fd_sc_hd__o21ai_1 _10371_ (.A1(_06290_),
    .A2(_03365_),
    .B1(_06291_),
    .Y(_03495_));
 sky130_fd_sc_hd__mux2_1 _10372_ (.A0(_06348_),
    .A1(_03495_),
    .S(net297),
    .X(_03496_));
 sky130_fd_sc_hd__nand2_1 _10373_ (.A(_06287_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__o211a_1 _10374_ (.A1(_06287_),
    .A2(_03496_),
    .B1(_03497_),
    .C1(net242),
    .X(_03498_));
 sky130_fd_sc_hd__o21ai_1 _10375_ (.A1(\div_res[7] ),
    .A2(_03377_),
    .B1(net152),
    .Y(_03499_));
 sky130_fd_sc_hd__xnor2_1 _10376_ (.A(\div_res[8] ),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__nor2_1 _10377_ (.A(reg1_val[8]),
    .B(net237),
    .Y(_03501_));
 sky130_fd_sc_hd__a221o_1 _10378_ (.A1(_06284_),
    .A2(_06455_),
    .B1(net273),
    .B2(_06285_),
    .C1(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__o21a_1 _10379_ (.A1(\div_shifter[39] ),
    .A2(_03381_),
    .B1(net235),
    .X(_03503_));
 sky130_fd_sc_hd__nor2_1 _10380_ (.A(\div_shifter[40] ),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__and2_1 _10381_ (.A(\div_shifter[40] ),
    .B(_03503_),
    .X(_03505_));
 sky130_fd_sc_hd__o32a_1 _10382_ (.A1(_02333_),
    .A2(_03504_),
    .A3(_03505_),
    .B1(net200),
    .B2(_06286_),
    .X(_03506_));
 sky130_fd_sc_hd__inv_2 _10383_ (.A(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__a211o_1 _10384_ (.A1(_06287_),
    .A2(net240),
    .B1(_03502_),
    .C1(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_1 _10385_ (.A0(_02277_),
    .A1(_02308_),
    .S(net222),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _10386_ (.A0(_03369_),
    .A1(_03509_),
    .S(net225),
    .X(_03510_));
 sky130_fd_sc_hd__a221o_1 _10387_ (.A1(_02330_),
    .A2(_03500_),
    .B1(_03510_),
    .B2(_02964_),
    .C1(_03508_),
    .X(_03511_));
 sky130_fd_sc_hd__o21a_1 _10388_ (.A1(_03387_),
    .A2(_03388_),
    .B1(_03389_),
    .X(_03512_));
 sky130_fd_sc_hd__nor2_1 _10389_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_1 _10390_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2b_1 _10391_ (.A_N(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__xor2_1 _10392_ (.A(_03512_),
    .B(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__o21a_1 _10393_ (.A1(net226),
    .A2(_03375_),
    .B1(_02338_),
    .X(_03517_));
 sky130_fd_sc_hd__a32o_1 _10394_ (.A1(net260),
    .A2(net210),
    .A3(_03516_),
    .B1(_03517_),
    .B2(net246),
    .X(_03518_));
 sky130_fd_sc_hd__or3_1 _10395_ (.A(_03498_),
    .B(_03511_),
    .C(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__a311o_1 _10396_ (.A1(_02317_),
    .A2(_03493_),
    .A3(_03494_),
    .B1(_03519_),
    .C1(_03492_),
    .X(_03520_));
 sky130_fd_sc_hd__and3_1 _10397_ (.A(curr_PC[7]),
    .B(curr_PC[8]),
    .C(_03264_),
    .X(_03521_));
 sky130_fd_sc_hd__a21oi_1 _10398_ (.A1(curr_PC[7]),
    .A2(_03264_),
    .B1(curr_PC[8]),
    .Y(_03522_));
 sky130_fd_sc_hd__nor2_1 _10399_ (.A(_03521_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__mux2_8 _10400_ (.A0(_03520_),
    .A1(_03523_),
    .S(net258),
    .X(dest_val[8]));
 sky130_fd_sc_hd__xor2_1 _10401_ (.A(curr_PC[9]),
    .B(_03521_),
    .X(_03524_));
 sky130_fd_sc_hd__nor3_1 _10402_ (.A(_03127_),
    .B(_03397_),
    .C(_03490_),
    .Y(_03525_));
 sky130_fd_sc_hd__or2_1 _10403_ (.A(net148),
    .B(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__a21oi_4 _10404_ (.A1(_03400_),
    .A2(_03479_),
    .B1(_03478_),
    .Y(_03527_));
 sky130_fd_sc_hd__o21ai_4 _10405_ (.A1(_03473_),
    .A2(_03474_),
    .B1(_03476_),
    .Y(_03528_));
 sky130_fd_sc_hd__o22a_1 _10406_ (.A1(net63),
    .A2(net48),
    .B1(net13),
    .B2(net78),
    .X(_03529_));
 sky130_fd_sc_hd__xnor2_1 _10407_ (.A(net87),
    .B(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__inv_2 _10408_ (.A(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__o22a_1 _10409_ (.A1(net22),
    .A2(net95),
    .B1(net54),
    .B2(net60),
    .X(_03532_));
 sky130_fd_sc_hd__xnor2_1 _10410_ (.A(net126),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__xnor2_1 _10411_ (.A(_03530_),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__o22a_1 _10412_ (.A1(net59),
    .A2(net52),
    .B1(net50),
    .B2(net64),
    .X(_03535_));
 sky130_fd_sc_hd__xnor2_1 _10413_ (.A(net88),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _10414_ (.A(_03534_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__or2_1 _10415_ (.A(_03534_),
    .B(_03536_),
    .X(_03538_));
 sky130_fd_sc_hd__and2_1 _10416_ (.A(_03537_),
    .B(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__a21o_1 _10417_ (.A1(_03402_),
    .A2(_03407_),
    .B1(_03405_),
    .X(_03540_));
 sky130_fd_sc_hd__xor2_1 _10418_ (.A(_03539_),
    .B(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__o21ai_1 _10419_ (.A1(_03418_),
    .A2(_03420_),
    .B1(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__or3_1 _10420_ (.A(_03418_),
    .B(_03420_),
    .C(_03541_),
    .X(_03543_));
 sky130_fd_sc_hd__and2_1 _10421_ (.A(_03542_),
    .B(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__o22a_1 _10422_ (.A1(net27),
    .A2(net91),
    .B1(net83),
    .B2(net25),
    .X(_03545_));
 sky130_fd_sc_hd__xnor2_1 _10423_ (.A(net67),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__o22a_1 _10424_ (.A1(net16),
    .A2(net81),
    .B1(net124),
    .B2(net7),
    .X(_03547_));
 sky130_fd_sc_hd__xnor2_1 _10425_ (.A(net43),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__o22a_1 _10426_ (.A1(net38),
    .A2(net57),
    .B1(net93),
    .B2(net36),
    .X(_03549_));
 sky130_fd_sc_hd__xnor2_1 _10427_ (.A(net120),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand2_1 _10428_ (.A(_03548_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__or2_1 _10429_ (.A(_03548_),
    .B(_03550_),
    .X(_03552_));
 sky130_fd_sc_hd__and2_1 _10430_ (.A(_03551_),
    .B(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__nand2b_1 _10431_ (.A_N(_03546_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__xnor2_1 _10432_ (.A(_03546_),
    .B(_03553_),
    .Y(_03555_));
 sky130_fd_sc_hd__or4_1 _10433_ (.A(net122),
    .B(net40),
    .C(_03439_),
    .D(_03441_),
    .X(_03556_));
 sky130_fd_sc_hd__a2bb2o_1 _10434_ (.A1_N(_03439_),
    .A2_N(_03441_),
    .B1(_00457_),
    .B2(net43),
    .X(_03557_));
 sky130_fd_sc_hd__and3_1 _10435_ (.A(_03415_),
    .B(_03556_),
    .C(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__a21oi_1 _10436_ (.A1(_03556_),
    .A2(_03557_),
    .B1(_03415_),
    .Y(_03559_));
 sky130_fd_sc_hd__o22a_1 _10437_ (.A1(net32),
    .A2(net104),
    .B1(net100),
    .B2(net29),
    .X(_03560_));
 sky130_fd_sc_hd__xnor2_2 _10438_ (.A(net116),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__o22a_1 _10439_ (.A1(net74),
    .A2(net47),
    .B1(net11),
    .B2(net71),
    .X(_03562_));
 sky130_fd_sc_hd__xnor2_2 _10440_ (.A(net112),
    .B(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__and2_1 _10441_ (.A(_03561_),
    .B(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__xor2_2 _10442_ (.A(_03561_),
    .B(_03563_),
    .X(_03565_));
 sky130_fd_sc_hd__o22a_1 _10443_ (.A1(net33),
    .A2(net108),
    .B1(net70),
    .B2(net79),
    .X(_03566_));
 sky130_fd_sc_hd__xnor2_2 _10444_ (.A(net113),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_1 _10445_ (.A(_03565_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__or3_2 _10446_ (.A(_03558_),
    .B(_03559_),
    .C(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__o21ai_1 _10447_ (.A1(_03558_),
    .A2(_03559_),
    .B1(_03568_),
    .Y(_03570_));
 sky130_fd_sc_hd__and3_1 _10448_ (.A(_03555_),
    .B(_03569_),
    .C(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__inv_2 _10449_ (.A(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__a21oi_1 _10450_ (.A1(_03569_),
    .A2(_03570_),
    .B1(_03555_),
    .Y(_03573_));
 sky130_fd_sc_hd__a21o_1 _10451_ (.A1(_03458_),
    .A2(_03460_),
    .B1(_03456_),
    .X(_03574_));
 sky130_fd_sc_hd__o22a_1 _10452_ (.A1(net103),
    .A2(net18),
    .B1(net9),
    .B2(net107),
    .X(_03575_));
 sky130_fd_sc_hd__xnor2_2 _10453_ (.A(_00146_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__inv_2 _10454_ (.A(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__o22a_1 _10455_ (.A1(net24),
    .A2(net56),
    .B1(net20),
    .B2(net98),
    .X(_03578_));
 sky130_fd_sc_hd__xnor2_2 _10456_ (.A(net129),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__and2b_1 _10457_ (.A_N(_03579_),
    .B(net186),
    .X(_03580_));
 sky130_fd_sc_hd__xor2_2 _10458_ (.A(net186),
    .B(_03579_),
    .X(_03581_));
 sky130_fd_sc_hd__xnor2_2 _10459_ (.A(_03576_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__o21a_1 _10460_ (.A1(_03426_),
    .A2(_03431_),
    .B1(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__nor3_1 _10461_ (.A(_03426_),
    .B(_03431_),
    .C(_03582_),
    .Y(_03584_));
 sky130_fd_sc_hd__nor2_1 _10462_ (.A(_03583_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__xnor2_1 _10463_ (.A(_03574_),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__or3_1 _10464_ (.A(_03571_),
    .B(_03573_),
    .C(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__o21ai_1 _10465_ (.A1(_03571_),
    .A2(_03573_),
    .B1(_03586_),
    .Y(_03588_));
 sky130_fd_sc_hd__and3_1 _10466_ (.A(_03544_),
    .B(_03587_),
    .C(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__a21oi_1 _10467_ (.A1(_03587_),
    .A2(_03588_),
    .B1(_03544_),
    .Y(_03590_));
 sky130_fd_sc_hd__nor2_2 _10468_ (.A(_03589_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__o21ai_4 _10469_ (.A1(_03450_),
    .A2(_03465_),
    .B1(_03448_),
    .Y(_03592_));
 sky130_fd_sc_hd__a21o_2 _10470_ (.A1(_03468_),
    .A2(_03472_),
    .B1(_03471_),
    .X(_03593_));
 sky130_fd_sc_hd__a21o_2 _10471_ (.A1(_03451_),
    .A2(_03464_),
    .B1(_03463_),
    .X(_03594_));
 sky130_fd_sc_hd__o21a_2 _10472_ (.A1(_03408_),
    .A2(_03435_),
    .B1(_03434_),
    .X(_03595_));
 sky130_fd_sc_hd__nor2_2 _10473_ (.A(_03443_),
    .B(_03446_),
    .Y(_03596_));
 sky130_fd_sc_hd__nor2_1 _10474_ (.A(_03595_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__xor2_4 _10475_ (.A(_03595_),
    .B(_03596_),
    .X(_03598_));
 sky130_fd_sc_hd__xor2_4 _10476_ (.A(_03594_),
    .B(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__xnor2_4 _10477_ (.A(_03593_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__and2b_1 _10478_ (.A_N(_03600_),
    .B(_03592_),
    .X(_03601_));
 sky130_fd_sc_hd__xnor2_4 _10479_ (.A(_03592_),
    .B(_03600_),
    .Y(_03602_));
 sky130_fd_sc_hd__and2_1 _10480_ (.A(_03591_),
    .B(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__xor2_4 _10481_ (.A(_03591_),
    .B(_03602_),
    .X(_03604_));
 sky130_fd_sc_hd__xnor2_4 _10482_ (.A(_03528_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__or2_1 _10483_ (.A(_03527_),
    .B(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__and2_1 _10484_ (.A(_03527_),
    .B(_03605_),
    .X(_03607_));
 sky130_fd_sc_hd__xnor2_4 _10485_ (.A(_03527_),
    .B(_03605_),
    .Y(_03608_));
 sky130_fd_sc_hd__nor2_1 _10486_ (.A(_03352_),
    .B(_03484_),
    .Y(_03609_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_03353_),
    .B(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__a21oi_1 _10488_ (.A1(_03350_),
    .A2(_03482_),
    .B1(_03483_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21o_1 _10489_ (.A1(_03357_),
    .A2(_03609_),
    .B1(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__o21ba_1 _10490_ (.A1(_03088_),
    .A2(_03610_),
    .B1_N(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__xnor2_4 _10491_ (.A(_03608_),
    .B(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__a21oi_1 _10492_ (.A1(_03526_),
    .A2(_03614_),
    .B1(_02242_),
    .Y(_03615_));
 sky130_fd_sc_hd__o21a_1 _10493_ (.A1(_03526_),
    .A2(_03614_),
    .B1(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__o21ai_1 _10494_ (.A1(net149),
    .A2(_02180_),
    .B1(_02182_),
    .Y(_03617_));
 sky130_fd_sc_hd__o31a_1 _10495_ (.A1(net149),
    .A2(_02180_),
    .A3(_02182_),
    .B1(_02317_),
    .X(_03618_));
 sky130_fd_sc_hd__a21boi_1 _10496_ (.A1(_06285_),
    .A2(_03495_),
    .B1_N(_06286_),
    .Y(_03619_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(_06350_),
    .A1(_03619_),
    .S(_04563_),
    .X(_03620_));
 sky130_fd_sc_hd__nor2_1 _10498_ (.A(_06282_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__a211o_1 _10499_ (.A1(_06282_),
    .A2(_03620_),
    .B1(_03621_),
    .C1(net241),
    .X(_03622_));
 sky130_fd_sc_hd__o21a_1 _10500_ (.A1(_03512_),
    .A2(_03513_),
    .B1(_03514_),
    .X(_03623_));
 sky130_fd_sc_hd__nor2_1 _10501_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_1 _10502_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2b_1 _10503_ (.A_N(_03624_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__xnor2_1 _10504_ (.A(_03623_),
    .B(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(_02485_),
    .A1(_02499_),
    .S(net222),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(_03236_),
    .A1(_03628_),
    .S(net225),
    .X(_03629_));
 sky130_fd_sc_hd__inv_2 _10507_ (.A(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(_03627_),
    .A1(_03630_),
    .S(net229),
    .X(_03631_));
 sky130_fd_sc_hd__or3_1 _10509_ (.A(\div_res[8] ),
    .B(\div_res[7] ),
    .C(_03377_),
    .X(_03632_));
 sky130_fd_sc_hd__a21oi_1 _10510_ (.A1(net152),
    .A2(_03632_),
    .B1(\div_res[9] ),
    .Y(_03633_));
 sky130_fd_sc_hd__a311o_1 _10511_ (.A1(\div_res[9] ),
    .A2(net152),
    .A3(_03632_),
    .B1(_03633_),
    .C1(net198),
    .X(_03634_));
 sky130_fd_sc_hd__o221a_1 _10512_ (.A1(_06279_),
    .A2(net252),
    .B1(net237),
    .B2(reg1_val[9]),
    .C1(net257),
    .X(_03635_));
 sky130_fd_sc_hd__o221a_1 _10513_ (.A1(_06281_),
    .A2(net200),
    .B1(_02323_),
    .B2(_06280_),
    .C1(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__or3_1 _10514_ (.A(\div_shifter[40] ),
    .B(\div_shifter[39] ),
    .C(_03381_),
    .X(_03637_));
 sky130_fd_sc_hd__a21oi_1 _10515_ (.A1(net235),
    .A2(_03637_),
    .B1(\div_shifter[41] ),
    .Y(_03638_));
 sky130_fd_sc_hd__a311o_1 _10516_ (.A1(\div_shifter[41] ),
    .A2(net235),
    .A3(_03637_),
    .B1(_03638_),
    .C1(net239),
    .X(_03639_));
 sky130_fd_sc_hd__o2111a_1 _10517_ (.A1(_06282_),
    .A2(_02327_),
    .B1(_03634_),
    .C1(_03636_),
    .D1(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__o21ai_1 _10518_ (.A1(net226),
    .A2(_03242_),
    .B1(_02338_),
    .Y(_03641_));
 sky130_fd_sc_hd__o221a_1 _10519_ (.A1(_02316_),
    .A2(_03630_),
    .B1(_03641_),
    .B2(_02247_),
    .C1(_03640_),
    .X(_03642_));
 sky130_fd_sc_hd__o211a_1 _10520_ (.A1(net209),
    .A2(_03631_),
    .B1(_03642_),
    .C1(_03622_),
    .X(_03643_));
 sky130_fd_sc_hd__a21bo_1 _10521_ (.A1(_03617_),
    .A2(_03618_),
    .B1_N(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__o22a_4 _10522_ (.A1(net253),
    .A2(_03524_),
    .B1(_03616_),
    .B2(_03644_),
    .X(dest_val[9]));
 sky130_fd_sc_hd__nor4b_1 _10523_ (.A(_03127_),
    .B(_03397_),
    .C(_03490_),
    .D_N(_03614_),
    .Y(_03645_));
 sky130_fd_sc_hd__nand2_2 _10524_ (.A(_03525_),
    .B(_03614_),
    .Y(_03646_));
 sky130_fd_sc_hd__a21oi_4 _10525_ (.A1(_03528_),
    .A2(_03604_),
    .B1(_03603_),
    .Y(_03647_));
 sky130_fd_sc_hd__a21o_2 _10526_ (.A1(_03593_),
    .A2(_03599_),
    .B1(_03601_),
    .X(_03648_));
 sky130_fd_sc_hd__nor2_2 _10527_ (.A(net103),
    .B(net9),
    .Y(_03649_));
 sky130_fd_sc_hd__xnor2_4 _10528_ (.A(net173),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21oi_4 _10529_ (.A1(_03565_),
    .A2(_03567_),
    .B1(_03564_),
    .Y(_03651_));
 sky130_fd_sc_hd__nor2_1 _10530_ (.A(_03650_),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__xnor2_4 _10531_ (.A(_03650_),
    .B(_03651_),
    .Y(_03653_));
 sky130_fd_sc_hd__o21a_2 _10532_ (.A1(_03531_),
    .A2(_03533_),
    .B1(_03537_),
    .X(_03654_));
 sky130_fd_sc_hd__xnor2_4 _10533_ (.A(_03653_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o22a_1 _10534_ (.A1(net27),
    .A2(net93),
    .B1(net91),
    .B2(net26),
    .X(_03656_));
 sky130_fd_sc_hd__xnor2_1 _10535_ (.A(net67),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__o22a_1 _10536_ (.A1(net32),
    .A2(net108),
    .B1(net104),
    .B2(net29),
    .X(_03658_));
 sky130_fd_sc_hd__xor2_1 _10537_ (.A(net116),
    .B(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__nor2_1 _10538_ (.A(_03657_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__and2_1 _10539_ (.A(_03657_),
    .B(_03659_),
    .X(_03661_));
 sky130_fd_sc_hd__or2_1 _10540_ (.A(_03660_),
    .B(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__a2bb2o_1 _10541_ (.A1_N(net36),
    .A2_N(net57),
    .B1(net99),
    .B2(_06486_),
    .X(_03663_));
 sky130_fd_sc_hd__xnor2_1 _10542_ (.A(_06472_),
    .B(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__and2b_1 _10543_ (.A_N(_03662_),
    .B(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__and2b_1 _10544_ (.A_N(_03664_),
    .B(_03662_),
    .X(_03666_));
 sky130_fd_sc_hd__or2_2 _10545_ (.A(_03665_),
    .B(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__o21ba_2 _10546_ (.A1(_03577_),
    .A2(_03581_),
    .B1_N(_03580_),
    .X(_03668_));
 sky130_fd_sc_hd__o22a_2 _10547_ (.A1(net16),
    .A2(net83),
    .B1(net81),
    .B2(net7),
    .X(_03669_));
 sky130_fd_sc_hd__xnor2_4 _10548_ (.A(net43),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__and2b_1 _10549_ (.A_N(_03668_),
    .B(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__xnor2_4 _10550_ (.A(_03668_),
    .B(_03670_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_2 _10551_ (.A(_00450_),
    .B(net43),
    .Y(_03673_));
 sky130_fd_sc_hd__xnor2_4 _10552_ (.A(_03672_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__or2_1 _10553_ (.A(net79),
    .B(net72),
    .X(_03675_));
 sky130_fd_sc_hd__a21o_1 _10554_ (.A1(_06514_),
    .A2(_06515_),
    .B1(net69),
    .X(_03676_));
 sky130_fd_sc_hd__and3_1 _10555_ (.A(net114),
    .B(_03675_),
    .C(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__a21oi_1 _10556_ (.A1(_03675_),
    .A2(_03676_),
    .B1(net114),
    .Y(_03678_));
 sky130_fd_sc_hd__or2_1 _10557_ (.A(net65),
    .B(net48),
    .X(_03679_));
 sky130_fd_sc_hd__a21o_1 _10558_ (.A1(_00438_),
    .A2(_00439_),
    .B1(net62),
    .X(_03680_));
 sky130_fd_sc_hd__and3_1 _10559_ (.A(net85),
    .B(_03679_),
    .C(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__a21oi_1 _10560_ (.A1(_03679_),
    .A2(_03680_),
    .B1(net85),
    .Y(_03682_));
 sky130_fd_sc_hd__o22a_1 _10561_ (.A1(_03677_),
    .A2(_03678_),
    .B1(_03681_),
    .B2(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__or4_1 _10562_ (.A(_03677_),
    .B(_03678_),
    .C(_03681_),
    .D(_03682_),
    .X(_03684_));
 sky130_fd_sc_hd__and2b_1 _10563_ (.A_N(_03683_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__o22a_1 _10564_ (.A1(net77),
    .A2(net46),
    .B1(net12),
    .B2(net74),
    .X(_03686_));
 sky130_fd_sc_hd__xnor2_1 _10565_ (.A(net111),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__and2_1 _10566_ (.A(_03685_),
    .B(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__nor2_1 _10567_ (.A(_03685_),
    .B(_03687_),
    .Y(_03689_));
 sky130_fd_sc_hd__nor2_2 _10568_ (.A(_03688_),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__nand2_1 _10569_ (.A(_03674_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__xnor2_4 _10570_ (.A(_03674_),
    .B(_03690_),
    .Y(_03692_));
 sky130_fd_sc_hd__xor2_4 _10571_ (.A(_03667_),
    .B(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__nand2b_1 _10572_ (.A_N(_03655_),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__xnor2_4 _10573_ (.A(_03655_),
    .B(_03693_),
    .Y(_03695_));
 sky130_fd_sc_hd__a21bo_2 _10574_ (.A1(_03415_),
    .A2(_03557_),
    .B1_N(_03556_),
    .X(_03696_));
 sky130_fd_sc_hd__o22a_1 _10575_ (.A1(net56),
    .A2(net20),
    .B1(net18),
    .B2(net98),
    .X(_03697_));
 sky130_fd_sc_hd__xnor2_1 _10576_ (.A(net129),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__o22a_1 _10577_ (.A1(net61),
    .A2(net53),
    .B1(net50),
    .B2(net58),
    .X(_03699_));
 sky130_fd_sc_hd__xnor2_2 _10578_ (.A(_00388_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__or2_1 _10579_ (.A(_03698_),
    .B(_03700_),
    .X(_03701_));
 sky130_fd_sc_hd__nand2_1 _10580_ (.A(_03698_),
    .B(_03700_),
    .Y(_03702_));
 sky130_fd_sc_hd__nand2_1 _10581_ (.A(_03701_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__o22a_1 _10582_ (.A1(net24),
    .A2(net95),
    .B1(net54),
    .B2(net22),
    .X(_03704_));
 sky130_fd_sc_hd__xnor2_1 _10583_ (.A(net126),
    .B(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__xnor2_1 _10584_ (.A(_03703_),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__a21oi_1 _10585_ (.A1(_03551_),
    .A2(_03554_),
    .B1(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__and3_1 _10586_ (.A(_03551_),
    .B(_03554_),
    .C(_03706_),
    .X(_03708_));
 sky130_fd_sc_hd__nor2_2 _10587_ (.A(_03707_),
    .B(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__xor2_4 _10588_ (.A(_03696_),
    .B(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__xnor2_4 _10589_ (.A(_03695_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__a21bo_2 _10590_ (.A1(_03544_),
    .A2(_03588_),
    .B1_N(_03587_),
    .X(_03712_));
 sky130_fd_sc_hd__a21bo_2 _10591_ (.A1(_03539_),
    .A2(_03540_),
    .B1_N(_03542_),
    .X(_03713_));
 sky130_fd_sc_hd__nand2_2 _10592_ (.A(_03569_),
    .B(_03572_),
    .Y(_03714_));
 sky130_fd_sc_hd__a21oi_4 _10593_ (.A1(_03574_),
    .A2(_03585_),
    .B1(_03583_),
    .Y(_03715_));
 sky130_fd_sc_hd__a21oi_1 _10594_ (.A1(_03569_),
    .A2(_03572_),
    .B1(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__xnor2_4 _10595_ (.A(_03714_),
    .B(_03715_),
    .Y(_03717_));
 sky130_fd_sc_hd__xnor2_4 _10596_ (.A(_03713_),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__a21oi_4 _10597_ (.A1(_03594_),
    .A2(_03598_),
    .B1(_03597_),
    .Y(_03719_));
 sky130_fd_sc_hd__nor2_1 _10598_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__xor2_4 _10599_ (.A(_03718_),
    .B(_03719_),
    .X(_03721_));
 sky130_fd_sc_hd__xnor2_4 _10600_ (.A(_03712_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__nor2_1 _10601_ (.A(_03711_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__xor2_4 _10602_ (.A(_03711_),
    .B(_03722_),
    .X(_03724_));
 sky130_fd_sc_hd__xnor2_4 _10603_ (.A(_03648_),
    .B(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__or2_1 _10604_ (.A(_03647_),
    .B(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__and2_1 _10605_ (.A(_03647_),
    .B(_03725_),
    .X(_03727_));
 sky130_fd_sc_hd__xnor2_4 _10606_ (.A(_03647_),
    .B(_03725_),
    .Y(_03728_));
 sky130_fd_sc_hd__nor2_1 _10607_ (.A(_03484_),
    .B(_03608_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _10608_ (.A(_03485_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand4b_2 _10609_ (.A_N(_02944_),
    .B(_03221_),
    .C(_03485_),
    .D(_03729_),
    .Y(_03731_));
 sky130_fd_sc_hd__a21oi_1 _10610_ (.A1(_03482_),
    .A2(_03606_),
    .B1(_03607_),
    .Y(_03732_));
 sky130_fd_sc_hd__a21oi_1 _10611_ (.A1(_03487_),
    .A2(_03729_),
    .B1(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__o221ai_4 _10612_ (.A1(_03224_),
    .A2(_03730_),
    .B1(_03731_),
    .B2(_02640_),
    .C1(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__xnor2_2 _10613_ (.A(_03728_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__a21oi_1 _10614_ (.A1(net151),
    .A2(_03646_),
    .B1(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__a31o_1 _10615_ (.A1(net151),
    .A2(_03646_),
    .A3(_03735_),
    .B1(_02242_),
    .X(_03737_));
 sky130_fd_sc_hd__o21ai_1 _10616_ (.A1(net148),
    .A2(_02183_),
    .B1(_02184_),
    .Y(_03738_));
 sky130_fd_sc_hd__or3_1 _10617_ (.A(net148),
    .B(_02183_),
    .C(_02184_),
    .X(_03739_));
 sky130_fd_sc_hd__nand2_1 _10618_ (.A(_03738_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__o21a_1 _10619_ (.A1(_06280_),
    .A2(_03619_),
    .B1(_06281_),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(_06352_),
    .A1(_03741_),
    .S(net297),
    .X(_03742_));
 sky130_fd_sc_hd__nor2_1 _10621_ (.A(_06276_),
    .B(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__a211o_1 _10622_ (.A1(_06276_),
    .A2(_03742_),
    .B1(_03743_),
    .C1(net241),
    .X(_03744_));
 sky130_fd_sc_hd__nand2_1 _10623_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03745_));
 sky130_fd_sc_hd__or2_1 _10624_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _10625_ (.A(_03745_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__o21ai_1 _10626_ (.A1(_03623_),
    .A2(_03624_),
    .B1(_03625_),
    .Y(_03748_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(_02655_),
    .A1(_02661_),
    .S(net223),
    .X(_03749_));
 sky130_fd_sc_hd__inv_2 _10628_ (.A(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__mux2_1 _10629_ (.A0(_03098_),
    .A1(_03750_),
    .S(net225),
    .X(_03751_));
 sky130_fd_sc_hd__xor2_1 _10630_ (.A(_03747_),
    .B(_03748_),
    .X(_03752_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(_03751_),
    .A1(_03752_),
    .S(net261),
    .X(_03753_));
 sky130_fd_sc_hd__or2_1 _10632_ (.A(\div_res[9] ),
    .B(_03632_),
    .X(_03754_));
 sky130_fd_sc_hd__a21oi_1 _10633_ (.A1(net154),
    .A2(_03754_),
    .B1(\div_res[10] ),
    .Y(_03755_));
 sky130_fd_sc_hd__a311o_1 _10634_ (.A1(\div_res[10] ),
    .A2(net154),
    .A3(_03754_),
    .B1(_03755_),
    .C1(net198),
    .X(_03756_));
 sky130_fd_sc_hd__or2_1 _10635_ (.A(\div_shifter[41] ),
    .B(_03637_),
    .X(_03757_));
 sky130_fd_sc_hd__a21oi_1 _10636_ (.A1(net235),
    .A2(_03757_),
    .B1(\div_shifter[42] ),
    .Y(_03758_));
 sky130_fd_sc_hd__a311o_1 _10637_ (.A1(\div_shifter[42] ),
    .A2(net234),
    .A3(_03757_),
    .B1(_03758_),
    .C1(net239),
    .X(_03759_));
 sky130_fd_sc_hd__nand2_1 _10638_ (.A(_06274_),
    .B(net273),
    .Y(_03760_));
 sky130_fd_sc_hd__o221a_1 _10639_ (.A1(_06273_),
    .A2(net252),
    .B1(net236),
    .B2(reg1_val[10]),
    .C1(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__o221a_1 _10640_ (.A1(_06275_),
    .A2(net200),
    .B1(_02327_),
    .B2(_06276_),
    .C1(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__and3_1 _10641_ (.A(_03756_),
    .B(_03759_),
    .C(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__o21ai_2 _10642_ (.A1(net226),
    .A2(_03104_),
    .B1(_02338_),
    .Y(_03764_));
 sky130_fd_sc_hd__o221a_1 _10643_ (.A1(_02316_),
    .A2(_03751_),
    .B1(_03764_),
    .B2(_02247_),
    .C1(_03763_),
    .X(_03765_));
 sky130_fd_sc_hd__o211a_1 _10644_ (.A1(net209),
    .A2(_03753_),
    .B1(_03765_),
    .C1(_03744_),
    .X(_03766_));
 sky130_fd_sc_hd__o221a_2 _10645_ (.A1(_03736_),
    .A2(_03737_),
    .B1(_03740_),
    .B2(_02318_),
    .C1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__and3_1 _10646_ (.A(curr_PC[9]),
    .B(curr_PC[10]),
    .C(_03521_),
    .X(_03768_));
 sky130_fd_sc_hd__a21oi_1 _10647_ (.A1(curr_PC[9]),
    .A2(_03521_),
    .B1(curr_PC[10]),
    .Y(_03769_));
 sky130_fd_sc_hd__or3_1 _10648_ (.A(net253),
    .B(_03768_),
    .C(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__o21ai_4 _10649_ (.A1(net258),
    .A2(_03767_),
    .B1(_03770_),
    .Y(dest_val[10]));
 sky130_fd_sc_hd__o21a_1 _10650_ (.A1(_03646_),
    .A2(_03735_),
    .B1(net151),
    .X(_03771_));
 sky130_fd_sc_hd__a21o_1 _10651_ (.A1(_03648_),
    .A2(_03724_),
    .B1(_03723_),
    .X(_03772_));
 sky130_fd_sc_hd__a21o_1 _10652_ (.A1(_03712_),
    .A2(_03721_),
    .B1(_03720_),
    .X(_03773_));
 sky130_fd_sc_hd__a31o_1 _10653_ (.A1(_00450_),
    .A2(net43),
    .A3(_03672_),
    .B1(_03671_),
    .X(_03774_));
 sky130_fd_sc_hd__o22a_1 _10654_ (.A1(net56),
    .A2(net18),
    .B1(net9),
    .B2(net98),
    .X(_03775_));
 sky130_fd_sc_hd__xnor2_1 _10655_ (.A(net129),
    .B(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__o22a_1 _10656_ (.A1(net24),
    .A2(net54),
    .B1(net20),
    .B2(net95),
    .X(_03777_));
 sky130_fd_sc_hd__xnor2_1 _10657_ (.A(net126),
    .B(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__xnor2_1 _10658_ (.A(net173),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__nand2b_1 _10659_ (.A_N(_03776_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__xnor2_1 _10660_ (.A(_03776_),
    .B(_03779_),
    .Y(_03781_));
 sky130_fd_sc_hd__o21a_1 _10661_ (.A1(_03660_),
    .A2(_03665_),
    .B1(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__nor3_1 _10662_ (.A(_03660_),
    .B(_03665_),
    .C(_03781_),
    .Y(_03783_));
 sky130_fd_sc_hd__nor2_1 _10663_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__xnor2_1 _10664_ (.A(_03774_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__o22a_1 _10665_ (.A1(net37),
    .A2(net104),
    .B1(net100),
    .B2(net35),
    .X(_03786_));
 sky130_fd_sc_hd__xnor2_1 _10666_ (.A(net120),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__o22a_1 _10667_ (.A1(net79),
    .A2(net74),
    .B1(net71),
    .B2(net33),
    .X(_03788_));
 sky130_fd_sc_hd__xnor2_1 _10668_ (.A(net113),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__and2_1 _10669_ (.A(_03787_),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__xor2_1 _10670_ (.A(_03787_),
    .B(_03789_),
    .X(_03791_));
 sky130_fd_sc_hd__o22a_1 _10671_ (.A1(net29),
    .A2(net108),
    .B1(net70),
    .B2(net32),
    .X(_03792_));
 sky130_fd_sc_hd__xnor2_1 _10672_ (.A(net117),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__and2_1 _10673_ (.A(_03791_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__nor2_1 _10674_ (.A(_03791_),
    .B(_03793_),
    .Y(_03795_));
 sky130_fd_sc_hd__nor2_1 _10675_ (.A(_03794_),
    .B(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__a21o_1 _10676_ (.A1(_00267_),
    .A2(_00269_),
    .B1(net52),
    .X(_03797_));
 sky130_fd_sc_hd__or2_1 _10677_ (.A(net61),
    .B(net50),
    .X(_03798_));
 sky130_fd_sc_hd__nand3_1 _10678_ (.A(net88),
    .B(_03797_),
    .C(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__a21o_1 _10679_ (.A1(_03797_),
    .A2(_03798_),
    .B1(net88),
    .X(_03800_));
 sky130_fd_sc_hd__o32a_1 _10680_ (.A1(net77),
    .A2(_00452_),
    .A3(_00453_),
    .B1(net62),
    .B2(net46),
    .X(_03801_));
 sky130_fd_sc_hd__xnor2_1 _10681_ (.A(net110),
    .B(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__a21o_1 _10682_ (.A1(_03799_),
    .A2(_03800_),
    .B1(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__nand3_1 _10683_ (.A(_03799_),
    .B(_03800_),
    .C(_03802_),
    .Y(_03804_));
 sky130_fd_sc_hd__o22a_1 _10684_ (.A1(net58),
    .A2(net48),
    .B1(net13),
    .B2(net64),
    .X(_03805_));
 sky130_fd_sc_hd__xnor2_1 _10685_ (.A(net87),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__and3_1 _10686_ (.A(_03803_),
    .B(_03804_),
    .C(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__a21oi_1 _10687_ (.A1(_03803_),
    .A2(_03804_),
    .B1(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__nor2_1 _10688_ (.A(_03807_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__o22a_1 _10689_ (.A1(net91),
    .A2(net16),
    .B1(net83),
    .B2(net6),
    .X(_03810_));
 sky130_fd_sc_hd__xnor2_1 _10690_ (.A(net42),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__o22a_1 _10691_ (.A1(net27),
    .A2(net57),
    .B1(net93),
    .B2(net26),
    .X(_03812_));
 sky130_fd_sc_hd__xor2_1 _10692_ (.A(net66),
    .B(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__nand2_1 _10693_ (.A(_00445_),
    .B(net42),
    .Y(_03814_));
 sky130_fd_sc_hd__and3_1 _10694_ (.A(_00445_),
    .B(net42),
    .C(_03813_),
    .X(_03815_));
 sky130_fd_sc_hd__xnor2_1 _10695_ (.A(_03813_),
    .B(_03814_),
    .Y(_03816_));
 sky130_fd_sc_hd__xor2_1 _10696_ (.A(_03811_),
    .B(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_03809_),
    .B(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__or2_1 _10698_ (.A(_03809_),
    .B(_03817_),
    .X(_03819_));
 sky130_fd_sc_hd__and3_1 _10699_ (.A(_03796_),
    .B(_03818_),
    .C(_03819_),
    .X(_03820_));
 sky130_fd_sc_hd__inv_2 _10700_ (.A(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__a21o_1 _10701_ (.A1(_03818_),
    .A2(_03819_),
    .B1(_03796_),
    .X(_03822_));
 sky130_fd_sc_hd__nand2_1 _10702_ (.A(_03821_),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__o21ai_2 _10703_ (.A1(_03703_),
    .A2(_03705_),
    .B1(_03701_),
    .Y(_03824_));
 sky130_fd_sc_hd__o21a_1 _10704_ (.A1(_03683_),
    .A2(_03688_),
    .B1(_03650_),
    .X(_03825_));
 sky130_fd_sc_hd__nor3_1 _10705_ (.A(_03650_),
    .B(_03683_),
    .C(_03688_),
    .Y(_03826_));
 sky130_fd_sc_hd__nor2_1 _10706_ (.A(_03825_),
    .B(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__xnor2_2 _10707_ (.A(_03824_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__xnor2_1 _10708_ (.A(_03823_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__or2_1 _10709_ (.A(_03785_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__nand2_1 _10710_ (.A(_03785_),
    .B(_03829_),
    .Y(_03831_));
 sky130_fd_sc_hd__and2_1 _10711_ (.A(_03830_),
    .B(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__a21bo_1 _10712_ (.A1(_03695_),
    .A2(_03710_),
    .B1_N(_03694_),
    .X(_03833_));
 sky130_fd_sc_hd__a21o_1 _10713_ (.A1(_03713_),
    .A2(_03717_),
    .B1(_03716_),
    .X(_03834_));
 sky130_fd_sc_hd__a21o_1 _10714_ (.A1(_03696_),
    .A2(_03709_),
    .B1(_03707_),
    .X(_03835_));
 sky130_fd_sc_hd__o21ba_1 _10715_ (.A1(_03653_),
    .A2(_03654_),
    .B1_N(_03652_),
    .X(_03836_));
 sky130_fd_sc_hd__o21ai_2 _10716_ (.A1(_03667_),
    .A2(_03692_),
    .B1(_03691_),
    .Y(_03837_));
 sky130_fd_sc_hd__and2b_1 _10717_ (.A_N(_03836_),
    .B(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__xnor2_2 _10718_ (.A(_03836_),
    .B(_03837_),
    .Y(_03839_));
 sky130_fd_sc_hd__xor2_2 _10719_ (.A(_03835_),
    .B(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__xnor2_2 _10720_ (.A(_03834_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2b_1 _10721_ (.A_N(_03841_),
    .B(_03833_),
    .Y(_03842_));
 sky130_fd_sc_hd__xnor2_2 _10722_ (.A(_03833_),
    .B(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__and2_1 _10723_ (.A(_03832_),
    .B(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__xor2_2 _10724_ (.A(_03832_),
    .B(_03843_),
    .X(_03845_));
 sky130_fd_sc_hd__xnor2_2 _10725_ (.A(_03773_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2b_1 _10726_ (.A_N(_03846_),
    .B(_03772_),
    .Y(_03847_));
 sky130_fd_sc_hd__and2b_1 _10727_ (.A_N(_03772_),
    .B(_03846_),
    .X(_03848_));
 sky130_fd_sc_hd__xnor2_2 _10728_ (.A(_03772_),
    .B(_03846_),
    .Y(_03849_));
 sky130_fd_sc_hd__a21oi_1 _10729_ (.A1(_03606_),
    .A2(_03726_),
    .B1(_03727_),
    .Y(_03850_));
 sky130_fd_sc_hd__nor2_1 _10730_ (.A(_03608_),
    .B(_03728_),
    .Y(_03851_));
 sky130_fd_sc_hd__a21oi_2 _10731_ (.A1(_03611_),
    .A2(_03851_),
    .B1(_03850_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _10732_ (.A(_03609_),
    .B(_03851_),
    .Y(_03853_));
 sky130_fd_sc_hd__a31o_2 _10733_ (.A1(_03355_),
    .A2(_03356_),
    .A3(_03358_),
    .B1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__and3_1 _10734_ (.A(_03849_),
    .B(_03852_),
    .C(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__a21oi_1 _10735_ (.A1(_03852_),
    .A2(_03854_),
    .B1(_03849_),
    .Y(_03856_));
 sky130_fd_sc_hd__or2_1 _10736_ (.A(_03855_),
    .B(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__o21ai_1 _10737_ (.A1(_03771_),
    .A2(_03857_),
    .B1(net202),
    .Y(_03858_));
 sky130_fd_sc_hd__a21oi_1 _10738_ (.A1(_03771_),
    .A2(_03857_),
    .B1(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__o21ai_1 _10739_ (.A1(net148),
    .A2(_02185_),
    .B1(_02186_),
    .Y(_03860_));
 sky130_fd_sc_hd__or3_1 _10740_ (.A(net150),
    .B(_02185_),
    .C(_02186_),
    .X(_03861_));
 sky130_fd_sc_hd__o21ai_1 _10741_ (.A1(_06276_),
    .A2(_03741_),
    .B1(_06275_),
    .Y(_03862_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(_06354_),
    .A1(_03862_),
    .S(net297),
    .X(_03863_));
 sky130_fd_sc_hd__nor2_1 _10743_ (.A(_06269_),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__a21o_1 _10744_ (.A1(_06269_),
    .A2(_03863_),
    .B1(net241),
    .X(_03865_));
 sky130_fd_sc_hd__and2_1 _10745_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03866_));
 sky130_fd_sc_hd__nor2_1 _10746_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .Y(_03867_));
 sky130_fd_sc_hd__or2_1 _10747_ (.A(_03866_),
    .B(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__a21bo_1 _10748_ (.A1(_03746_),
    .A2(_03748_),
    .B1_N(_03745_),
    .X(_03869_));
 sky130_fd_sc_hd__and2b_1 _10749_ (.A_N(_03868_),
    .B(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(_02803_),
    .A1(_02809_),
    .S(net222),
    .X(_03871_));
 sky130_fd_sc_hd__inv_2 _10751_ (.A(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(_02956_),
    .A1(_03872_),
    .S(net225),
    .X(_03873_));
 sky130_fd_sc_hd__xor2_1 _10753_ (.A(_03868_),
    .B(_03869_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(_03873_),
    .A1(_03874_),
    .S(net261),
    .X(_03875_));
 sky130_fd_sc_hd__or2_1 _10755_ (.A(\div_res[10] ),
    .B(_03754_),
    .X(_03876_));
 sky130_fd_sc_hd__a21oi_1 _10756_ (.A1(net154),
    .A2(_03876_),
    .B1(\div_res[11] ),
    .Y(_03877_));
 sky130_fd_sc_hd__a31o_1 _10757_ (.A1(\div_res[11] ),
    .A2(net154),
    .A3(_03876_),
    .B1(net199),
    .X(_03878_));
 sky130_fd_sc_hd__or2_1 _10758_ (.A(\div_shifter[42] ),
    .B(_03757_),
    .X(_03879_));
 sky130_fd_sc_hd__a21oi_1 _10759_ (.A1(net235),
    .A2(_03879_),
    .B1(\div_shifter[43] ),
    .Y(_03880_));
 sky130_fd_sc_hd__a31o_1 _10760_ (.A1(\div_shifter[43] ),
    .A2(net235),
    .A3(_03879_),
    .B1(net239),
    .X(_03881_));
 sky130_fd_sc_hd__o21ai_1 _10761_ (.A1(reg1_val[11]),
    .A2(_06238_),
    .B1(net273),
    .Y(_03882_));
 sky130_fd_sc_hd__o221a_1 _10762_ (.A1(_06247_),
    .A2(net252),
    .B1(net236),
    .B2(reg1_val[11]),
    .C1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__a21boi_1 _10763_ (.A1(_06263_),
    .A2(net201),
    .B1_N(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__o221a_1 _10764_ (.A1(_06270_),
    .A2(_02327_),
    .B1(_03880_),
    .B2(_03881_),
    .C1(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__o21ai_2 _10765_ (.A1(net226),
    .A2(_02962_),
    .B1(_02338_),
    .Y(_03886_));
 sky130_fd_sc_hd__o221a_1 _10766_ (.A1(_03877_),
    .A2(_03878_),
    .B1(_03886_),
    .B2(_02247_),
    .C1(_03885_),
    .X(_03887_));
 sky130_fd_sc_hd__o221a_1 _10767_ (.A1(_02316_),
    .A2(_03873_),
    .B1(_03875_),
    .B2(_06447_),
    .C1(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__o21ai_1 _10768_ (.A1(_03864_),
    .A2(_03865_),
    .B1(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__a311o_2 _10769_ (.A1(_02317_),
    .A2(_03860_),
    .A3(_03861_),
    .B1(_03889_),
    .C1(_03859_),
    .X(_03890_));
 sky130_fd_sc_hd__or2_1 _10770_ (.A(curr_PC[11]),
    .B(_03768_),
    .X(_03891_));
 sky130_fd_sc_hd__and2_1 _10771_ (.A(curr_PC[11]),
    .B(_03768_),
    .X(_03892_));
 sky130_fd_sc_hd__nor2_1 _10772_ (.A(net254),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__a22o_4 _10773_ (.A1(net253),
    .A2(_03890_),
    .B1(_03891_),
    .B2(_03893_),
    .X(dest_val[11]));
 sky130_fd_sc_hd__or2_1 _10774_ (.A(_03735_),
    .B(_03857_),
    .X(_03894_));
 sky130_fd_sc_hd__o21ai_1 _10775_ (.A1(_03646_),
    .A2(_03894_),
    .B1(net151),
    .Y(_03895_));
 sky130_fd_sc_hd__inv_2 _10776_ (.A(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__a21bo_1 _10777_ (.A1(_03834_),
    .A2(_03840_),
    .B1_N(_03842_),
    .X(_03897_));
 sky130_fd_sc_hd__o22a_1 _10778_ (.A1(net27),
    .A2(net100),
    .B1(net57),
    .B2(net25),
    .X(_03898_));
 sky130_fd_sc_hd__xnor2_1 _10779_ (.A(net67),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__o22a_1 _10780_ (.A1(net93),
    .A2(net16),
    .B1(net6),
    .B2(net91),
    .X(_03900_));
 sky130_fd_sc_hd__xnor2_1 _10781_ (.A(net42),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2b_1 _10782_ (.A_N(_03899_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__xnor2_1 _10783_ (.A(_03899_),
    .B(_03901_),
    .Y(_03903_));
 sky130_fd_sc_hd__o22a_1 _10784_ (.A1(net23),
    .A2(net52),
    .B1(net50),
    .B2(net21),
    .X(_03904_));
 sky130_fd_sc_hd__xnor2_1 _10785_ (.A(net88),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__o22a_1 _10786_ (.A1(net64),
    .A2(net47),
    .B1(net11),
    .B2(net63),
    .X(_03906_));
 sky130_fd_sc_hd__xnor2_1 _10787_ (.A(net112),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_1 _10788_ (.A(_03905_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__xor2_1 _10789_ (.A(_03905_),
    .B(_03907_),
    .X(_03909_));
 sky130_fd_sc_hd__o22a_1 _10790_ (.A1(net60),
    .A2(net48),
    .B1(net13),
    .B2(net59),
    .X(_03910_));
 sky130_fd_sc_hd__xnor2_1 _10791_ (.A(net87),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand2_1 _10792_ (.A(_03909_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__xor2_1 _10793_ (.A(_03909_),
    .B(_03911_),
    .X(_03913_));
 sky130_fd_sc_hd__and2_1 _10794_ (.A(_03903_),
    .B(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__xnor2_1 _10795_ (.A(_03903_),
    .B(_03913_),
    .Y(_03915_));
 sky130_fd_sc_hd__o22a_1 _10796_ (.A1(net37),
    .A2(net108),
    .B1(net104),
    .B2(net35),
    .X(_03916_));
 sky130_fd_sc_hd__xnor2_1 _10797_ (.A(net120),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__o22a_1 _10798_ (.A1(net79),
    .A2(net78),
    .B1(net74),
    .B2(net33),
    .X(_03918_));
 sky130_fd_sc_hd__xnor2_1 _10799_ (.A(net113),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__and2_1 _10800_ (.A(_03917_),
    .B(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__nor2_1 _10801_ (.A(_03917_),
    .B(_03919_),
    .Y(_03921_));
 sky130_fd_sc_hd__nor2_1 _10802_ (.A(_03920_),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__o22a_1 _10803_ (.A1(net32),
    .A2(net71),
    .B1(net70),
    .B2(net29),
    .X(_03923_));
 sky130_fd_sc_hd__xnor2_1 _10804_ (.A(net116),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__xor2_1 _10805_ (.A(_03922_),
    .B(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__and2b_1 _10806_ (.A_N(_03915_),
    .B(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__xnor2_1 _10807_ (.A(_03915_),
    .B(_03925_),
    .Y(_03927_));
 sky130_fd_sc_hd__o21ai_2 _10808_ (.A1(_00146_),
    .A2(_03778_),
    .B1(_03780_),
    .Y(_03928_));
 sky130_fd_sc_hd__a21bo_1 _10809_ (.A1(_03804_),
    .A2(_03806_),
    .B1_N(_03803_),
    .X(_03929_));
 sky130_fd_sc_hd__nand2_1 _10810_ (.A(_00436_),
    .B(net42),
    .Y(_03930_));
 sky130_fd_sc_hd__and3_1 _10811_ (.A(_00436_),
    .B(net42),
    .C(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__xnor2_1 _10812_ (.A(_03929_),
    .B(_03930_),
    .Y(_03932_));
 sky130_fd_sc_hd__xor2_1 _10813_ (.A(_03928_),
    .B(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(_03927_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__or2_1 _10815_ (.A(_03927_),
    .B(_03933_),
    .X(_03935_));
 sky130_fd_sc_hd__nand2_1 _10816_ (.A(_03934_),
    .B(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__a21o_1 _10817_ (.A1(_03811_),
    .A2(_03816_),
    .B1(_03815_),
    .X(_03937_));
 sky130_fd_sc_hd__o22a_1 _10818_ (.A1(net54),
    .A2(net20),
    .B1(net18),
    .B2(net95),
    .X(_03938_));
 sky130_fd_sc_hd__xnor2_2 _10819_ (.A(_00319_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__a21oi_1 _10820_ (.A1(_00303_),
    .A2(_00567_),
    .B1(net130),
    .Y(_03940_));
 sky130_fd_sc_hd__a31o_2 _10821_ (.A1(net130),
    .A2(_00304_),
    .A3(_00567_),
    .B1(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__xnor2_1 _10822_ (.A(_03939_),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__o21ai_1 _10823_ (.A1(_03790_),
    .A2(_03794_),
    .B1(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__or3_1 _10824_ (.A(_03790_),
    .B(_03794_),
    .C(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__and2_1 _10825_ (.A(_03943_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__xnor2_1 _10826_ (.A(_03937_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__xor2_1 _10827_ (.A(_03936_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__o21ai_2 _10828_ (.A1(_03823_),
    .A2(_03828_),
    .B1(_03830_),
    .Y(_03948_));
 sky130_fd_sc_hd__a21o_1 _10829_ (.A1(_03774_),
    .A2(_03784_),
    .B1(_03782_),
    .X(_03949_));
 sky130_fd_sc_hd__a21oi_1 _10830_ (.A1(_03824_),
    .A2(_03827_),
    .B1(_03825_),
    .Y(_03950_));
 sky130_fd_sc_hd__a21oi_1 _10831_ (.A1(_03818_),
    .A2(_03821_),
    .B1(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand3_1 _10832_ (.A(_03818_),
    .B(_03821_),
    .C(_03950_),
    .Y(_03952_));
 sky130_fd_sc_hd__and2b_1 _10833_ (.A_N(_03951_),
    .B(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__xnor2_1 _10834_ (.A(_03949_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21oi_1 _10835_ (.A1(_03835_),
    .A2(_03839_),
    .B1(_03838_),
    .Y(_03955_));
 sky130_fd_sc_hd__or2_1 _10836_ (.A(_03954_),
    .B(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__xnor2_1 _10837_ (.A(_03954_),
    .B(_03955_),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2b_1 _10838_ (.A_N(_03957_),
    .B(_03948_),
    .Y(_03958_));
 sky130_fd_sc_hd__xnor2_1 _10839_ (.A(_03948_),
    .B(_03957_),
    .Y(_03959_));
 sky130_fd_sc_hd__and2_1 _10840_ (.A(_03947_),
    .B(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__or2_1 _10841_ (.A(_03947_),
    .B(_03959_),
    .X(_03961_));
 sky130_fd_sc_hd__xor2_1 _10842_ (.A(_03947_),
    .B(_03959_),
    .X(_03962_));
 sky130_fd_sc_hd__xnor2_1 _10843_ (.A(_03897_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__a21oi_1 _10844_ (.A1(_03773_),
    .A2(_03845_),
    .B1(_03844_),
    .Y(_03964_));
 sky130_fd_sc_hd__or2_1 _10845_ (.A(_03963_),
    .B(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__and2_1 _10846_ (.A(_03963_),
    .B(_03964_),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _10847_ (.A(_03963_),
    .B(_03964_),
    .Y(_03967_));
 sky130_fd_sc_hd__nand2_1 _10848_ (.A(_03965_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__and2b_1 _10849_ (.A_N(_03728_),
    .B(_03849_),
    .X(_03969_));
 sky130_fd_sc_hd__nand2_1 _10850_ (.A(_03729_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2b_1 _10851_ (.A_N(_03970_),
    .B(_03488_),
    .Y(_03971_));
 sky130_fd_sc_hd__a21oi_2 _10852_ (.A1(_03726_),
    .A2(_03847_),
    .B1(_03848_),
    .Y(_03972_));
 sky130_fd_sc_hd__a21oi_1 _10853_ (.A1(_03732_),
    .A2(_03969_),
    .B1(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__o311a_2 _10854_ (.A1(_02945_),
    .A2(_03486_),
    .A3(_03970_),
    .B1(_03971_),
    .C1(_03973_),
    .X(_03974_));
 sky130_fd_sc_hd__xor2_2 _10855_ (.A(_03968_),
    .B(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__a21oi_1 _10856_ (.A1(_03896_),
    .A2(_03975_),
    .B1(_02242_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ai_1 _10857_ (.A1(_03896_),
    .A2(_03975_),
    .B1(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__a21oi_1 _10858_ (.A1(_02185_),
    .A2(_02186_),
    .B1(net150),
    .Y(_03978_));
 sky130_fd_sc_hd__xnor2_1 _10859_ (.A(_02187_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _10860_ (.A(_02317_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__a21oi_1 _10861_ (.A1(_06269_),
    .A2(_03862_),
    .B1(_06263_),
    .Y(_03981_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(_06356_),
    .A1(_03981_),
    .S(net297),
    .X(_03982_));
 sky130_fd_sc_hd__nor2_1 _10863_ (.A(_06221_),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__a211o_1 _10864_ (.A1(_06221_),
    .A2(_03982_),
    .B1(_03983_),
    .C1(net241),
    .X(_03984_));
 sky130_fd_sc_hd__or2_1 _10865_ (.A(net224),
    .B(_02961_),
    .X(_03985_));
 sky130_fd_sc_hd__o211a_1 _10866_ (.A1(net222),
    .A2(_02959_),
    .B1(_03985_),
    .C1(net225),
    .X(_03986_));
 sky130_fd_sc_hd__a21oi_2 _10867_ (.A1(net226),
    .A2(_02820_),
    .B1(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _10868_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .Y(_03988_));
 sky130_fd_sc_hd__or2_1 _10869_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .X(_03989_));
 sky130_fd_sc_hd__o211a_1 _10870_ (.A1(_03866_),
    .A2(_03870_),
    .B1(_03988_),
    .C1(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__a211o_1 _10871_ (.A1(_03988_),
    .A2(_03989_),
    .B1(_03866_),
    .C1(_03870_),
    .X(_03991_));
 sky130_fd_sc_hd__or3b_1 _10872_ (.A(net229),
    .B(_03990_),
    .C_N(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__o21a_1 _10873_ (.A1(net261),
    .A2(_03987_),
    .B1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__or2_1 _10874_ (.A(\div_res[11] ),
    .B(_03876_),
    .X(_03994_));
 sky130_fd_sc_hd__a21oi_1 _10875_ (.A1(net156),
    .A2(_03994_),
    .B1(\div_res[12] ),
    .Y(_03995_));
 sky130_fd_sc_hd__a31o_1 _10876_ (.A1(\div_res[12] ),
    .A2(net156),
    .A3(_03994_),
    .B1(net198),
    .X(_03996_));
 sky130_fd_sc_hd__or2_1 _10877_ (.A(\div_shifter[43] ),
    .B(_03879_),
    .X(_03997_));
 sky130_fd_sc_hd__a21oi_1 _10878_ (.A1(net234),
    .A2(_03997_),
    .B1(\div_shifter[44] ),
    .Y(_03998_));
 sky130_fd_sc_hd__a31o_1 _10879_ (.A1(\div_shifter[44] ),
    .A2(net234),
    .A3(_03997_),
    .B1(net239),
    .X(_03999_));
 sky130_fd_sc_hd__o2bb2a_1 _10880_ (.A1_N(_06194_),
    .A2_N(_06455_),
    .B1(net236),
    .B2(reg1_val[12]),
    .X(_04000_));
 sky130_fd_sc_hd__o221a_1 _10881_ (.A1(_06212_),
    .A2(_02320_),
    .B1(_02323_),
    .B2(_06203_),
    .C1(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__o221a_1 _10882_ (.A1(_06221_),
    .A2(_02327_),
    .B1(_03998_),
    .B2(_03999_),
    .C1(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__o21ai_2 _10883_ (.A1(net226),
    .A2(_02810_),
    .B1(_02338_),
    .Y(_04003_));
 sky130_fd_sc_hd__o221a_1 _10884_ (.A1(_03995_),
    .A2(_03996_),
    .B1(_04003_),
    .B2(_02247_),
    .C1(_04002_),
    .X(_04004_));
 sky130_fd_sc_hd__o221a_1 _10885_ (.A1(_02316_),
    .A2(_03987_),
    .B1(_03993_),
    .B2(net209),
    .C1(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__a41o_1 _10886_ (.A1(_03977_),
    .A2(_03980_),
    .A3(_03984_),
    .A4(_04005_),
    .B1(net259),
    .X(_04006_));
 sky130_fd_sc_hd__and3_2 _10887_ (.A(curr_PC[11]),
    .B(curr_PC[12]),
    .C(_03768_),
    .X(_04007_));
 sky130_fd_sc_hd__o21ai_2 _10888_ (.A1(curr_PC[12]),
    .A2(_03892_),
    .B1(net258),
    .Y(_04008_));
 sky130_fd_sc_hd__o21ai_4 _10889_ (.A1(_04007_),
    .A2(_04008_),
    .B1(_04006_),
    .Y(dest_val[12]));
 sky130_fd_sc_hd__o31a_1 _10890_ (.A1(_03646_),
    .A2(_03894_),
    .A3(_03975_),
    .B1(net151),
    .X(_04009_));
 sky130_fd_sc_hd__o22a_1 _10891_ (.A1(_00349_),
    .A2(net52),
    .B1(net50),
    .B2(net24),
    .X(_04010_));
 sky130_fd_sc_hd__xnor2_1 _10892_ (.A(net88),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_1 _10893_ (.A(net129),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__xor2_1 _10894_ (.A(net129),
    .B(_04011_),
    .X(_04013_));
 sky130_fd_sc_hd__o22a_1 _10895_ (.A1(net54),
    .A2(net18),
    .B1(net9),
    .B2(net95),
    .X(_04014_));
 sky130_fd_sc_hd__xnor2_1 _10896_ (.A(net126),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2b_1 _10897_ (.A_N(_04015_),
    .B(_04013_),
    .Y(_04016_));
 sky130_fd_sc_hd__xor2_1 _10898_ (.A(_04013_),
    .B(_04015_),
    .X(_04017_));
 sky130_fd_sc_hd__o22a_1 _10899_ (.A1(net104),
    .A2(net27),
    .B1(net25),
    .B2(net100),
    .X(_04018_));
 sky130_fd_sc_hd__xnor2_1 _10900_ (.A(net67),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__o22a_1 _10901_ (.A1(net32),
    .A2(net74),
    .B1(net71),
    .B2(net29),
    .X(_04020_));
 sky130_fd_sc_hd__xnor2_1 _10902_ (.A(net117),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__and2b_1 _10903_ (.A_N(_04019_),
    .B(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__xor2_1 _10904_ (.A(_04019_),
    .B(_04021_),
    .X(_04023_));
 sky130_fd_sc_hd__o22a_1 _10905_ (.A1(net35),
    .A2(net108),
    .B1(net70),
    .B2(net37),
    .X(_04024_));
 sky130_fd_sc_hd__xnor2_1 _10906_ (.A(net120),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__and2b_1 _10907_ (.A_N(_04023_),
    .B(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__xor2_1 _10908_ (.A(_04023_),
    .B(_04025_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_1 _10909_ (.A(_04017_),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__xor2_1 _10910_ (.A(_04017_),
    .B(_04027_),
    .X(_04029_));
 sky130_fd_sc_hd__o22a_1 _10911_ (.A1(net33),
    .A2(net78),
    .B1(net63),
    .B2(net79),
    .X(_04030_));
 sky130_fd_sc_hd__xnor2_1 _10912_ (.A(net113),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__o22a_1 _10913_ (.A1(net21),
    .A2(net48),
    .B1(net13),
    .B2(net60),
    .X(_04032_));
 sky130_fd_sc_hd__xnor2_1 _10914_ (.A(net87),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__and2_1 _10915_ (.A(_04031_),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__nor2_1 _10916_ (.A(_04031_),
    .B(_04033_),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_1 _10917_ (.A(_04034_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__o22a_1 _10918_ (.A1(net59),
    .A2(net47),
    .B1(net11),
    .B2(net64),
    .X(_04037_));
 sky130_fd_sc_hd__xnor2_1 _10919_ (.A(net112),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__xor2_1 _10920_ (.A(_04036_),
    .B(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__xnor2_1 _10921_ (.A(_04029_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__o22a_1 _10922_ (.A1(net57),
    .A2(net15),
    .B1(net7),
    .B2(net93),
    .X(_04041_));
 sky130_fd_sc_hd__xnor2_1 _10923_ (.A(net42),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__o21ai_1 _10924_ (.A1(_03939_),
    .A2(_03941_),
    .B1(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__or3_1 _10925_ (.A(_03939_),
    .B(_03941_),
    .C(_04042_),
    .X(_04044_));
 sky130_fd_sc_hd__nand2_1 _10926_ (.A(_04043_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__or2_1 _10927_ (.A(net91),
    .B(net40),
    .X(_04046_));
 sky130_fd_sc_hd__xnor2_1 _10928_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__nor2_1 _10929_ (.A(_04040_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__nand2_1 _10930_ (.A(_04040_),
    .B(_04047_),
    .Y(_04049_));
 sky130_fd_sc_hd__nand2b_1 _10931_ (.A_N(_04048_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__a21o_1 _10932_ (.A1(_03922_),
    .A2(_03924_),
    .B1(_03920_),
    .X(_04051_));
 sky130_fd_sc_hd__a21oi_1 _10933_ (.A1(_03908_),
    .A2(_03912_),
    .B1(_03902_),
    .Y(_04052_));
 sky130_fd_sc_hd__and3_1 _10934_ (.A(_03902_),
    .B(_03908_),
    .C(_03912_),
    .X(_04053_));
 sky130_fd_sc_hd__or2_1 _10935_ (.A(_04052_),
    .B(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__and2b_1 _10936_ (.A_N(_04054_),
    .B(_04051_),
    .X(_04055_));
 sky130_fd_sc_hd__xnor2_1 _10937_ (.A(_04051_),
    .B(_04054_),
    .Y(_04056_));
 sky130_fd_sc_hd__xnor2_1 _10938_ (.A(_04050_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__o21ai_1 _10939_ (.A1(_03936_),
    .A2(_03946_),
    .B1(_03934_),
    .Y(_04058_));
 sky130_fd_sc_hd__a21bo_1 _10940_ (.A1(_03937_),
    .A2(_03944_),
    .B1_N(_03943_),
    .X(_04059_));
 sky130_fd_sc_hd__a21oi_1 _10941_ (.A1(_03928_),
    .A2(_03932_),
    .B1(_03931_),
    .Y(_04060_));
 sky130_fd_sc_hd__o21ba_1 _10942_ (.A1(_03914_),
    .A2(_03926_),
    .B1_N(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__or3b_1 _10943_ (.A(_03914_),
    .B(_03926_),
    .C_N(_04060_),
    .X(_04062_));
 sky130_fd_sc_hd__and2b_1 _10944_ (.A_N(_04061_),
    .B(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__xnor2_1 _10945_ (.A(_04059_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__a21oi_1 _10946_ (.A1(_03949_),
    .A2(_03952_),
    .B1(_03951_),
    .Y(_04065_));
 sky130_fd_sc_hd__xnor2_1 _10947_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2b_1 _10948_ (.A_N(_04066_),
    .B(_04058_),
    .Y(_04067_));
 sky130_fd_sc_hd__xnor2_1 _10949_ (.A(_04058_),
    .B(_04066_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand2_1 _10950_ (.A(_04057_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__xnor2_1 _10951_ (.A(_04057_),
    .B(_04068_),
    .Y(_04070_));
 sky130_fd_sc_hd__a21o_1 _10952_ (.A1(_03956_),
    .A2(_03958_),
    .B1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__nand3_1 _10953_ (.A(_03956_),
    .B(_03958_),
    .C(_04070_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _10954_ (.A(_04071_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__a21oi_2 _10955_ (.A1(_03897_),
    .A2(_03961_),
    .B1(_03960_),
    .Y(_04074_));
 sky130_fd_sc_hd__or2_1 _10956_ (.A(_04073_),
    .B(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__and2_1 _10957_ (.A(_04073_),
    .B(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__xnor2_2 _10958_ (.A(_04073_),
    .B(_04074_),
    .Y(_04077_));
 sky130_fd_sc_hd__and3_1 _10959_ (.A(_03849_),
    .B(_03965_),
    .C(_03967_),
    .X(_04078_));
 sky130_fd_sc_hd__nand2_1 _10960_ (.A(_03851_),
    .B(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2b_1 _10961_ (.A_N(_04079_),
    .B(_03612_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21oi_1 _10962_ (.A1(_03847_),
    .A2(_03965_),
    .B1(_03966_),
    .Y(_04081_));
 sky130_fd_sc_hd__a21oi_1 _10963_ (.A1(_03850_),
    .A2(_04078_),
    .B1(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__o311a_2 _10964_ (.A1(_03088_),
    .A2(_03610_),
    .A3(_04079_),
    .B1(_04080_),
    .C1(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__xor2_2 _10965_ (.A(_04077_),
    .B(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__o21ai_1 _10966_ (.A1(_04009_),
    .A2(_04084_),
    .B1(net202),
    .Y(_04085_));
 sky130_fd_sc_hd__a21o_1 _10967_ (.A1(_04009_),
    .A2(_04084_),
    .B1(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__o21a_1 _10968_ (.A1(net150),
    .A2(_02188_),
    .B1(_02189_),
    .X(_04087_));
 sky130_fd_sc_hd__o31ai_1 _10969_ (.A1(net150),
    .A2(_02188_),
    .A3(_02189_),
    .B1(_02317_),
    .Y(_04088_));
 sky130_fd_sc_hd__o21a_1 _10970_ (.A1(_06221_),
    .A2(_03981_),
    .B1(_06212_),
    .X(_04089_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(_06358_),
    .A1(_04089_),
    .S(net297),
    .X(_04090_));
 sky130_fd_sc_hd__nor2_1 _10972_ (.A(_06176_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a211o_1 _10973_ (.A1(_06176_),
    .A2(_04090_),
    .B1(_04091_),
    .C1(net241),
    .X(_04092_));
 sky130_fd_sc_hd__nand2_1 _10974_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .Y(_04093_));
 sky130_fd_sc_hd__or2_1 _10975_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .X(_04094_));
 sky130_fd_sc_hd__nand2_1 _10976_ (.A(_04093_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__a21oi_1 _10977_ (.A1(reg1_val[12]),
    .A2(curr_PC[12]),
    .B1(_03990_),
    .Y(_04096_));
 sky130_fd_sc_hd__xnor2_1 _10978_ (.A(_04095_),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__or2_1 _10979_ (.A(net224),
    .B(_03103_),
    .X(_04098_));
 sky130_fd_sc_hd__o211a_1 _10980_ (.A1(net223),
    .A2(_03101_),
    .B1(_04098_),
    .C1(net225),
    .X(_04099_));
 sky130_fd_sc_hd__a21oi_2 _10981_ (.A1(net227),
    .A2(_02648_),
    .B1(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(_04097_),
    .A1(_04100_),
    .S(net229),
    .X(_04101_));
 sky130_fd_sc_hd__or2_1 _10983_ (.A(\div_res[12] ),
    .B(_03994_),
    .X(_04102_));
 sky130_fd_sc_hd__a21oi_1 _10984_ (.A1(net154),
    .A2(_04102_),
    .B1(\div_res[13] ),
    .Y(_04103_));
 sky130_fd_sc_hd__a31o_1 _10985_ (.A1(\div_res[13] ),
    .A2(net154),
    .A3(_04102_),
    .B1(net198),
    .X(_04104_));
 sky130_fd_sc_hd__or2_1 _10986_ (.A(\div_shifter[44] ),
    .B(_03997_),
    .X(_04105_));
 sky130_fd_sc_hd__a21oi_1 _10987_ (.A1(net234),
    .A2(_04105_),
    .B1(\div_shifter[45] ),
    .Y(_04106_));
 sky130_fd_sc_hd__a31o_1 _10988_ (.A1(\div_shifter[45] ),
    .A2(net234),
    .A3(_04105_),
    .B1(net239),
    .X(_04107_));
 sky130_fd_sc_hd__o2bb2a_1 _10989_ (.A1_N(_06149_),
    .A2_N(_06455_),
    .B1(net236),
    .B2(reg1_val[13]),
    .X(_04108_));
 sky130_fd_sc_hd__o221a_1 _10990_ (.A1(_06167_),
    .A2(_02320_),
    .B1(_02323_),
    .B2(_06158_),
    .C1(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__o221a_1 _10991_ (.A1(_06176_),
    .A2(_02327_),
    .B1(_04106_),
    .B2(_04107_),
    .C1(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__o21ai_2 _10992_ (.A1(net227),
    .A2(_02662_),
    .B1(_02338_),
    .Y(_04111_));
 sky130_fd_sc_hd__o221a_1 _10993_ (.A1(_04103_),
    .A2(_04104_),
    .B1(_04111_),
    .B2(_02247_),
    .C1(_04110_),
    .X(_04112_));
 sky130_fd_sc_hd__o221a_1 _10994_ (.A1(_02316_),
    .A2(_04100_),
    .B1(_04101_),
    .B2(net209),
    .C1(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__o211a_1 _10995_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04092_),
    .C1(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__a21oi_1 _10996_ (.A1(_04086_),
    .A2(_04114_),
    .B1(net259),
    .Y(_04115_));
 sky130_fd_sc_hd__or2_1 _10997_ (.A(curr_PC[13]),
    .B(_04007_),
    .X(_04116_));
 sky130_fd_sc_hd__nand2_1 _10998_ (.A(curr_PC[13]),
    .B(_04007_),
    .Y(_04117_));
 sky130_fd_sc_hd__a31o_4 _10999_ (.A1(net258),
    .A2(_04116_),
    .A3(_04117_),
    .B1(_04115_),
    .X(dest_val[13]));
 sky130_fd_sc_hd__or4_1 _11000_ (.A(_03646_),
    .B(_03894_),
    .C(_03975_),
    .D(_04084_),
    .X(_04118_));
 sky130_fd_sc_hd__o21ai_1 _11001_ (.A1(_04064_),
    .A2(_04065_),
    .B1(_04067_),
    .Y(_04119_));
 sky130_fd_sc_hd__a21o_1 _11002_ (.A1(_04036_),
    .A2(_04038_),
    .B1(_04034_),
    .X(_04120_));
 sky130_fd_sc_hd__nor2_1 _11003_ (.A(_04022_),
    .B(_04026_),
    .Y(_04121_));
 sky130_fd_sc_hd__a21oi_1 _11004_ (.A1(_04012_),
    .A2(_04016_),
    .B1(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__and3_1 _11005_ (.A(_04012_),
    .B(_04016_),
    .C(_04121_),
    .X(_04123_));
 sky130_fd_sc_hd__nor2_1 _11006_ (.A(_04122_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_2 _11007_ (.A(_04120_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__o22a_1 _11008_ (.A1(net100),
    .A2(net15),
    .B1(net7),
    .B2(net57),
    .X(_04126_));
 sky130_fd_sc_hd__xnor2_1 _11009_ (.A(net40),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__o22a_1 _11010_ (.A1(net108),
    .A2(net27),
    .B1(net26),
    .B2(net104),
    .X(_04128_));
 sky130_fd_sc_hd__xnor2_1 _11011_ (.A(net66),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_2 _11012_ (.A(_00323_),
    .B(net45),
    .Y(_04130_));
 sky130_fd_sc_hd__nor2_1 _11013_ (.A(_04129_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__and2_1 _11014_ (.A(_04129_),
    .B(_04130_),
    .X(_04132_));
 sky130_fd_sc_hd__or2_1 _11015_ (.A(_04131_),
    .B(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__nor2_1 _11016_ (.A(_04127_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _11017_ (.A(_04127_),
    .B(_04133_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand2b_1 _11018_ (.A_N(_04134_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__o22a_1 _11019_ (.A1(net23),
    .A2(net48),
    .B1(net13),
    .B2(net21),
    .X(_04137_));
 sky130_fd_sc_hd__xnor2_1 _11020_ (.A(net87),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__o22a_1 _11021_ (.A1(net79),
    .A2(net64),
    .B1(net63),
    .B2(net33),
    .X(_04139_));
 sky130_fd_sc_hd__xnor2_1 _11022_ (.A(net113),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__and2_1 _11023_ (.A(_04138_),
    .B(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__nor2_1 _11024_ (.A(_04138_),
    .B(_04140_),
    .Y(_04142_));
 sky130_fd_sc_hd__nor2_1 _11025_ (.A(_04141_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__o22a_1 _11026_ (.A1(net60),
    .A2(net47),
    .B1(net11),
    .B2(net59),
    .X(_04144_));
 sky130_fd_sc_hd__xnor2_2 _11027_ (.A(net112),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__xor2_2 _11028_ (.A(_04143_),
    .B(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__o22a_1 _11029_ (.A1(net32),
    .A2(net78),
    .B1(net74),
    .B2(net29),
    .X(_04147_));
 sky130_fd_sc_hd__xnor2_1 _11030_ (.A(net116),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__o22a_1 _11031_ (.A1(net37),
    .A2(net71),
    .B1(net70),
    .B2(net35),
    .X(_04149_));
 sky130_fd_sc_hd__xnor2_1 _11032_ (.A(net120),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__and2_1 _11033_ (.A(_04148_),
    .B(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__nor2_1 _11034_ (.A(_04148_),
    .B(_04150_),
    .Y(_04152_));
 sky130_fd_sc_hd__nor2_1 _11035_ (.A(_04151_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__o22a_1 _11036_ (.A1(net17),
    .A2(net52),
    .B1(net50),
    .B2(_00349_),
    .X(_04154_));
 sky130_fd_sc_hd__xnor2_1 _11037_ (.A(net88),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__a31o_1 _11038_ (.A1(net130),
    .A2(_00321_),
    .A3(_00567_),
    .B1(net127),
    .X(_04156_));
 sky130_fd_sc_hd__o21ai_4 _11039_ (.A1(_00326_),
    .A2(net9),
    .B1(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__nor2_1 _11040_ (.A(_04155_),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__and2_1 _11041_ (.A(_04155_),
    .B(_04157_),
    .X(_04159_));
 sky130_fd_sc_hd__nor2_1 _11042_ (.A(_04158_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__and2b_1 _11043_ (.A_N(_04160_),
    .B(_04153_),
    .X(_04161_));
 sky130_fd_sc_hd__xnor2_2 _11044_ (.A(_04153_),
    .B(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__xnor2_2 _11045_ (.A(_04146_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__xor2_2 _11046_ (.A(_04136_),
    .B(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__and2b_1 _11047_ (.A_N(_04125_),
    .B(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__xnor2_2 _11048_ (.A(_04125_),
    .B(_04164_),
    .Y(_04166_));
 sky130_fd_sc_hd__a21oi_1 _11049_ (.A1(_04049_),
    .A2(_04056_),
    .B1(_04048_),
    .Y(_04167_));
 sky130_fd_sc_hd__a21o_1 _11050_ (.A1(_04029_),
    .A2(_04039_),
    .B1(_04028_),
    .X(_04168_));
 sky130_fd_sc_hd__o21ai_1 _11051_ (.A1(_04045_),
    .A2(_04046_),
    .B1(_04043_),
    .Y(_04169_));
 sky130_fd_sc_hd__xor2_1 _11052_ (.A(_04168_),
    .B(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__o21ai_1 _11053_ (.A1(_04052_),
    .A2(_04055_),
    .B1(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__or3_1 _11054_ (.A(_04052_),
    .B(_04055_),
    .C(_04170_),
    .X(_04172_));
 sky130_fd_sc_hd__nand2_1 _11055_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__a21o_1 _11056_ (.A1(_04059_),
    .A2(_04063_),
    .B1(_04061_),
    .X(_04174_));
 sky130_fd_sc_hd__nand2b_1 _11057_ (.A_N(_04173_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__xnor2_1 _11058_ (.A(_04173_),
    .B(_04174_),
    .Y(_04176_));
 sky130_fd_sc_hd__nand2b_1 _11059_ (.A_N(_04167_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__xnor2_1 _11060_ (.A(_04167_),
    .B(_04176_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand2_1 _11061_ (.A(_04166_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__xnor2_1 _11062_ (.A(_04166_),
    .B(_04178_),
    .Y(_04180_));
 sky130_fd_sc_hd__nand2b_1 _11063_ (.A_N(_04180_),
    .B(_04119_),
    .Y(_04181_));
 sky130_fd_sc_hd__xor2_1 _11064_ (.A(_04119_),
    .B(_04180_),
    .X(_04182_));
 sky130_fd_sc_hd__a21oi_2 _11065_ (.A1(_04069_),
    .A2(_04071_),
    .B1(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__inv_2 _11066_ (.A(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__and3_1 _11067_ (.A(_04069_),
    .B(_04071_),
    .C(_04182_),
    .X(_04185_));
 sky130_fd_sc_hd__or2_2 _11068_ (.A(_04183_),
    .B(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__a21oi_1 _11069_ (.A1(_03965_),
    .A2(_04075_),
    .B1(_04076_),
    .Y(_04187_));
 sky130_fd_sc_hd__nor2_1 _11070_ (.A(_03968_),
    .B(_04077_),
    .Y(_04188_));
 sky130_fd_sc_hd__a21o_1 _11071_ (.A1(_03972_),
    .A2(_04188_),
    .B1(_04187_),
    .X(_04189_));
 sky130_fd_sc_hd__a31o_1 _11072_ (.A1(_03734_),
    .A2(_03969_),
    .A3(_04188_),
    .B1(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__xnor2_2 _11073_ (.A(_04186_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__a21oi_1 _11074_ (.A1(net151),
    .A2(_04118_),
    .B1(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__a31o_1 _11075_ (.A1(net151),
    .A2(_04118_),
    .A3(_04191_),
    .B1(_02242_),
    .X(_04193_));
 sky130_fd_sc_hd__or2_4 _11076_ (.A(_04192_),
    .B(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__a21o_1 _11077_ (.A1(_02188_),
    .A2(_02189_),
    .B1(net150),
    .X(_04195_));
 sky130_fd_sc_hd__a21oi_1 _11078_ (.A1(_02190_),
    .A2(_04195_),
    .B1(_02318_),
    .Y(_04196_));
 sky130_fd_sc_hd__o21ai_1 _11079_ (.A1(_02190_),
    .A2(_04195_),
    .B1(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__o21ai_1 _11080_ (.A1(_06176_),
    .A2(_04089_),
    .B1(_06167_),
    .Y(_04198_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(_06360_),
    .A1(_04198_),
    .S(net297),
    .X(_04199_));
 sky130_fd_sc_hd__o21ai_1 _11082_ (.A1(_06125_),
    .A2(_04199_),
    .B1(net242),
    .Y(_04200_));
 sky130_fd_sc_hd__a21o_1 _11083_ (.A1(_06125_),
    .A2(_04199_),
    .B1(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__nand2_1 _11084_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .Y(_04202_));
 sky130_fd_sc_hd__or2_1 _11085_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .X(_04203_));
 sky130_fd_sc_hd__nand2_1 _11086_ (.A(_04202_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21a_1 _11087_ (.A1(_04095_),
    .A2(_04096_),
    .B1(_04093_),
    .X(_04205_));
 sky130_fd_sc_hd__xnor2_1 _11088_ (.A(_04204_),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__or2_1 _11089_ (.A(net224),
    .B(_03241_),
    .X(_04207_));
 sky130_fd_sc_hd__o211a_1 _11090_ (.A1(net222),
    .A2(_03240_),
    .B1(_04207_),
    .C1(net225),
    .X(_04208_));
 sky130_fd_sc_hd__a21oi_2 _11091_ (.A1(net226),
    .A2(_02526_),
    .B1(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__inv_2 _11092_ (.A(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(_04206_),
    .A1(_04209_),
    .S(net229),
    .X(_04211_));
 sky130_fd_sc_hd__o21ai_1 _11094_ (.A1(\div_res[13] ),
    .A2(_04102_),
    .B1(net156),
    .Y(_04212_));
 sky130_fd_sc_hd__xnor2_1 _11095_ (.A(\div_res[14] ),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__o21a_1 _11096_ (.A1(\div_shifter[45] ),
    .A2(_04105_),
    .B1(net234),
    .X(_04214_));
 sky130_fd_sc_hd__o21ai_1 _11097_ (.A1(\div_shifter[46] ),
    .A2(_04214_),
    .B1(_02332_),
    .Y(_04215_));
 sky130_fd_sc_hd__a21oi_1 _11098_ (.A1(\div_shifter[46] ),
    .A2(_04214_),
    .B1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__nor2_1 _11099_ (.A(reg1_val[14]),
    .B(net236),
    .Y(_04217_));
 sky130_fd_sc_hd__a221o_1 _11100_ (.A1(_06101_),
    .A2(_06455_),
    .B1(net273),
    .B2(_06113_),
    .C1(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__a221o_1 _11101_ (.A1(_06119_),
    .A2(net201),
    .B1(net240),
    .B2(_06125_),
    .C1(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__a211o_1 _11102_ (.A1(_02330_),
    .A2(_04213_),
    .B1(_04216_),
    .C1(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__o21a_1 _11103_ (.A1(net227),
    .A2(_02500_),
    .B1(_02338_),
    .X(_04221_));
 sky130_fd_sc_hd__a21oi_1 _11104_ (.A1(net246),
    .A2(_04221_),
    .B1(_04220_),
    .Y(_04222_));
 sky130_fd_sc_hd__o221a_1 _11105_ (.A1(_02316_),
    .A2(_04209_),
    .B1(_04211_),
    .B2(net209),
    .C1(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__a41o_2 _11106_ (.A1(_04194_),
    .A2(_04197_),
    .A3(_04201_),
    .A4(_04223_),
    .B1(_06427_),
    .X(_04224_));
 sky130_fd_sc_hd__and3_1 _11107_ (.A(curr_PC[13]),
    .B(curr_PC[14]),
    .C(_04007_),
    .X(_04225_));
 sky130_fd_sc_hd__a21oi_1 _11108_ (.A1(curr_PC[13]),
    .A2(_04007_),
    .B1(curr_PC[14]),
    .Y(_04226_));
 sky130_fd_sc_hd__o31ai_4 _11109_ (.A1(net253),
    .A2(_04225_),
    .A3(_04226_),
    .B1(_04224_),
    .Y(dest_val[14]));
 sky130_fd_sc_hd__o21a_1 _11110_ (.A1(_04118_),
    .A2(_04191_),
    .B1(net151),
    .X(_04227_));
 sky130_fd_sc_hd__o22a_1 _11111_ (.A1(net29),
    .A2(net78),
    .B1(net63),
    .B2(net32),
    .X(_04228_));
 sky130_fd_sc_hd__xnor2_1 _11112_ (.A(net116),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__o22a_1 _11113_ (.A1(net21),
    .A2(net47),
    .B1(net11),
    .B2(net60),
    .X(_04230_));
 sky130_fd_sc_hd__xnor2_1 _11114_ (.A(net112),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__and2_1 _11115_ (.A(_04229_),
    .B(_04231_),
    .X(_04232_));
 sky130_fd_sc_hd__xor2_1 _11116_ (.A(_04229_),
    .B(_04231_),
    .X(_04233_));
 sky130_fd_sc_hd__o22a_1 _11117_ (.A1(net33),
    .A2(net64),
    .B1(net59),
    .B2(net79),
    .X(_04234_));
 sky130_fd_sc_hd__xnor2_1 _11118_ (.A(net113),
    .B(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__xor2_1 _11119_ (.A(_04233_),
    .B(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__and2_1 _11120_ (.A(_04151_),
    .B(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__xnor2_1 _11121_ (.A(_04151_),
    .B(_04236_),
    .Y(_04238_));
 sky130_fd_sc_hd__o22a_1 _11122_ (.A1(net19),
    .A2(net48),
    .B1(net13),
    .B2(net23),
    .X(_04239_));
 sky130_fd_sc_hd__xnor2_1 _11123_ (.A(net87),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__and2_1 _11124_ (.A(net126),
    .B(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__nor2_1 _11125_ (.A(net126),
    .B(_04240_),
    .Y(_04242_));
 sky130_fd_sc_hd__nor2_1 _11126_ (.A(_04241_),
    .B(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__o22a_1 _11127_ (.A1(net17),
    .A2(net50),
    .B1(net8),
    .B2(net52),
    .X(_04244_));
 sky130_fd_sc_hd__xnor2_1 _11128_ (.A(net88),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__xnor2_1 _11129_ (.A(_04243_),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__nor2_1 _11130_ (.A(_04238_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__and2_1 _11131_ (.A(_04238_),
    .B(_04246_),
    .X(_04248_));
 sky130_fd_sc_hd__o22a_1 _11132_ (.A1(net70),
    .A2(net27),
    .B1(net26),
    .B2(net108),
    .X(_04249_));
 sky130_fd_sc_hd__xnor2_1 _11133_ (.A(net67),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__o22a_1 _11134_ (.A1(net104),
    .A2(net15),
    .B1(net6),
    .B2(net100),
    .X(_04251_));
 sky130_fd_sc_hd__xnor2_1 _11135_ (.A(net42),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o22a_1 _11136_ (.A1(net37),
    .A2(net74),
    .B1(net71),
    .B2(net35),
    .X(_04253_));
 sky130_fd_sc_hd__xnor2_1 _11137_ (.A(net120),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__and2_1 _11138_ (.A(_04252_),
    .B(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__nor2_1 _11139_ (.A(_04252_),
    .B(_04254_),
    .Y(_04256_));
 sky130_fd_sc_hd__nor2_1 _11140_ (.A(_04255_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__and2b_1 _11141_ (.A_N(_04250_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__xor2_1 _11142_ (.A(_04250_),
    .B(_04257_),
    .X(_04259_));
 sky130_fd_sc_hd__nor3_1 _11143_ (.A(_04247_),
    .B(_04248_),
    .C(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__o21ai_1 _11144_ (.A1(_04247_),
    .A2(_04248_),
    .B1(_04259_),
    .Y(_04261_));
 sky130_fd_sc_hd__nand2b_1 _11145_ (.A_N(_04260_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21oi_1 _11146_ (.A1(_04143_),
    .A2(_04145_),
    .B1(_04141_),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_2 _11147_ (.A(_00310_),
    .B(net45),
    .Y(_04264_));
 sky130_fd_sc_hd__xnor2_1 _11148_ (.A(_04263_),
    .B(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__nor2_1 _11149_ (.A(_04158_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__and2_1 _11150_ (.A(_04158_),
    .B(_04265_),
    .X(_04267_));
 sky130_fd_sc_hd__nor2_1 _11151_ (.A(_04266_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__xnor2_1 _11152_ (.A(_04262_),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__o21ba_1 _11153_ (.A1(_04136_),
    .A2(_04163_),
    .B1_N(_04165_),
    .X(_04270_));
 sky130_fd_sc_hd__a21bo_1 _11154_ (.A1(_04168_),
    .A2(_04169_),
    .B1_N(_04171_),
    .X(_04271_));
 sky130_fd_sc_hd__a21o_1 _11155_ (.A1(_04120_),
    .A2(_04124_),
    .B1(_04122_),
    .X(_04272_));
 sky130_fd_sc_hd__a21oi_1 _11156_ (.A1(_04146_),
    .A2(_04162_),
    .B1(_04161_),
    .Y(_04273_));
 sky130_fd_sc_hd__o21bai_1 _11157_ (.A1(_04131_),
    .A2(_04134_),
    .B1_N(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__or3b_1 _11158_ (.A(_04131_),
    .B(_04134_),
    .C_N(_04273_),
    .X(_04275_));
 sky130_fd_sc_hd__and2_1 _11159_ (.A(_04274_),
    .B(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__xnor2_1 _11160_ (.A(_04272_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2b_1 _11161_ (.A_N(_04277_),
    .B(_04271_),
    .Y(_04278_));
 sky130_fd_sc_hd__xnor2_1 _11162_ (.A(_04271_),
    .B(_04277_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2b_1 _11163_ (.A_N(_04270_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__xnor2_1 _11164_ (.A(_04270_),
    .B(_04279_),
    .Y(_04281_));
 sky130_fd_sc_hd__and2_1 _11165_ (.A(_04269_),
    .B(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__xnor2_1 _11166_ (.A(_04269_),
    .B(_04281_),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_1 _11167_ (.A(_04175_),
    .B(_04177_),
    .Y(_04284_));
 sky130_fd_sc_hd__and2b_1 _11168_ (.A_N(_04283_),
    .B(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__xor2_1 _11169_ (.A(_04283_),
    .B(_04284_),
    .X(_04286_));
 sky130_fd_sc_hd__a21oi_1 _11170_ (.A1(_04179_),
    .A2(_04181_),
    .B1(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__nand3_1 _11171_ (.A(_04179_),
    .B(_04181_),
    .C(_04286_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2b_1 _11172_ (.A_N(_04287_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_1 _11173_ (.A(_04077_),
    .B(_04186_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _11174_ (.A(_04078_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__a21oi_1 _11175_ (.A1(_04075_),
    .A2(_04184_),
    .B1(_04185_),
    .Y(_04292_));
 sky130_fd_sc_hd__a21oi_1 _11176_ (.A1(_04081_),
    .A2(_04290_),
    .B1(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__o21a_1 _11177_ (.A1(_03852_),
    .A2(_04291_),
    .B1(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__o21ai_4 _11178_ (.A1(_03854_),
    .A2(_04291_),
    .B1(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__xnor2_1 _11179_ (.A(_04289_),
    .B(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_1 _11180_ (.A1(_04227_),
    .A2(_04296_),
    .B1(net202),
    .Y(_04297_));
 sky130_fd_sc_hd__a21o_1 _11181_ (.A1(_04227_),
    .A2(_04296_),
    .B1(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__o21a_1 _11182_ (.A1(_02135_),
    .A2(_02191_),
    .B1(_02192_),
    .X(_04299_));
 sky130_fd_sc_hd__or3_1 _11183_ (.A(_02135_),
    .B(_02191_),
    .C(_02192_),
    .X(_04300_));
 sky130_fd_sc_hd__or3b_1 _11184_ (.A(_02318_),
    .B(_04299_),
    .C_N(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__a21oi_1 _11185_ (.A1(_06125_),
    .A2(_04198_),
    .B1(_06119_),
    .Y(_04302_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(_06362_),
    .A1(_04302_),
    .S(net297),
    .X(_04303_));
 sky130_fd_sc_hd__nor2_1 _11187_ (.A(_06089_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__a211o_1 _11188_ (.A1(_06089_),
    .A2(_04303_),
    .B1(_04304_),
    .C1(net241),
    .X(_04305_));
 sky130_fd_sc_hd__nand2_1 _11189_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .Y(_04306_));
 sky130_fd_sc_hd__or2_1 _11190_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .X(_04307_));
 sky130_fd_sc_hd__nand2_1 _11191_ (.A(_04306_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__o21a_1 _11192_ (.A1(_04204_),
    .A2(_04205_),
    .B1(_04202_),
    .X(_04309_));
 sky130_fd_sc_hd__xnor2_1 _11193_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(_03372_),
    .A1(_03374_),
    .S(net223),
    .X(_04311_));
 sky130_fd_sc_hd__and3_1 _11195_ (.A(net227),
    .B(_02343_),
    .C(_02345_),
    .X(_04312_));
 sky130_fd_sc_hd__a21oi_2 _11196_ (.A1(net225),
    .A2(_04311_),
    .B1(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(_04310_),
    .A1(_04313_),
    .S(net229),
    .X(_04314_));
 sky130_fd_sc_hd__or3_1 _11198_ (.A(\div_shifter[46] ),
    .B(\div_shifter[45] ),
    .C(_04105_),
    .X(_04315_));
 sky130_fd_sc_hd__and3_1 _11199_ (.A(\div_shifter[47] ),
    .B(net233),
    .C(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__a21oi_1 _11200_ (.A1(net233),
    .A2(_04315_),
    .B1(\div_shifter[47] ),
    .Y(_04317_));
 sky130_fd_sc_hd__or3_1 _11201_ (.A(\div_res[14] ),
    .B(\div_res[13] ),
    .C(_04102_),
    .X(_04318_));
 sky130_fd_sc_hd__a21oi_1 _11202_ (.A1(net155),
    .A2(_04318_),
    .B1(\div_res[15] ),
    .Y(_04319_));
 sky130_fd_sc_hd__a31o_1 _11203_ (.A1(\div_res[15] ),
    .A2(net155),
    .A3(_04318_),
    .B1(net199),
    .X(_04320_));
 sky130_fd_sc_hd__o2bb2a_1 _11204_ (.A1_N(_06071_),
    .A2_N(_06455_),
    .B1(net236),
    .B2(reg1_val[15]),
    .X(_04321_));
 sky130_fd_sc_hd__o221a_1 _11205_ (.A1(_06083_),
    .A2(_02320_),
    .B1(_02323_),
    .B2(_06077_),
    .C1(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__o221a_1 _11206_ (.A1(_06089_),
    .A2(_02327_),
    .B1(_04319_),
    .B2(_04320_),
    .C1(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__o31a_1 _11207_ (.A1(net238),
    .A2(_04316_),
    .A3(_04317_),
    .B1(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__o21a_1 _11208_ (.A1(net226),
    .A2(_02309_),
    .B1(_02338_),
    .X(_04325_));
 sky130_fd_sc_hd__o2bb2a_1 _11209_ (.A1_N(net246),
    .A2_N(_04325_),
    .B1(_04313_),
    .B2(_02316_),
    .X(_04326_));
 sky130_fd_sc_hd__o211a_1 _11210_ (.A1(net209),
    .A2(_04314_),
    .B1(_04324_),
    .C1(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__a41o_2 _11211_ (.A1(_04298_),
    .A2(_04301_),
    .A3(_04305_),
    .A4(_04327_),
    .B1(_06427_),
    .X(_04328_));
 sky130_fd_sc_hd__nor2_1 _11212_ (.A(curr_PC[15]),
    .B(_04225_),
    .Y(_04329_));
 sky130_fd_sc_hd__and2_2 _11213_ (.A(curr_PC[15]),
    .B(_04225_),
    .X(_04330_));
 sky130_fd_sc_hd__o31ai_4 _11214_ (.A1(net254),
    .A2(_04329_),
    .A3(_04330_),
    .B1(_04328_),
    .Y(dest_val[15]));
 sky130_fd_sc_hd__or4_1 _11215_ (.A(_03975_),
    .B(_04084_),
    .C(_04191_),
    .D(_04296_),
    .X(_04331_));
 sky130_fd_sc_hd__o31a_1 _11216_ (.A1(_03646_),
    .A2(_03894_),
    .A3(_04331_),
    .B1(net151),
    .X(_04332_));
 sky130_fd_sc_hd__nand2_1 _11217_ (.A(_04278_),
    .B(_04280_),
    .Y(_04333_));
 sky130_fd_sc_hd__a21o_1 _11218_ (.A1(_04243_),
    .A2(_04245_),
    .B1(_04241_),
    .X(_04334_));
 sky130_fd_sc_hd__o22a_1 _11219_ (.A1(net108),
    .A2(net15),
    .B1(net6),
    .B2(net104),
    .X(_04335_));
 sky130_fd_sc_hd__xnor2_1 _11220_ (.A(net41),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__xor2_1 _11221_ (.A(_04334_),
    .B(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__and3_1 _11222_ (.A(net99),
    .B(net41),
    .C(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__a21oi_1 _11223_ (.A1(net99),
    .A2(net41),
    .B1(_04337_),
    .Y(_04339_));
 sky130_fd_sc_hd__nor2_1 _11224_ (.A(_04338_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__o22a_1 _11225_ (.A1(net71),
    .A2(net27),
    .B1(net25),
    .B2(net70),
    .X(_04341_));
 sky130_fd_sc_hd__xnor2_1 _11226_ (.A(net66),
    .B(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__o22a_1 _11227_ (.A1(net32),
    .A2(net64),
    .B1(net63),
    .B2(net29),
    .X(_04343_));
 sky130_fd_sc_hd__xnor2_1 _11228_ (.A(net116),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__and2b_1 _11229_ (.A_N(_04342_),
    .B(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__and2b_1 _11230_ (.A_N(_04344_),
    .B(_04342_),
    .X(_04346_));
 sky130_fd_sc_hd__or2_1 _11231_ (.A(_04345_),
    .B(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__o22a_1 _11232_ (.A1(net37),
    .A2(net78),
    .B1(net74),
    .B2(net35),
    .X(_04348_));
 sky130_fd_sc_hd__xnor2_1 _11233_ (.A(net120),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__and2b_1 _11234_ (.A_N(_04347_),
    .B(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__and2b_1 _11235_ (.A_N(_04349_),
    .B(_04347_),
    .X(_04351_));
 sky130_fd_sc_hd__or2_1 _11236_ (.A(_04350_),
    .B(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__o22a_1 _11237_ (.A1(net79),
    .A2(net60),
    .B1(net59),
    .B2(net33),
    .X(_04353_));
 sky130_fd_sc_hd__xnor2_1 _11238_ (.A(net113),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__o22a_1 _11239_ (.A1(net23),
    .A2(net47),
    .B1(net11),
    .B2(net21),
    .X(_04355_));
 sky130_fd_sc_hd__xnor2_2 _11240_ (.A(net112),
    .B(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__xor2_1 _11241_ (.A(_04354_),
    .B(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__a21oi_1 _11242_ (.A1(_04233_),
    .A2(_04235_),
    .B1(_04232_),
    .Y(_04358_));
 sky130_fd_sc_hd__and2b_1 _11243_ (.A_N(_04358_),
    .B(_04357_),
    .X(_04359_));
 sky130_fd_sc_hd__xnor2_1 _11244_ (.A(_04357_),
    .B(_04358_),
    .Y(_04360_));
 sky130_fd_sc_hd__o22a_1 _11245_ (.A1(net17),
    .A2(net48),
    .B1(net13),
    .B2(net19),
    .X(_04361_));
 sky130_fd_sc_hd__xnor2_1 _11246_ (.A(net87),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__o21a_1 _11247_ (.A1(_00391_),
    .A2(net8),
    .B1(net88),
    .X(_04363_));
 sky130_fd_sc_hd__a21o_1 _11248_ (.A1(_00393_),
    .A2(net10),
    .B1(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__nor2_1 _11249_ (.A(_04362_),
    .B(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__and2_1 _11250_ (.A(_04362_),
    .B(_04364_),
    .X(_04366_));
 sky130_fd_sc_hd__nor2_1 _11251_ (.A(_04365_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__and2b_1 _11252_ (.A_N(_04367_),
    .B(_04360_),
    .X(_04368_));
 sky130_fd_sc_hd__and2b_1 _11253_ (.A_N(_04360_),
    .B(_04367_),
    .X(_04369_));
 sky130_fd_sc_hd__nor2_1 _11254_ (.A(_04368_),
    .B(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2b_1 _11255_ (.A_N(_04352_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__xnor2_2 _11256_ (.A(_04352_),
    .B(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__xor2_2 _11257_ (.A(_04340_),
    .B(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__a21oi_1 _11258_ (.A1(_04261_),
    .A2(_04268_),
    .B1(_04260_),
    .Y(_04374_));
 sky130_fd_sc_hd__a21bo_1 _11259_ (.A1(_04272_),
    .A2(_04275_),
    .B1_N(_04274_),
    .X(_04375_));
 sky130_fd_sc_hd__o21bai_2 _11260_ (.A1(_04263_),
    .A2(_04264_),
    .B1_N(_04266_),
    .Y(_04376_));
 sky130_fd_sc_hd__o22a_1 _11261_ (.A1(_04237_),
    .A2(_04247_),
    .B1(_04255_),
    .B2(_04258_),
    .X(_04377_));
 sky130_fd_sc_hd__or4_1 _11262_ (.A(_04237_),
    .B(_04247_),
    .C(_04255_),
    .D(_04258_),
    .X(_04378_));
 sky130_fd_sc_hd__and2b_1 _11263_ (.A_N(_04377_),
    .B(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__xnor2_1 _11264_ (.A(_04376_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2b_1 _11265_ (.A_N(_04380_),
    .B(_04375_),
    .Y(_04381_));
 sky130_fd_sc_hd__xnor2_1 _11266_ (.A(_04375_),
    .B(_04380_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2b_1 _11267_ (.A_N(_04374_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__xnor2_1 _11268_ (.A(_04374_),
    .B(_04382_),
    .Y(_04384_));
 sky130_fd_sc_hd__nand2_1 _11269_ (.A(_04373_),
    .B(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__xnor2_1 _11270_ (.A(_04373_),
    .B(_04384_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand2b_1 _11271_ (.A_N(_04386_),
    .B(_04333_),
    .Y(_04387_));
 sky130_fd_sc_hd__xnor2_1 _11272_ (.A(_04333_),
    .B(_04386_),
    .Y(_04388_));
 sky130_fd_sc_hd__o21a_1 _11273_ (.A1(_04282_),
    .A2(_04285_),
    .B1(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__nor3_1 _11274_ (.A(_04282_),
    .B(_04285_),
    .C(_04388_),
    .Y(_04390_));
 sky130_fd_sc_hd__or2_1 _11275_ (.A(_04389_),
    .B(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__o21ai_1 _11276_ (.A1(_04183_),
    .A2(_04287_),
    .B1(_04288_),
    .Y(_04392_));
 sky130_fd_sc_hd__nor2_1 _11277_ (.A(_04186_),
    .B(_04289_),
    .Y(_04393_));
 sky130_fd_sc_hd__a21bo_1 _11278_ (.A1(_04187_),
    .A2(_04393_),
    .B1_N(_04392_),
    .X(_04394_));
 sky130_fd_sc_hd__nand2_1 _11279_ (.A(_04188_),
    .B(_04393_),
    .Y(_04395_));
 sky130_fd_sc_hd__o21bai_1 _11280_ (.A1(_03974_),
    .A2(_04395_),
    .B1_N(_04394_),
    .Y(_04396_));
 sky130_fd_sc_hd__xnor2_1 _11281_ (.A(_04391_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__a21oi_1 _11282_ (.A1(_04332_),
    .A2(_04397_),
    .B1(_02242_),
    .Y(_04398_));
 sky130_fd_sc_hd__o21a_1 _11283_ (.A1(_04332_),
    .A2(_04397_),
    .B1(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__a21o_1 _11284_ (.A1(_02191_),
    .A2(_02192_),
    .B1(_02135_),
    .X(_04401_));
 sky130_fd_sc_hd__or2_1 _11285_ (.A(_02193_),
    .B(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__a21oi_1 _11286_ (.A1(_02193_),
    .A2(_04401_),
    .B1(_02318_),
    .Y(_04403_));
 sky130_fd_sc_hd__o21ai_1 _11287_ (.A1(_06089_),
    .A2(_04302_),
    .B1(_06083_),
    .Y(_04404_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(_06364_),
    .A1(_04404_),
    .S(net297),
    .X(_04405_));
 sky130_fd_sc_hd__xor2_1 _11289_ (.A(_06059_),
    .B(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__o21a_1 _11290_ (.A1(_04308_),
    .A2(_04309_),
    .B1(_04306_),
    .X(_04407_));
 sky130_fd_sc_hd__nor2_1 _11291_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04408_));
 sky130_fd_sc_hd__nand2_1 _11292_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04409_));
 sky130_fd_sc_hd__and2b_1 _11293_ (.A_N(_04408_),
    .B(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__xnor2_1 _11294_ (.A(_04407_),
    .B(_04410_),
    .Y(_04412_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(_04325_),
    .A1(_04412_),
    .S(net261),
    .X(_04413_));
 sky130_fd_sc_hd__or2_1 _11296_ (.A(\div_shifter[47] ),
    .B(_04315_),
    .X(_04414_));
 sky130_fd_sc_hd__a21o_1 _11297_ (.A1(net233),
    .A2(_04414_),
    .B1(\div_shifter[48] ),
    .X(_04415_));
 sky130_fd_sc_hd__a31oi_2 _11298_ (.A1(\div_shifter[48] ),
    .A2(net233),
    .A3(_04414_),
    .B1(net238),
    .Y(_04416_));
 sky130_fd_sc_hd__a2bb2o_1 _11299_ (.A1_N(reg1_val[16]),
    .A2_N(net236),
    .B1(_06020_),
    .B2(_06455_),
    .X(_04417_));
 sky130_fd_sc_hd__a221o_1 _11300_ (.A1(_06053_),
    .A2(net201),
    .B1(_02322_),
    .B2(_06042_),
    .C1(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__a221o_1 _11301_ (.A1(_06059_),
    .A2(net240),
    .B1(_04415_),
    .B2(_04416_),
    .C1(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__or2_1 _11302_ (.A(\div_res[15] ),
    .B(_04318_),
    .X(_04420_));
 sky130_fd_sc_hd__a21oi_1 _11303_ (.A1(net155),
    .A2(_04420_),
    .B1(\div_res[16] ),
    .Y(_04421_));
 sky130_fd_sc_hd__a31o_1 _11304_ (.A1(\div_res[16] ),
    .A2(net155),
    .A3(_04420_),
    .B1(net199),
    .X(_04423_));
 sky130_fd_sc_hd__o2bb2a_1 _11305_ (.A1_N(_02315_),
    .A2_N(_04325_),
    .B1(_04421_),
    .B2(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__o21ai_1 _11306_ (.A1(_02247_),
    .A2(_04313_),
    .B1(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__a211o_1 _11307_ (.A1(net210),
    .A2(_04413_),
    .B1(_04419_),
    .C1(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__a221o_2 _11308_ (.A1(_04402_),
    .A2(_04403_),
    .B1(_04406_),
    .B2(net242),
    .C1(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__o21a_1 _11309_ (.A1(_04399_),
    .A2(_04427_),
    .B1(net255),
    .X(_04428_));
 sky130_fd_sc_hd__nand2_1 _11310_ (.A(curr_PC[16]),
    .B(_04330_),
    .Y(_04429_));
 sky130_fd_sc_hd__or2_1 _11311_ (.A(curr_PC[16]),
    .B(_04330_),
    .X(_04430_));
 sky130_fd_sc_hd__a31o_4 _11312_ (.A1(net258),
    .A2(_04429_),
    .A3(_04430_),
    .B1(_04428_),
    .X(dest_val[16]));
 sky130_fd_sc_hd__a21oi_1 _11313_ (.A1(curr_PC[16]),
    .A2(_04330_),
    .B1(curr_PC[17]),
    .Y(_04431_));
 sky130_fd_sc_hd__and3_1 _11314_ (.A(curr_PC[16]),
    .B(curr_PC[17]),
    .C(_04330_),
    .X(_04433_));
 sky130_fd_sc_hd__o21ai_1 _11315_ (.A1(_04431_),
    .A2(_04433_),
    .B1(net258),
    .Y(_04434_));
 sky130_fd_sc_hd__or4b_2 _11316_ (.A(_03894_),
    .B(_04397_),
    .C(_04331_),
    .D_N(_03645_),
    .X(_04435_));
 sky130_fd_sc_hd__and2_1 _11317_ (.A(net157),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__o22a_1 _11318_ (.A1(net19),
    .A2(net47),
    .B1(net11),
    .B2(net23),
    .X(_04437_));
 sky130_fd_sc_hd__xnor2_1 _11319_ (.A(net110),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__nor2_1 _11320_ (.A(net88),
    .B(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__xnor2_1 _11321_ (.A(net88),
    .B(_04438_),
    .Y(_04440_));
 sky130_fd_sc_hd__o22a_1 _11322_ (.A1(net17),
    .A2(net13),
    .B1(net8),
    .B2(net48),
    .X(_04441_));
 sky130_fd_sc_hd__xor2_1 _11323_ (.A(net87),
    .B(_04441_),
    .X(_04442_));
 sky130_fd_sc_hd__nor2_1 _11324_ (.A(_04440_),
    .B(_04442_),
    .Y(_04444_));
 sky130_fd_sc_hd__xnor2_1 _11325_ (.A(_04440_),
    .B(_04442_),
    .Y(_04445_));
 sky130_fd_sc_hd__nor2_1 _11326_ (.A(_04365_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__xor2_1 _11327_ (.A(_04365_),
    .B(_04445_),
    .X(_04447_));
 sky130_fd_sc_hd__and3_1 _11328_ (.A(_04354_),
    .B(_04356_),
    .C(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__a21oi_1 _11329_ (.A1(_04354_),
    .A2(_04356_),
    .B1(_04447_),
    .Y(_04449_));
 sky130_fd_sc_hd__nor2_1 _11330_ (.A(_04448_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__o22a_1 _11331_ (.A1(net35),
    .A2(net78),
    .B1(net63),
    .B2(net37),
    .X(_04451_));
 sky130_fd_sc_hd__xnor2_1 _11332_ (.A(net120),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__o22a_1 _11333_ (.A1(net79),
    .A2(net21),
    .B1(net60),
    .B2(net33),
    .X(_04453_));
 sky130_fd_sc_hd__xnor2_1 _11334_ (.A(net113),
    .B(_04453_),
    .Y(_04455_));
 sky130_fd_sc_hd__and2_1 _11335_ (.A(_04452_),
    .B(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__nor2_1 _11336_ (.A(_04452_),
    .B(_04455_),
    .Y(_04457_));
 sky130_fd_sc_hd__nor2_1 _11337_ (.A(_04456_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__o22a_1 _11338_ (.A1(net29),
    .A2(net64),
    .B1(net59),
    .B2(net32),
    .X(_04459_));
 sky130_fd_sc_hd__xnor2_2 _11339_ (.A(net116),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__xor2_2 _11340_ (.A(_04458_),
    .B(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__nand2_1 _11341_ (.A(_04450_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__xnor2_2 _11342_ (.A(_04450_),
    .B(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__o22a_1 _11343_ (.A1(net70),
    .A2(net15),
    .B1(net6),
    .B2(net108),
    .X(_04464_));
 sky130_fd_sc_hd__xnor2_2 _11344_ (.A(net41),
    .B(_04464_),
    .Y(_04466_));
 sky130_fd_sc_hd__o22a_1 _11345_ (.A1(net74),
    .A2(net27),
    .B1(net25),
    .B2(net71),
    .X(_04467_));
 sky130_fd_sc_hd__xnor2_1 _11346_ (.A(net66),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__or3_1 _11347_ (.A(net104),
    .B(net39),
    .C(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__o21ai_1 _11348_ (.A1(net104),
    .A2(net39),
    .B1(_04468_),
    .Y(_04470_));
 sky130_fd_sc_hd__and2_1 _11349_ (.A(_04469_),
    .B(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__xnor2_2 _11350_ (.A(_04466_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__xor2_2 _11351_ (.A(_04463_),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__a21bo_1 _11352_ (.A1(_04340_),
    .A2(_04372_),
    .B1_N(_04371_),
    .X(_04474_));
 sky130_fd_sc_hd__a21o_1 _11353_ (.A1(_04334_),
    .A2(_04336_),
    .B1(_04338_),
    .X(_04475_));
 sky130_fd_sc_hd__or2_1 _11354_ (.A(_04345_),
    .B(_04350_),
    .X(_04477_));
 sky130_fd_sc_hd__o21a_1 _11355_ (.A1(_04359_),
    .A2(_04368_),
    .B1(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__or3_1 _11356_ (.A(_04359_),
    .B(_04368_),
    .C(_04477_),
    .X(_04479_));
 sky130_fd_sc_hd__and2b_1 _11357_ (.A_N(_04478_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__xnor2_1 _11358_ (.A(_04475_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__a21oi_1 _11359_ (.A1(_04376_),
    .A2(_04379_),
    .B1(_04377_),
    .Y(_04482_));
 sky130_fd_sc_hd__xnor2_1 _11360_ (.A(_04481_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__and2b_1 _11361_ (.A_N(_04483_),
    .B(_04474_),
    .X(_04484_));
 sky130_fd_sc_hd__xnor2_1 _11362_ (.A(_04474_),
    .B(_04483_),
    .Y(_04485_));
 sky130_fd_sc_hd__nand2_1 _11363_ (.A(_04473_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__xnor2_1 _11364_ (.A(_04473_),
    .B(_04485_),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_1 _11365_ (.A(_04381_),
    .B(_04383_),
    .Y(_04489_));
 sky130_fd_sc_hd__nand2b_1 _11366_ (.A_N(_04488_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__xor2_1 _11367_ (.A(_04488_),
    .B(_04489_),
    .X(_04491_));
 sky130_fd_sc_hd__a21oi_1 _11368_ (.A1(_04385_),
    .A2(_04387_),
    .B1(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__nand3_1 _11369_ (.A(_04385_),
    .B(_04387_),
    .C(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2b_2 _11370_ (.A_N(_04492_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__o21ba_1 _11371_ (.A1(_04287_),
    .A2(_04389_),
    .B1_N(_04390_),
    .X(_04495_));
 sky130_fd_sc_hd__nor2_1 _11372_ (.A(_04289_),
    .B(_04391_),
    .Y(_04496_));
 sky130_fd_sc_hd__a21oi_1 _11373_ (.A1(_04292_),
    .A2(_04496_),
    .B1(_04495_),
    .Y(_04497_));
 sky130_fd_sc_hd__nand2_1 _11374_ (.A(_04290_),
    .B(_04496_),
    .Y(_04499_));
 sky130_fd_sc_hd__o21ai_2 _11375_ (.A1(_04083_),
    .A2(_04499_),
    .B1(_04497_),
    .Y(_04500_));
 sky130_fd_sc_hd__xnor2_2 _11376_ (.A(_04494_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__o21ai_1 _11377_ (.A1(_04436_),
    .A2(_04501_),
    .B1(net202),
    .Y(_04502_));
 sky130_fd_sc_hd__a21oi_1 _11378_ (.A1(_04436_),
    .A2(_04501_),
    .B1(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__or3_1 _11379_ (.A(_02135_),
    .B(_02194_),
    .C(_02195_),
    .X(_04504_));
 sky130_fd_sc_hd__o21ai_1 _11380_ (.A1(_02135_),
    .A2(_02194_),
    .B1(_02195_),
    .Y(_04505_));
 sky130_fd_sc_hd__and3_2 _11381_ (.A(_02317_),
    .B(_04504_),
    .C(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__a21o_1 _11382_ (.A1(_06042_),
    .A2(_04404_),
    .B1(_06053_),
    .X(_04507_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(_06366_),
    .A1(_04507_),
    .S(net297),
    .X(_04508_));
 sky130_fd_sc_hd__a21oi_1 _11384_ (.A1(_05976_),
    .A2(_04508_),
    .B1(net241),
    .Y(_04510_));
 sky130_fd_sc_hd__o21a_1 _11385_ (.A1(_05976_),
    .A2(_04508_),
    .B1(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__o21a_1 _11386_ (.A1(_04407_),
    .A2(_04408_),
    .B1(_04409_),
    .X(_04512_));
 sky130_fd_sc_hd__nor2_1 _11387_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04513_));
 sky130_fd_sc_hd__nand2_1 _11388_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2b_1 _11389_ (.A_N(_04513_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__xor2_1 _11390_ (.A(_04512_),
    .B(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__or2_1 _11391_ (.A(net261),
    .B(_04221_),
    .X(_04517_));
 sky130_fd_sc_hd__o211a_1 _11392_ (.A1(net229),
    .A2(_04516_),
    .B1(_04517_),
    .C1(_06446_),
    .X(_04518_));
 sky130_fd_sc_hd__o21ai_1 _11393_ (.A1(reg1_val[17]),
    .A2(net236),
    .B1(net257),
    .Y(_04519_));
 sky130_fd_sc_hd__a221o_1 _11394_ (.A1(_05935_),
    .A2(_06455_),
    .B1(_02322_),
    .B2(_05954_),
    .C1(_04519_),
    .X(_04521_));
 sky130_fd_sc_hd__a221o_1 _11395_ (.A1(_05965_),
    .A2(net201),
    .B1(net240),
    .B2(_05976_),
    .C1(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__a221o_1 _11396_ (.A1(net246),
    .A2(_04210_),
    .B1(_04221_),
    .B2(_02315_),
    .C1(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__or2_1 _11397_ (.A(\div_shifter[48] ),
    .B(_04414_),
    .X(_04524_));
 sky130_fd_sc_hd__and3_1 _11398_ (.A(\div_shifter[49] ),
    .B(net233),
    .C(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__a21oi_1 _11399_ (.A1(net233),
    .A2(_04524_),
    .B1(\div_shifter[49] ),
    .Y(_04526_));
 sky130_fd_sc_hd__or3_1 _11400_ (.A(net238),
    .B(_04525_),
    .C(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__o21a_1 _11401_ (.A1(\div_res[16] ),
    .A2(_04420_),
    .B1(net154),
    .X(_04528_));
 sky130_fd_sc_hd__xnor2_1 _11402_ (.A(\div_res[17] ),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__o21ai_1 _11403_ (.A1(net198),
    .A2(_04529_),
    .B1(_04527_),
    .Y(_04530_));
 sky130_fd_sc_hd__or4_2 _11404_ (.A(_04511_),
    .B(_04518_),
    .C(_04523_),
    .D(_04530_),
    .X(_04532_));
 sky130_fd_sc_hd__o31a_4 _11405_ (.A1(_04503_),
    .A2(_04506_),
    .A3(_04532_),
    .B1(_04434_),
    .X(dest_val[17]));
 sky130_fd_sc_hd__o21a_1 _11406_ (.A1(_04435_),
    .A2(_04501_),
    .B1(net157),
    .X(_04533_));
 sky130_fd_sc_hd__o21bai_1 _11407_ (.A1(_04481_),
    .A2(_04482_),
    .B1_N(_04484_),
    .Y(_04534_));
 sky130_fd_sc_hd__o22a_1 _11408_ (.A1(net78),
    .A2(net27),
    .B1(net25),
    .B2(net74),
    .X(_04535_));
 sky130_fd_sc_hd__xnor2_2 _11409_ (.A(net66),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__o22a_1 _11410_ (.A1(net71),
    .A2(net15),
    .B1(net6),
    .B2(net70),
    .X(_04537_));
 sky130_fd_sc_hd__xnor2_2 _11411_ (.A(net41),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__o22a_1 _11412_ (.A1(net37),
    .A2(net64),
    .B1(net63),
    .B2(net35),
    .X(_04539_));
 sky130_fd_sc_hd__xnor2_2 _11413_ (.A(net120),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__xor2_2 _11414_ (.A(_04538_),
    .B(_04540_),
    .X(_04542_));
 sky130_fd_sc_hd__nand2b_1 _11415_ (.A_N(_04536_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__xor2_2 _11416_ (.A(_04536_),
    .B(_04542_),
    .X(_04544_));
 sky130_fd_sc_hd__o22a_1 _11417_ (.A1(net32),
    .A2(net60),
    .B1(net59),
    .B2(net29),
    .X(_04545_));
 sky130_fd_sc_hd__xnor2_1 _11418_ (.A(net116),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__o22a_1 _11419_ (.A1(net17),
    .A2(net47),
    .B1(net11),
    .B2(net19),
    .X(_04547_));
 sky130_fd_sc_hd__xnor2_1 _11420_ (.A(net112),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand2_1 _11421_ (.A(_04546_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__or2_1 _11422_ (.A(_04546_),
    .B(_04548_),
    .X(_04550_));
 sky130_fd_sc_hd__and2_1 _11423_ (.A(_04549_),
    .B(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__o22a_1 _11424_ (.A1(net79),
    .A2(net23),
    .B1(net21),
    .B2(net33),
    .X(_04553_));
 sky130_fd_sc_hd__xnor2_1 _11425_ (.A(net113),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nand2_1 _11426_ (.A(_04551_),
    .B(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__or2_1 _11427_ (.A(_04551_),
    .B(_04554_),
    .X(_04556_));
 sky130_fd_sc_hd__and2_1 _11428_ (.A(_04555_),
    .B(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__or3_1 _11429_ (.A(net88),
    .B(_00432_),
    .C(net9),
    .X(_04558_));
 sky130_fd_sc_hd__a2bb2o_2 _11430_ (.A1_N(_00439_),
    .A2_N(net9),
    .B1(_04558_),
    .B2(net85),
    .X(_04559_));
 sky130_fd_sc_hd__nor2_1 _11431_ (.A(net108),
    .B(net39),
    .Y(_04560_));
 sky130_fd_sc_hd__xnor2_1 _11432_ (.A(_04559_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__o21ai_1 _11433_ (.A1(_04439_),
    .A2(_04444_),
    .B1(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__or3_1 _11434_ (.A(_04439_),
    .B(_04444_),
    .C(_04561_),
    .X(_04564_));
 sky130_fd_sc_hd__and2_1 _11435_ (.A(_04562_),
    .B(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__nand2_1 _11436_ (.A(_04557_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__or2_1 _11437_ (.A(_04557_),
    .B(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__nand2_1 _11438_ (.A(_04566_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__xnor2_1 _11439_ (.A(_04544_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__o21ai_1 _11440_ (.A1(_04463_),
    .A2(_04472_),
    .B1(_04462_),
    .Y(_04570_));
 sky130_fd_sc_hd__a21bo_1 _11441_ (.A1(_04466_),
    .A2(_04471_),
    .B1_N(_04469_),
    .X(_04571_));
 sky130_fd_sc_hd__a21oi_1 _11442_ (.A1(_04458_),
    .A2(_04460_),
    .B1(_04456_),
    .Y(_04572_));
 sky130_fd_sc_hd__o21ba_1 _11443_ (.A1(_04446_),
    .A2(_04448_),
    .B1_N(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__or3b_1 _11444_ (.A(_04446_),
    .B(_04448_),
    .C_N(_04572_),
    .X(_04575_));
 sky130_fd_sc_hd__and2b_1 _11445_ (.A_N(_04573_),
    .B(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__xnor2_1 _11446_ (.A(_04571_),
    .B(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__a21o_1 _11447_ (.A1(_04475_),
    .A2(_04479_),
    .B1(_04478_),
    .X(_04578_));
 sky130_fd_sc_hd__and2b_1 _11448_ (.A_N(_04577_),
    .B(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__xnor2_1 _11449_ (.A(_04577_),
    .B(_04578_),
    .Y(_04580_));
 sky130_fd_sc_hd__and2_1 _11450_ (.A(_04570_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__xnor2_1 _11451_ (.A(_04570_),
    .B(_04580_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _11452_ (.A(_04569_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__xor2_1 _11453_ (.A(_04569_),
    .B(_04582_),
    .X(_04584_));
 sky130_fd_sc_hd__and2_1 _11454_ (.A(_04534_),
    .B(_04584_),
    .X(_04586_));
 sky130_fd_sc_hd__xnor2_1 _11455_ (.A(_04534_),
    .B(_04584_),
    .Y(_04587_));
 sky130_fd_sc_hd__a21oi_1 _11456_ (.A1(_04486_),
    .A2(_04490_),
    .B1(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__nand3_1 _11457_ (.A(_04486_),
    .B(_04490_),
    .C(_04587_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2b_2 _11458_ (.A_N(_04588_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21ai_1 _11459_ (.A1(_04389_),
    .A2(_04492_),
    .B1(_04493_),
    .Y(_04591_));
 sky130_fd_sc_hd__or2_1 _11460_ (.A(_04391_),
    .B(_04494_),
    .X(_04592_));
 sky130_fd_sc_hd__o21ai_1 _11461_ (.A1(_04392_),
    .A2(_04592_),
    .B1(_04591_),
    .Y(_04593_));
 sky130_fd_sc_hd__nor3_1 _11462_ (.A(_04186_),
    .B(_04289_),
    .C(_04592_),
    .Y(_04594_));
 sky130_fd_sc_hd__a21o_1 _11463_ (.A1(_04190_),
    .A2(_04594_),
    .B1(_04593_),
    .X(_04595_));
 sky130_fd_sc_hd__xnor2_2 _11464_ (.A(_04590_),
    .B(_04595_),
    .Y(_04597_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(_04533_),
    .A2(_04597_),
    .B1(net202),
    .Y(_04598_));
 sky130_fd_sc_hd__a21o_1 _11466_ (.A1(_04533_),
    .A2(_04597_),
    .B1(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__a21o_1 _11467_ (.A1(_02194_),
    .A2(_02195_),
    .B1(net150),
    .X(_04600_));
 sky130_fd_sc_hd__xnor2_1 _11468_ (.A(_02196_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__a21o_1 _11469_ (.A1(_05954_),
    .A2(_04507_),
    .B1(_05965_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_1 _11470_ (.A(net297),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__o21ai_1 _11471_ (.A1(net297),
    .A2(_06368_),
    .B1(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__o21ai_1 _11472_ (.A1(_05905_),
    .A2(_04604_),
    .B1(net242),
    .Y(_04605_));
 sky130_fd_sc_hd__a21o_1 _11473_ (.A1(_05905_),
    .A2(_04604_),
    .B1(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2_1 _11474_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04608_));
 sky130_fd_sc_hd__or2_1 _11475_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .X(_04609_));
 sky130_fd_sc_hd__nand2_1 _11476_ (.A(_04608_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__o21ai_1 _11477_ (.A1(_04512_),
    .A2(_04513_),
    .B1(_04514_),
    .Y(_04611_));
 sky130_fd_sc_hd__xor2_1 _11478_ (.A(_04610_),
    .B(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(_04111_),
    .A1(_04612_),
    .S(net261),
    .X(_04613_));
 sky130_fd_sc_hd__or3_1 _11480_ (.A(\div_res[17] ),
    .B(\div_res[16] ),
    .C(_04420_),
    .X(_04614_));
 sky130_fd_sc_hd__a21oi_1 _11481_ (.A1(net154),
    .A2(_04614_),
    .B1(\div_res[18] ),
    .Y(_04615_));
 sky130_fd_sc_hd__a311o_1 _11482_ (.A1(\div_res[18] ),
    .A2(net154),
    .A3(_04614_),
    .B1(_04615_),
    .C1(net199),
    .X(_04616_));
 sky130_fd_sc_hd__or2_1 _11483_ (.A(\div_shifter[49] ),
    .B(_04524_),
    .X(_04617_));
 sky130_fd_sc_hd__a21oi_1 _11484_ (.A1(net232),
    .A2(_04617_),
    .B1(\div_shifter[50] ),
    .Y(_04619_));
 sky130_fd_sc_hd__a311o_1 _11485_ (.A1(\div_shifter[50] ),
    .A2(net232),
    .A3(_04617_),
    .B1(_04619_),
    .C1(net238),
    .X(_04620_));
 sky130_fd_sc_hd__a21oi_1 _11486_ (.A1(_05890_),
    .A2(net240),
    .B1(net273),
    .Y(_04621_));
 sky130_fd_sc_hd__o22a_1 _11487_ (.A1(_05863_),
    .A2(net252),
    .B1(net237),
    .B2(reg1_val[18]),
    .X(_04622_));
 sky130_fd_sc_hd__o221a_1 _11488_ (.A1(_05890_),
    .A2(_02320_),
    .B1(_04621_),
    .B2(_05899_),
    .C1(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__o221a_1 _11489_ (.A1(_02247_),
    .A2(_04100_),
    .B1(_04111_),
    .B2(_02316_),
    .C1(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__and3_1 _11490_ (.A(_04616_),
    .B(_04620_),
    .C(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__o211a_1 _11491_ (.A1(net209),
    .A2(_04613_),
    .B1(_04625_),
    .C1(_04606_),
    .X(_04626_));
 sky130_fd_sc_hd__o211a_1 _11492_ (.A1(_02318_),
    .A2(_04601_),
    .B1(_04626_),
    .C1(_04599_),
    .X(_04627_));
 sky130_fd_sc_hd__and2_2 _11493_ (.A(curr_PC[18]),
    .B(_04433_),
    .X(_04628_));
 sky130_fd_sc_hd__o21ai_2 _11494_ (.A1(curr_PC[18]),
    .A2(_04433_),
    .B1(net258),
    .Y(_04630_));
 sky130_fd_sc_hd__o22ai_4 _11495_ (.A1(net258),
    .A2(_04627_),
    .B1(_04628_),
    .B2(_04630_),
    .Y(dest_val[18]));
 sky130_fd_sc_hd__o22a_1 _11496_ (.A1(net33),
    .A2(net23),
    .B1(net19),
    .B2(net79),
    .X(_04631_));
 sky130_fd_sc_hd__xor2_1 _11497_ (.A(net113),
    .B(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__nor2_1 _11498_ (.A(net87),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__and2_1 _11499_ (.A(net87),
    .B(_04632_),
    .X(_04634_));
 sky130_fd_sc_hd__or2_1 _11500_ (.A(_04633_),
    .B(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__o22a_1 _11501_ (.A1(net17),
    .A2(net11),
    .B1(net8),
    .B2(net47),
    .X(_04636_));
 sky130_fd_sc_hd__xnor2_1 _11502_ (.A(net112),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__and2b_1 _11503_ (.A_N(_04635_),
    .B(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__and2b_1 _11504_ (.A_N(_04637_),
    .B(_04635_),
    .X(_04640_));
 sky130_fd_sc_hd__or2_1 _11505_ (.A(_04638_),
    .B(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__o22a_1 _11506_ (.A1(net74),
    .A2(net15),
    .B1(net6),
    .B2(net71),
    .X(_04642_));
 sky130_fd_sc_hd__xnor2_1 _11507_ (.A(net41),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__and2_1 _11508_ (.A(_04559_),
    .B(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__nor2_1 _11509_ (.A(_04559_),
    .B(_04643_),
    .Y(_04645_));
 sky130_fd_sc_hd__or2_1 _11510_ (.A(_04644_),
    .B(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(_00211_),
    .B(net41),
    .Y(_04647_));
 sky130_fd_sc_hd__nor2_1 _11512_ (.A(_04646_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__and2_1 _11513_ (.A(_04646_),
    .B(_04647_),
    .X(_04649_));
 sky130_fd_sc_hd__nor2_1 _11514_ (.A(_04648_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__and2b_1 _11515_ (.A_N(_04641_),
    .B(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__xnor2_1 _11516_ (.A(_04641_),
    .B(_04650_),
    .Y(_04652_));
 sky130_fd_sc_hd__o22a_1 _11517_ (.A1(net78),
    .A2(net25),
    .B1(net63),
    .B2(net27),
    .X(_04653_));
 sky130_fd_sc_hd__xnor2_1 _11518_ (.A(net66),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o22a_1 _11519_ (.A1(net32),
    .A2(net21),
    .B1(net60),
    .B2(net29),
    .X(_04655_));
 sky130_fd_sc_hd__xnor2_1 _11520_ (.A(net116),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__and2b_1 _11521_ (.A_N(_04654_),
    .B(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__xor2_1 _11522_ (.A(_04654_),
    .B(_04656_),
    .X(_04658_));
 sky130_fd_sc_hd__o22a_1 _11523_ (.A1(net35),
    .A2(net64),
    .B1(net59),
    .B2(net37),
    .X(_04659_));
 sky130_fd_sc_hd__xnor2_1 _11524_ (.A(net120),
    .B(_04659_),
    .Y(_04661_));
 sky130_fd_sc_hd__and2b_1 _11525_ (.A_N(_04658_),
    .B(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__and2b_1 _11526_ (.A_N(_04661_),
    .B(_04658_),
    .X(_04663_));
 sky130_fd_sc_hd__or2_1 _11527_ (.A(_04662_),
    .B(_04663_),
    .X(_04664_));
 sky130_fd_sc_hd__inv_2 _11528_ (.A(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__xnor2_1 _11529_ (.A(_04652_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__o21ai_1 _11530_ (.A1(_04544_),
    .A2(_04568_),
    .B1(_04566_),
    .Y(_04667_));
 sky130_fd_sc_hd__a21bo_1 _11531_ (.A1(_04538_),
    .A2(_04540_),
    .B1_N(_04543_),
    .X(_04668_));
 sky130_fd_sc_hd__nand2_1 _11532_ (.A(_04549_),
    .B(_04555_),
    .Y(_04669_));
 sky130_fd_sc_hd__o31a_1 _11533_ (.A1(net108),
    .A2(net39),
    .A3(_04559_),
    .B1(_04562_),
    .X(_04670_));
 sky130_fd_sc_hd__a21oi_1 _11534_ (.A1(_04549_),
    .A2(_04555_),
    .B1(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__xnor2_1 _11535_ (.A(_04669_),
    .B(_04670_),
    .Y(_04672_));
 sky130_fd_sc_hd__xnor2_1 _11536_ (.A(_04668_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__a21oi_1 _11537_ (.A1(_04571_),
    .A2(_04575_),
    .B1(_04573_),
    .Y(_04674_));
 sky130_fd_sc_hd__nor2_1 _11538_ (.A(_04673_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__xor2_1 _11539_ (.A(_04673_),
    .B(_04674_),
    .X(_04676_));
 sky130_fd_sc_hd__xnor2_1 _11540_ (.A(_04667_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__or2_1 _11541_ (.A(_04666_),
    .B(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__xor2_1 _11542_ (.A(_04666_),
    .B(_04677_),
    .X(_04679_));
 sky130_fd_sc_hd__o21ai_1 _11543_ (.A1(_04579_),
    .A2(_04581_),
    .B1(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__or3_1 _11544_ (.A(_04579_),
    .B(_04581_),
    .C(_04679_),
    .X(_04682_));
 sky130_fd_sc_hd__and2_1 _11545_ (.A(_04680_),
    .B(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__o21a_1 _11546_ (.A1(_04583_),
    .A2(_04586_),
    .B1(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__nor3_1 _11547_ (.A(_04583_),
    .B(_04586_),
    .C(_04683_),
    .Y(_04685_));
 sky130_fd_sc_hd__or2_1 _11548_ (.A(_04684_),
    .B(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__o21a_1 _11549_ (.A1(_04492_),
    .A2(_04588_),
    .B1(_04589_),
    .X(_04687_));
 sky130_fd_sc_hd__nor2_1 _11550_ (.A(_04494_),
    .B(_04590_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21o_1 _11551_ (.A1(_04495_),
    .A2(_04688_),
    .B1(_04687_),
    .X(_04689_));
 sky130_fd_sc_hd__and2_1 _11552_ (.A(_04496_),
    .B(_04688_),
    .X(_04690_));
 sky130_fd_sc_hd__a21o_1 _11553_ (.A1(_04295_),
    .A2(_04690_),
    .B1(_04689_),
    .X(_04691_));
 sky130_fd_sc_hd__xnor2_1 _11554_ (.A(_04686_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__o31a_1 _11555_ (.A1(_04435_),
    .A2(_04501_),
    .A3(_04597_),
    .B1(net157),
    .X(_04693_));
 sky130_fd_sc_hd__a21oi_1 _11556_ (.A1(_04692_),
    .A2(_04693_),
    .B1(_02242_),
    .Y(_04694_));
 sky130_fd_sc_hd__o21a_1 _11557_ (.A1(_04692_),
    .A2(_04693_),
    .B1(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__a21o_1 _11558_ (.A1(net155),
    .A2(_02197_),
    .B1(_02198_),
    .X(_04696_));
 sky130_fd_sc_hd__nand3_1 _11559_ (.A(net156),
    .B(_02197_),
    .C(_02198_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21o_1 _11560_ (.A1(_05905_),
    .A2(_04602_),
    .B1(_05881_),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(_06370_),
    .A1(_04698_),
    .S(net297),
    .X(_04699_));
 sky130_fd_sc_hd__o21ai_1 _11562_ (.A1(_05836_),
    .A2(_04699_),
    .B1(net242),
    .Y(_04700_));
 sky130_fd_sc_hd__a21o_1 _11563_ (.A1(_05836_),
    .A2(_04699_),
    .B1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__nand2_1 _11564_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04703_));
 sky130_fd_sc_hd__or2_1 _11565_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .X(_04704_));
 sky130_fd_sc_hd__nand2_1 _11566_ (.A(_04703_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__a21boi_1 _11567_ (.A1(_04609_),
    .A2(_04611_),
    .B1_N(_04608_),
    .Y(_04706_));
 sky130_fd_sc_hd__xnor2_1 _11568_ (.A(_04705_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__mux2_1 _11569_ (.A0(_04003_),
    .A1(_04707_),
    .S(net261),
    .X(_04708_));
 sky130_fd_sc_hd__or2_1 _11570_ (.A(\div_shifter[50] ),
    .B(_04617_),
    .X(_04709_));
 sky130_fd_sc_hd__a21oi_1 _11571_ (.A1(net232),
    .A2(_04709_),
    .B1(\div_shifter[51] ),
    .Y(_04710_));
 sky130_fd_sc_hd__a311o_1 _11572_ (.A1(\div_shifter[51] ),
    .A2(net232),
    .A3(_04709_),
    .B1(_04710_),
    .C1(net238),
    .X(_04711_));
 sky130_fd_sc_hd__or2_1 _11573_ (.A(\div_res[18] ),
    .B(_04614_),
    .X(_04712_));
 sky130_fd_sc_hd__a21oi_1 _11574_ (.A1(net154),
    .A2(_04712_),
    .B1(\div_res[19] ),
    .Y(_04713_));
 sky130_fd_sc_hd__a31o_1 _11575_ (.A1(\div_res[19] ),
    .A2(net156),
    .A3(_04712_),
    .B1(net199),
    .X(_04714_));
 sky130_fd_sc_hd__o21a_1 _11576_ (.A1(_05810_),
    .A2(_02327_),
    .B1(_02323_),
    .X(_04715_));
 sky130_fd_sc_hd__o22a_1 _11577_ (.A1(_05800_),
    .A2(net251),
    .B1(net236),
    .B2(reg1_val[19]),
    .X(_04716_));
 sky130_fd_sc_hd__o221a_1 _11578_ (.A1(_05819_),
    .A2(net200),
    .B1(_04715_),
    .B2(_05828_),
    .C1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__o221a_1 _11579_ (.A1(_02247_),
    .A2(_03987_),
    .B1(_04003_),
    .B2(_02316_),
    .C1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__o211a_1 _11580_ (.A1(_04713_),
    .A2(_04714_),
    .B1(_04718_),
    .C1(_04711_),
    .X(_04719_));
 sky130_fd_sc_hd__o211ai_1 _11581_ (.A1(net209),
    .A2(_04708_),
    .B1(_04719_),
    .C1(_04701_),
    .Y(_04720_));
 sky130_fd_sc_hd__a311o_2 _11582_ (.A1(_02317_),
    .A2(_04696_),
    .A3(_04697_),
    .B1(_04720_),
    .C1(_04695_),
    .X(_04721_));
 sky130_fd_sc_hd__or2_1 _11583_ (.A(curr_PC[19]),
    .B(_04628_),
    .X(_04722_));
 sky130_fd_sc_hd__a21oi_1 _11584_ (.A1(curr_PC[19]),
    .A2(_04628_),
    .B1(net253),
    .Y(_04724_));
 sky130_fd_sc_hd__a22o_4 _11585_ (.A1(net255),
    .A2(_04721_),
    .B1(_04722_),
    .B2(_04724_),
    .X(dest_val[19]));
 sky130_fd_sc_hd__or2_1 _11586_ (.A(_04597_),
    .B(_04692_),
    .X(_04725_));
 sky130_fd_sc_hd__nor3_1 _11587_ (.A(_04435_),
    .B(_04501_),
    .C(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__nor2_1 _11588_ (.A(net149),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__a21o_1 _11589_ (.A1(_04667_),
    .A2(_04676_),
    .B1(_04675_),
    .X(_04728_));
 sky130_fd_sc_hd__o22a_1 _11590_ (.A1(net27),
    .A2(net64),
    .B1(net63),
    .B2(net25),
    .X(_04729_));
 sky130_fd_sc_hd__xnor2_1 _11591_ (.A(net66),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__o22a_1 _11592_ (.A1(net32),
    .A2(net23),
    .B1(net21),
    .B2(net29),
    .X(_04731_));
 sky130_fd_sc_hd__xnor2_1 _11593_ (.A(net116),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__and2b_1 _11594_ (.A_N(_04730_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__xor2_1 _11595_ (.A(_04730_),
    .B(_04732_),
    .X(_04734_));
 sky130_fd_sc_hd__o22a_1 _11596_ (.A1(net37),
    .A2(net60),
    .B1(net59),
    .B2(net35),
    .X(_04735_));
 sky130_fd_sc_hd__xnor2_1 _11597_ (.A(net120),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__and2b_1 _11598_ (.A_N(_04734_),
    .B(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__and2b_1 _11599_ (.A_N(_04736_),
    .B(_04734_),
    .X(_04738_));
 sky130_fd_sc_hd__or2_1 _11600_ (.A(_04737_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__o22a_1 _11601_ (.A1(net33),
    .A2(net19),
    .B1(net17),
    .B2(net79),
    .X(_04740_));
 sky130_fd_sc_hd__xnor2_1 _11602_ (.A(net113),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_1 _11603_ (.A(net11),
    .B(net8),
    .Y(_04742_));
 sky130_fd_sc_hd__xnor2_1 _11604_ (.A(net112),
    .B(_04742_),
    .Y(_04744_));
 sky130_fd_sc_hd__and2b_1 _11605_ (.A_N(_04741_),
    .B(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__and2b_1 _11606_ (.A_N(_04744_),
    .B(_04741_),
    .X(_04746_));
 sky130_fd_sc_hd__or2_1 _11607_ (.A(_04745_),
    .B(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__o22a_1 _11608_ (.A1(net78),
    .A2(net15),
    .B1(net6),
    .B2(net74),
    .X(_04748_));
 sky130_fd_sc_hd__nand2_1 _11609_ (.A(net71),
    .B(net41),
    .Y(_04749_));
 sky130_fd_sc_hd__xor2_1 _11610_ (.A(_04748_),
    .B(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__nand2_1 _11611_ (.A(_04747_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__or2_1 _11612_ (.A(_04747_),
    .B(_04750_),
    .X(_04752_));
 sky130_fd_sc_hd__nand2_1 _11613_ (.A(_04751_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__xor2_1 _11614_ (.A(_04739_),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a21o_1 _11615_ (.A1(_04652_),
    .A2(_04665_),
    .B1(_04651_),
    .X(_04755_));
 sky130_fd_sc_hd__or2_1 _11616_ (.A(_04657_),
    .B(_04662_),
    .X(_04756_));
 sky130_fd_sc_hd__o22ai_1 _11617_ (.A1(_04633_),
    .A2(_04638_),
    .B1(_04644_),
    .B2(_04648_),
    .Y(_04757_));
 sky130_fd_sc_hd__or4_1 _11618_ (.A(_04633_),
    .B(_04638_),
    .C(_04644_),
    .D(_04648_),
    .X(_04758_));
 sky130_fd_sc_hd__and2_1 _11619_ (.A(_04757_),
    .B(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__xnor2_1 _11620_ (.A(_04756_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__a21oi_1 _11621_ (.A1(_04668_),
    .A2(_04672_),
    .B1(_04671_),
    .Y(_04761_));
 sky130_fd_sc_hd__xnor2_1 _11622_ (.A(_04760_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__and2b_1 _11623_ (.A_N(_04762_),
    .B(_04755_),
    .X(_04763_));
 sky130_fd_sc_hd__xnor2_1 _11624_ (.A(_04755_),
    .B(_04762_),
    .Y(_04765_));
 sky130_fd_sc_hd__and2_1 _11625_ (.A(_04754_),
    .B(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__nor2_1 _11626_ (.A(_04754_),
    .B(_04765_),
    .Y(_04767_));
 sky130_fd_sc_hd__or2_1 _11627_ (.A(_04766_),
    .B(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__and2b_1 _11628_ (.A_N(_04768_),
    .B(_04728_),
    .X(_04769_));
 sky130_fd_sc_hd__xor2_1 _11629_ (.A(_04728_),
    .B(_04768_),
    .X(_04770_));
 sky130_fd_sc_hd__a21o_1 _11630_ (.A1(_04678_),
    .A2(_04680_),
    .B1(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__inv_2 _11631_ (.A(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand3_1 _11632_ (.A(_04678_),
    .B(_04680_),
    .C(_04770_),
    .Y(_04773_));
 sky130_fd_sc_hd__and2_1 _11633_ (.A(_04771_),
    .B(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__o21bai_1 _11634_ (.A1(_04588_),
    .A2(_04684_),
    .B1_N(_04685_),
    .Y(_04775_));
 sky130_fd_sc_hd__or2_1 _11635_ (.A(_04590_),
    .B(_04686_),
    .X(_04776_));
 sky130_fd_sc_hd__nor2_1 _11636_ (.A(_04592_),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__inv_2 _11637_ (.A(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(_04394_),
    .B(_04777_),
    .Y(_04779_));
 sky130_fd_sc_hd__o211a_1 _11639_ (.A1(_04591_),
    .A2(_04776_),
    .B1(_04779_),
    .C1(_04775_),
    .X(_04780_));
 sky130_fd_sc_hd__o31a_1 _11640_ (.A1(_03974_),
    .A2(_04395_),
    .A3(_04778_),
    .B1(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__xnor2_1 _11641_ (.A(_04774_),
    .B(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__o21ai_1 _11642_ (.A1(_04727_),
    .A2(_04782_),
    .B1(net202),
    .Y(_04783_));
 sky130_fd_sc_hd__a21o_2 _11643_ (.A1(_04727_),
    .A2(_04782_),
    .B1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__a21oi_1 _11644_ (.A1(net155),
    .A2(_02199_),
    .B1(_02200_),
    .Y(_04785_));
 sky130_fd_sc_hd__a31o_1 _11645_ (.A1(net155),
    .A2(_02199_),
    .A3(_02200_),
    .B1(_02318_),
    .X(_04786_));
 sky130_fd_sc_hd__a21o_1 _11646_ (.A1(_05836_),
    .A2(_04698_),
    .B1(_05810_),
    .X(_04787_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(_06372_),
    .A1(_04787_),
    .S(_04563_),
    .X(_04788_));
 sky130_fd_sc_hd__o21ai_1 _11648_ (.A1(_05709_),
    .A2(_04788_),
    .B1(net242),
    .Y(_04789_));
 sky130_fd_sc_hd__a21o_1 _11649_ (.A1(_05709_),
    .A2(_04788_),
    .B1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__nand2_1 _11650_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .Y(_04791_));
 sky130_fd_sc_hd__or2_1 _11651_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .X(_04792_));
 sky130_fd_sc_hd__nand2_1 _11652_ (.A(_04791_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__o21ai_1 _11653_ (.A1(_04705_),
    .A2(_04706_),
    .B1(_04703_),
    .Y(_04794_));
 sky130_fd_sc_hd__xnor2_1 _11654_ (.A(_04793_),
    .B(_04794_),
    .Y(_04796_));
 sky130_fd_sc_hd__nor2_1 _11655_ (.A(_06300_),
    .B(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__a211o_1 _11656_ (.A1(_06300_),
    .A2(_03886_),
    .B1(_04797_),
    .C1(_06447_),
    .X(_04798_));
 sky130_fd_sc_hd__or2_1 _11657_ (.A(\div_res[19] ),
    .B(_04712_),
    .X(_04799_));
 sky130_fd_sc_hd__a21oi_1 _11658_ (.A1(net154),
    .A2(_04799_),
    .B1(\div_res[20] ),
    .Y(_04800_));
 sky130_fd_sc_hd__a31o_1 _11659_ (.A1(\div_res[20] ),
    .A2(net156),
    .A3(_04799_),
    .B1(net199),
    .X(_04801_));
 sky130_fd_sc_hd__a21o_1 _11660_ (.A1(_05690_),
    .A2(net240),
    .B1(net273),
    .X(_04802_));
 sky130_fd_sc_hd__o21ai_1 _11661_ (.A1(reg1_val[20]),
    .A2(_05681_),
    .B1(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__o221a_1 _11662_ (.A1(_05690_),
    .A2(net200),
    .B1(net236),
    .B2(reg1_val[20]),
    .C1(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__o221a_1 _11663_ (.A1(_02247_),
    .A2(_03873_),
    .B1(_03886_),
    .B2(_02316_),
    .C1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__or2_1 _11664_ (.A(\div_shifter[51] ),
    .B(_04709_),
    .X(_04807_));
 sky130_fd_sc_hd__a21oi_1 _11665_ (.A1(net232),
    .A2(_04807_),
    .B1(\div_shifter[52] ),
    .Y(_04808_));
 sky130_fd_sc_hd__a311o_1 _11666_ (.A1(\div_shifter[52] ),
    .A2(net232),
    .A3(_04807_),
    .B1(_04808_),
    .C1(net238),
    .X(_04809_));
 sky130_fd_sc_hd__o21a_1 _11667_ (.A1(_04800_),
    .A2(_04801_),
    .B1(_04805_),
    .X(_04810_));
 sky130_fd_sc_hd__and4_1 _11668_ (.A(_04790_),
    .B(_04798_),
    .C(_04809_),
    .D(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__o211a_1 _11669_ (.A1(_04785_),
    .A2(_04786_),
    .B1(_04811_),
    .C1(_04784_),
    .X(_04812_));
 sky130_fd_sc_hd__o22a_1 _11670_ (.A1(_05671_),
    .A2(net251),
    .B1(_06457_),
    .B2(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__and3_1 _11671_ (.A(curr_PC[19]),
    .B(curr_PC[20]),
    .C(_04628_),
    .X(_04814_));
 sky130_fd_sc_hd__a21oi_1 _11672_ (.A1(curr_PC[19]),
    .A2(_04628_),
    .B1(curr_PC[20]),
    .Y(_04815_));
 sky130_fd_sc_hd__or3_2 _11673_ (.A(net254),
    .B(_04814_),
    .C(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__o21ai_4 _11674_ (.A1(net259),
    .A2(_04813_),
    .B1(_04816_),
    .Y(dest_val[20]));
 sky130_fd_sc_hd__o22a_1 _11675_ (.A1(net63),
    .A2(net15),
    .B1(net6),
    .B2(net78),
    .X(_04818_));
 sky130_fd_sc_hd__xnor2_1 _11676_ (.A(net41),
    .B(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__o22a_1 _11677_ (.A1(net37),
    .A2(net21),
    .B1(net60),
    .B2(net35),
    .X(_04820_));
 sky130_fd_sc_hd__xnor2_1 _11678_ (.A(net120),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(_04819_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__or2_1 _11680_ (.A(_04819_),
    .B(_04821_),
    .X(_04823_));
 sky130_fd_sc_hd__and2_1 _11681_ (.A(_04822_),
    .B(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__o22a_1 _11682_ (.A1(net25),
    .A2(net64),
    .B1(net59),
    .B2(net28),
    .X(_04825_));
 sky130_fd_sc_hd__xnor2_1 _11683_ (.A(net66),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__inv_2 _11684_ (.A(_04826_),
    .Y(_04828_));
 sky130_fd_sc_hd__nand2_1 _11685_ (.A(_04824_),
    .B(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__or2_1 _11686_ (.A(_04824_),
    .B(_04828_),
    .X(_04830_));
 sky130_fd_sc_hd__nand2_1 _11687_ (.A(_04829_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__or3b_1 _11688_ (.A(net71),
    .B(net39),
    .C_N(_04748_),
    .X(_04832_));
 sky130_fd_sc_hd__or2_1 _11689_ (.A(_04831_),
    .B(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__nand2_1 _11690_ (.A(_04831_),
    .B(_04832_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand2_1 _11691_ (.A(_04833_),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__o22a_1 _11692_ (.A1(net29),
    .A2(net23),
    .B1(net19),
    .B2(net32),
    .X(_04836_));
 sky130_fd_sc_hd__xnor2_1 _11693_ (.A(net116),
    .B(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__and2_1 _11694_ (.A(net110),
    .B(_04837_),
    .X(_04839_));
 sky130_fd_sc_hd__xnor2_1 _11695_ (.A(net110),
    .B(_04837_),
    .Y(_04840_));
 sky130_fd_sc_hd__o22a_1 _11696_ (.A1(net33),
    .A2(net17),
    .B1(net8),
    .B2(net79),
    .X(_04841_));
 sky130_fd_sc_hd__xnor2_1 _11697_ (.A(net113),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__and2b_1 _11698_ (.A_N(_04840_),
    .B(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__and2b_1 _11699_ (.A_N(_04842_),
    .B(_04840_),
    .X(_04844_));
 sky130_fd_sc_hd__or2_1 _11700_ (.A(_04843_),
    .B(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__xnor2_1 _11701_ (.A(_04835_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__o21ai_1 _11702_ (.A1(_04739_),
    .A2(_04753_),
    .B1(_04751_),
    .Y(_04847_));
 sky130_fd_sc_hd__a21bo_1 _11703_ (.A1(_04756_),
    .A2(_04758_),
    .B1_N(_04757_),
    .X(_04848_));
 sky130_fd_sc_hd__nor2_1 _11704_ (.A(net74),
    .B(net39),
    .Y(_04850_));
 sky130_fd_sc_hd__o21a_1 _11705_ (.A1(_04733_),
    .A2(_04737_),
    .B1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__or3_1 _11706_ (.A(_04733_),
    .B(_04737_),
    .C(_04850_),
    .X(_04852_));
 sky130_fd_sc_hd__nand2b_1 _11707_ (.A_N(_04851_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__nor2_1 _11708_ (.A(_04745_),
    .B(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__and2_1 _11709_ (.A(_04745_),
    .B(_04853_),
    .X(_04855_));
 sky130_fd_sc_hd__or2_1 _11710_ (.A(_04854_),
    .B(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__and2b_1 _11711_ (.A_N(_04856_),
    .B(_04848_),
    .X(_04857_));
 sky130_fd_sc_hd__xnor2_1 _11712_ (.A(_04848_),
    .B(_04856_),
    .Y(_04858_));
 sky130_fd_sc_hd__xnor2_1 _11713_ (.A(_04847_),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__or2_1 _11714_ (.A(_04846_),
    .B(_04859_),
    .X(_04861_));
 sky130_fd_sc_hd__nand2_1 _11715_ (.A(_04846_),
    .B(_04859_),
    .Y(_04862_));
 sky130_fd_sc_hd__and2_1 _11716_ (.A(_04861_),
    .B(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__o21ba_1 _11717_ (.A1(_04760_),
    .A2(_04761_),
    .B1_N(_04763_),
    .X(_04864_));
 sky130_fd_sc_hd__nand2b_1 _11718_ (.A_N(_04864_),
    .B(_04863_),
    .Y(_04865_));
 sky130_fd_sc_hd__xnor2_1 _11719_ (.A(_04863_),
    .B(_04864_),
    .Y(_04866_));
 sky130_fd_sc_hd__o21ai_2 _11720_ (.A1(_04766_),
    .A2(_04769_),
    .B1(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__inv_2 _11721_ (.A(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__nor3_1 _11722_ (.A(_04766_),
    .B(_04769_),
    .C(_04866_),
    .Y(_04869_));
 sky130_fd_sc_hd__nor2_2 _11723_ (.A(_04868_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__nand2b_1 _11724_ (.A_N(_04686_),
    .B(_04774_),
    .Y(_04872_));
 sky130_fd_sc_hd__inv_2 _11725_ (.A(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__o21ai_1 _11726_ (.A1(_04684_),
    .A2(_04772_),
    .B1(_04773_),
    .Y(_04874_));
 sky130_fd_sc_hd__a21bo_1 _11727_ (.A1(_04687_),
    .A2(_04873_),
    .B1_N(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__a31o_1 _11728_ (.A1(_04500_),
    .A2(_04688_),
    .A3(_04873_),
    .B1(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__xnor2_2 _11729_ (.A(_04870_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__or4_1 _11730_ (.A(_04435_),
    .B(_04501_),
    .C(_04725_),
    .D(_04782_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _11731_ (.A(net157),
    .B(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__a21oi_1 _11732_ (.A1(_04877_),
    .A2(_04879_),
    .B1(_02242_),
    .Y(_04880_));
 sky130_fd_sc_hd__o21ai_2 _11733_ (.A1(_04877_),
    .A2(_04879_),
    .B1(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__a21oi_1 _11734_ (.A1(net156),
    .A2(_02201_),
    .B1(_02204_),
    .Y(_04883_));
 sky130_fd_sc_hd__a311o_1 _11735_ (.A1(net155),
    .A2(_02201_),
    .A3(_02204_),
    .B1(_02318_),
    .C1(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__o21a_1 _11736_ (.A1(_05709_),
    .A2(_06372_),
    .B1(_06375_),
    .X(_04885_));
 sky130_fd_sc_hd__a21bo_1 _11737_ (.A1(_05709_),
    .A2(_04787_),
    .B1_N(_05690_),
    .X(_04886_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(_04885_),
    .A1(_04886_),
    .S(net297),
    .X(_04887_));
 sky130_fd_sc_hd__nor2_1 _11739_ (.A(_05764_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__a21o_1 _11740_ (.A1(_05764_),
    .A2(_04887_),
    .B1(net241),
    .X(_04889_));
 sky130_fd_sc_hd__nand2_1 _11741_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_04890_));
 sky130_fd_sc_hd__or2_1 _11742_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_1 _11743_ (.A(_04890_),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21bo_1 _11744_ (.A1(_04792_),
    .A2(_04794_),
    .B1_N(_04791_),
    .X(_04894_));
 sky130_fd_sc_hd__xnor2_1 _11745_ (.A(_04892_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__nor2_1 _11746_ (.A(_06300_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__a211o_1 _11747_ (.A1(_06300_),
    .A2(_03764_),
    .B1(_04896_),
    .C1(net209),
    .X(_04897_));
 sky130_fd_sc_hd__or2_1 _11748_ (.A(\div_shifter[52] ),
    .B(_04807_),
    .X(_04898_));
 sky130_fd_sc_hd__a21oi_1 _11749_ (.A1(net232),
    .A2(_04898_),
    .B1(\div_shifter[53] ),
    .Y(_04899_));
 sky130_fd_sc_hd__a31o_1 _11750_ (.A1(\div_shifter[53] ),
    .A2(net232),
    .A3(_04898_),
    .B1(net238),
    .X(_04900_));
 sky130_fd_sc_hd__or3_1 _11751_ (.A(\div_res[20] ),
    .B(\div_res[19] ),
    .C(_04712_),
    .X(_04901_));
 sky130_fd_sc_hd__a21oi_1 _11752_ (.A1(net154),
    .A2(_04901_),
    .B1(\div_res[21] ),
    .Y(_04902_));
 sky130_fd_sc_hd__a31o_1 _11753_ (.A1(\div_res[21] ),
    .A2(net154),
    .A3(_04901_),
    .B1(net199),
    .X(_04903_));
 sky130_fd_sc_hd__or2_1 _11754_ (.A(_04902_),
    .B(_04903_),
    .X(_04905_));
 sky130_fd_sc_hd__o21a_1 _11755_ (.A1(_05747_),
    .A2(_02327_),
    .B1(_02323_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_1 _11756_ (.A(_05747_),
    .B(net201),
    .Y(_04907_));
 sky130_fd_sc_hd__o221a_1 _11757_ (.A1(reg1_val[21]),
    .A2(net236),
    .B1(_04906_),
    .B2(_05755_),
    .C1(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__o221a_1 _11758_ (.A1(_02247_),
    .A2(_03751_),
    .B1(_03764_),
    .B2(_02316_),
    .C1(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__o211a_1 _11759_ (.A1(_04899_),
    .A2(_04900_),
    .B1(_04905_),
    .C1(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__o211a_1 _11760_ (.A1(_04888_),
    .A2(_04889_),
    .B1(_04897_),
    .C1(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__a31o_1 _11761_ (.A1(_04881_),
    .A2(_04884_),
    .A3(_04911_),
    .B1(_06457_),
    .X(_04912_));
 sky130_fd_sc_hd__o21a_1 _11762_ (.A1(_05737_),
    .A2(net251),
    .B1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__nor2_1 _11763_ (.A(curr_PC[21]),
    .B(_04814_),
    .Y(_04914_));
 sky130_fd_sc_hd__and2_1 _11764_ (.A(curr_PC[21]),
    .B(_04814_),
    .X(_04916_));
 sky130_fd_sc_hd__or3_2 _11765_ (.A(net254),
    .B(_04914_),
    .C(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__o21ai_4 _11766_ (.A1(net258),
    .A2(_04913_),
    .B1(_04917_),
    .Y(dest_val[21]));
 sky130_fd_sc_hd__and2b_1 _11767_ (.A_N(_04782_),
    .B(_04877_),
    .X(_04918_));
 sky130_fd_sc_hd__a21o_1 _11768_ (.A1(_04726_),
    .A2(_04918_),
    .B1(net149),
    .X(_04919_));
 sky130_fd_sc_hd__o22a_1 _11769_ (.A1(net28),
    .A2(net60),
    .B1(net59),
    .B2(net25),
    .X(_04920_));
 sky130_fd_sc_hd__xnor2_1 _11770_ (.A(net66),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__o22a_1 _11771_ (.A1(net37),
    .A2(net23),
    .B1(net21),
    .B2(net35),
    .X(_04922_));
 sky130_fd_sc_hd__xnor2_1 _11772_ (.A(net120),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2b_1 _11773_ (.A_N(_04921_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand2b_1 _11774_ (.A_N(_04923_),
    .B(_04921_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand2_1 _11775_ (.A(_04924_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__a21o_1 _11776_ (.A1(_04822_),
    .A2(_04829_),
    .B1(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__nand3_1 _11777_ (.A(_04822_),
    .B(_04829_),
    .C(_04927_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _11778_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__o22a_1 _11779_ (.A1(net29),
    .A2(net20),
    .B1(net18),
    .B2(net32),
    .X(_04931_));
 sky130_fd_sc_hd__xnor2_1 _11780_ (.A(net117),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__o31a_1 _11781_ (.A1(net111),
    .A2(_06507_),
    .A3(net9),
    .B1(net114),
    .X(_04933_));
 sky130_fd_sc_hd__nor2_1 _11782_ (.A(_06515_),
    .B(net8),
    .Y(_04934_));
 sky130_fd_sc_hd__nor3_2 _11783_ (.A(_04932_),
    .B(_04933_),
    .C(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__o21a_1 _11784_ (.A1(_04933_),
    .A2(_04934_),
    .B1(_04932_),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_2 _11785_ (.A(_04935_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__xor2_1 _11786_ (.A(_04930_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__o21a_1 _11787_ (.A1(_04835_),
    .A2(_04845_),
    .B1(_04833_),
    .X(_04940_));
 sky130_fd_sc_hd__o22a_1 _11788_ (.A1(net64),
    .A2(net15),
    .B1(net6),
    .B2(net63),
    .X(_04941_));
 sky130_fd_sc_hd__xnor2_1 _11789_ (.A(net41),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__o21ai_1 _11790_ (.A1(_04839_),
    .A2(_04843_),
    .B1(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__or3_1 _11791_ (.A(_04839_),
    .B(_04843_),
    .C(_04942_),
    .X(_04944_));
 sky130_fd_sc_hd__and2_1 _11792_ (.A(_04943_),
    .B(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_00186_),
    .B(net42),
    .Y(_04946_));
 sky130_fd_sc_hd__or3b_1 _11794_ (.A(net78),
    .B(net39),
    .C_N(_04945_),
    .X(_04948_));
 sky130_fd_sc_hd__xnor2_1 _11795_ (.A(_04945_),
    .B(_04946_),
    .Y(_04949_));
 sky130_fd_sc_hd__o21ai_1 _11796_ (.A1(_04851_),
    .A2(_04854_),
    .B1(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__or3_1 _11797_ (.A(_04851_),
    .B(_04854_),
    .C(_04949_),
    .X(_04951_));
 sky130_fd_sc_hd__and2_1 _11798_ (.A(_04950_),
    .B(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__nand2b_1 _11799_ (.A_N(_04940_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__xnor2_1 _11800_ (.A(_04940_),
    .B(_04952_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _11801_ (.A(_04939_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__xnor2_1 _11802_ (.A(_04939_),
    .B(_04954_),
    .Y(_04956_));
 sky130_fd_sc_hd__a21oi_1 _11803_ (.A1(_04847_),
    .A2(_04858_),
    .B1(_04857_),
    .Y(_04957_));
 sky130_fd_sc_hd__or2_1 _11804_ (.A(_04956_),
    .B(_04957_),
    .X(_04959_));
 sky130_fd_sc_hd__nand2_1 _11805_ (.A(_04956_),
    .B(_04957_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_1 _11806_ (.A(_04959_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__a21o_1 _11807_ (.A1(_04861_),
    .A2(_04865_),
    .B1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__inv_2 _11808_ (.A(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__and3_1 _11809_ (.A(_04861_),
    .B(_04865_),
    .C(_04961_),
    .X(_04964_));
 sky130_fd_sc_hd__nor2_2 _11810_ (.A(_04963_),
    .B(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__a21o_1 _11811_ (.A1(_04771_),
    .A2(_04867_),
    .B1(_04869_),
    .X(_04966_));
 sky130_fd_sc_hd__nand2_1 _11812_ (.A(_04774_),
    .B(_04870_),
    .Y(_04967_));
 sky130_fd_sc_hd__o21ai_1 _11813_ (.A1(_04775_),
    .A2(_04967_),
    .B1(_04966_),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _11814_ (.A(_04776_),
    .B(_04967_),
    .Y(_04970_));
 sky130_fd_sc_hd__a21o_1 _11815_ (.A1(_04595_),
    .A2(_04970_),
    .B1(_04968_),
    .X(_04971_));
 sky130_fd_sc_hd__xnor2_2 _11816_ (.A(_04965_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__o21ai_1 _11817_ (.A1(_04919_),
    .A2(_04972_),
    .B1(net202),
    .Y(_04973_));
 sky130_fd_sc_hd__a21o_1 _11818_ (.A1(_04919_),
    .A2(_04972_),
    .B1(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__a21oi_1 _11819_ (.A1(net153),
    .A2(_02205_),
    .B1(_02206_),
    .Y(_04975_));
 sky130_fd_sc_hd__and3_1 _11820_ (.A(net153),
    .B(_02205_),
    .C(_02206_),
    .X(_04976_));
 sky130_fd_sc_hd__a21o_1 _11821_ (.A1(_05764_),
    .A2(_04886_),
    .B1(_05747_),
    .X(_04977_));
 sky130_fd_sc_hd__o21a_1 _11822_ (.A1(_05764_),
    .A2(_04885_),
    .B1(_06374_),
    .X(_04978_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(_04977_),
    .A1(_04978_),
    .S(net304),
    .X(_04979_));
 sky130_fd_sc_hd__nor2_1 _11824_ (.A(_05643_),
    .B(_04979_),
    .Y(_04981_));
 sky130_fd_sc_hd__a21o_1 _11825_ (.A1(_05643_),
    .A2(_04979_),
    .B1(_02325_),
    .X(_04982_));
 sky130_fd_sc_hd__nand2_1 _11826_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_04983_));
 sky130_fd_sc_hd__or2_1 _11827_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .X(_04984_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(_04983_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__a21boi_1 _11829_ (.A1(_04891_),
    .A2(_04894_),
    .B1_N(_04890_),
    .Y(_04986_));
 sky130_fd_sc_hd__xnor2_1 _11830_ (.A(_04985_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(_03641_),
    .A1(_04987_),
    .S(net261),
    .X(_04988_));
 sky130_fd_sc_hd__or2_1 _11832_ (.A(\div_shifter[53] ),
    .B(_04898_),
    .X(_04989_));
 sky130_fd_sc_hd__a21oi_1 _11833_ (.A1(net232),
    .A2(_04989_),
    .B1(\div_shifter[54] ),
    .Y(_04990_));
 sky130_fd_sc_hd__a311o_1 _11834_ (.A1(\div_shifter[54] ),
    .A2(net232),
    .A3(_04989_),
    .B1(_04990_),
    .C1(net238),
    .X(_04992_));
 sky130_fd_sc_hd__or2_1 _11835_ (.A(\div_res[21] ),
    .B(_04901_),
    .X(_04993_));
 sky130_fd_sc_hd__a21oi_1 _11836_ (.A1(net156),
    .A2(_04993_),
    .B1(\div_res[22] ),
    .Y(_04994_));
 sky130_fd_sc_hd__a31o_1 _11837_ (.A1(\div_res[22] ),
    .A2(net156),
    .A3(_04993_),
    .B1(net199),
    .X(_04995_));
 sky130_fd_sc_hd__a21oi_1 _11838_ (.A1(_05614_),
    .A2(net240),
    .B1(net273),
    .Y(_04996_));
 sky130_fd_sc_hd__o22a_1 _11839_ (.A1(_05595_),
    .A2(net252),
    .B1(net237),
    .B2(reg1_val[22]),
    .X(_04997_));
 sky130_fd_sc_hd__o221a_1 _11840_ (.A1(_05614_),
    .A2(net200),
    .B1(_04996_),
    .B2(_05633_),
    .C1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__o221a_1 _11841_ (.A1(_02247_),
    .A2(_03630_),
    .B1(_03641_),
    .B2(_02316_),
    .C1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__o211a_1 _11842_ (.A1(_04994_),
    .A2(_04995_),
    .B1(_04999_),
    .C1(_04992_),
    .X(_05000_));
 sky130_fd_sc_hd__o221a_1 _11843_ (.A1(_04981_),
    .A2(_04982_),
    .B1(_04988_),
    .B2(net209),
    .C1(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__o311a_1 _11844_ (.A1(_02318_),
    .A2(_04975_),
    .A3(_04976_),
    .B1(_05001_),
    .C1(_04974_),
    .X(_05003_));
 sky130_fd_sc_hd__a21oi_1 _11845_ (.A1(curr_PC[22]),
    .A2(_04916_),
    .B1(net254),
    .Y(_05004_));
 sky130_fd_sc_hd__o21ai_2 _11846_ (.A1(curr_PC[22]),
    .A2(_04916_),
    .B1(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__o21ai_4 _11847_ (.A1(net258),
    .A2(_05003_),
    .B1(_05005_),
    .Y(dest_val[22]));
 sky130_fd_sc_hd__a31o_1 _11848_ (.A1(_04726_),
    .A2(_04918_),
    .A3(_04972_),
    .B1(net149),
    .X(_05006_));
 sky130_fd_sc_hd__nand2_1 _11849_ (.A(_04950_),
    .B(_04953_),
    .Y(_05007_));
 sky130_fd_sc_hd__o22a_1 _11850_ (.A1(net35),
    .A2(net23),
    .B1(net19),
    .B2(net37),
    .X(_05008_));
 sky130_fd_sc_hd__xnor2_1 _11851_ (.A(_06472_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__nor2_1 _11852_ (.A(net113),
    .B(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__and2_1 _11853_ (.A(net113),
    .B(_05009_),
    .X(_05011_));
 sky130_fd_sc_hd__or2_1 _11854_ (.A(_05010_),
    .B(_05011_),
    .X(_05013_));
 sky130_fd_sc_hd__o22a_1 _11855_ (.A1(net29),
    .A2(net17),
    .B1(net8),
    .B2(net32),
    .X(_05014_));
 sky130_fd_sc_hd__xor2_1 _11856_ (.A(net116),
    .B(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__nor2_1 _11857_ (.A(_05013_),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__and2_1 _11858_ (.A(_05013_),
    .B(_05015_),
    .X(_05017_));
 sky130_fd_sc_hd__or2_1 _11859_ (.A(_05016_),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__nor2_1 _11860_ (.A(_04935_),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__and2_1 _11861_ (.A(_04935_),
    .B(_05018_),
    .X(_05020_));
 sky130_fd_sc_hd__nor2_1 _11862_ (.A(_05019_),
    .B(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__and2b_1 _11863_ (.A_N(_04924_),
    .B(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__xnor2_1 _11864_ (.A(_04924_),
    .B(_05021_),
    .Y(_05024_));
 sky130_fd_sc_hd__o21ai_1 _11865_ (.A1(_04930_),
    .A2(_04938_),
    .B1(_04928_),
    .Y(_05025_));
 sky130_fd_sc_hd__o22a_1 _11866_ (.A1(net59),
    .A2(net15),
    .B1(net6),
    .B2(net64),
    .X(_05026_));
 sky130_fd_sc_hd__xnor2_1 _11867_ (.A(net41),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__or2_1 _11868_ (.A(net63),
    .B(net39),
    .X(_05028_));
 sky130_fd_sc_hd__o22a_1 _11869_ (.A1(net27),
    .A2(net21),
    .B1(net60),
    .B2(net25),
    .X(_05029_));
 sky130_fd_sc_hd__xnor2_1 _11870_ (.A(net66),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__nor2_1 _11871_ (.A(_05028_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__and2_1 _11872_ (.A(_05028_),
    .B(_05030_),
    .X(_05032_));
 sky130_fd_sc_hd__nor2_1 _11873_ (.A(_05031_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__and2_1 _11874_ (.A(_05027_),
    .B(_05033_),
    .X(_05035_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(_05027_),
    .B(_05033_),
    .Y(_05036_));
 sky130_fd_sc_hd__or2_1 _11876_ (.A(_05035_),
    .B(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__a21oi_1 _11877_ (.A1(_04943_),
    .A2(_04948_),
    .B1(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__and3_1 _11878_ (.A(_04943_),
    .B(_04948_),
    .C(_05037_),
    .X(_05039_));
 sky130_fd_sc_hd__or2_1 _11879_ (.A(_05038_),
    .B(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__and2b_1 _11880_ (.A_N(_05040_),
    .B(_05025_),
    .X(_05041_));
 sky130_fd_sc_hd__xnor2_1 _11881_ (.A(_05025_),
    .B(_05040_),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _11882_ (.A(_05024_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__or2_1 _11883_ (.A(_05024_),
    .B(_05042_),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_1 _11884_ (.A(_05043_),
    .B(_05044_),
    .Y(_05046_));
 sky130_fd_sc_hd__nand2b_1 _11885_ (.A_N(_05046_),
    .B(_05007_),
    .Y(_05047_));
 sky130_fd_sc_hd__xor2_1 _11886_ (.A(_05007_),
    .B(_05046_),
    .X(_05048_));
 sky130_fd_sc_hd__a21o_1 _11887_ (.A1(_04955_),
    .A2(_04959_),
    .B1(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__and3_1 _11888_ (.A(_04955_),
    .B(_04959_),
    .C(_05048_),
    .X(_05050_));
 sky130_fd_sc_hd__inv_2 _11889_ (.A(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand2_2 _11890_ (.A(_05049_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__inv_2 _11891_ (.A(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__nand2_1 _11892_ (.A(_04870_),
    .B(_04965_),
    .Y(_05054_));
 sky130_fd_sc_hd__nor2_1 _11893_ (.A(_04872_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__nor2_1 _11894_ (.A(_04874_),
    .B(_05054_),
    .Y(_05057_));
 sky130_fd_sc_hd__a21oi_1 _11895_ (.A1(_04867_),
    .A2(_04962_),
    .B1(_04964_),
    .Y(_05058_));
 sky130_fd_sc_hd__a211o_1 _11896_ (.A1(_04689_),
    .A2(_05055_),
    .B1(_05057_),
    .C1(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__a31oi_4 _11897_ (.A1(_04295_),
    .A2(_04690_),
    .A3(_05055_),
    .B1(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__xnor2_2 _11898_ (.A(_05052_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21ai_1 _11899_ (.A1(_05006_),
    .A2(_05061_),
    .B1(net202),
    .Y(_05062_));
 sky130_fd_sc_hd__a21oi_2 _11900_ (.A1(_05006_),
    .A2(_05061_),
    .B1(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__o21ai_1 _11901_ (.A1(net150),
    .A2(_02207_),
    .B1(_02208_),
    .Y(_05064_));
 sky130_fd_sc_hd__o311a_1 _11902_ (.A1(net150),
    .A2(_02207_),
    .A3(_02208_),
    .B1(_02317_),
    .C1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__o211a_1 _11903_ (.A1(_05643_),
    .A2(_04978_),
    .B1(_06378_),
    .C1(net304),
    .X(_05066_));
 sky130_fd_sc_hd__a21o_1 _11904_ (.A1(_05643_),
    .A2(_04977_),
    .B1(_05623_),
    .X(_05068_));
 sky130_fd_sc_hd__a21o_1 _11905_ (.A1(net297),
    .A2(_05068_),
    .B1(_05066_),
    .X(_05069_));
 sky130_fd_sc_hd__nand2_1 _11906_ (.A(_05565_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__o211a_1 _11907_ (.A1(_05565_),
    .A2(_05069_),
    .B1(_05070_),
    .C1(net242),
    .X(_05071_));
 sky130_fd_sc_hd__and2_1 _11908_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .X(_05072_));
 sky130_fd_sc_hd__nor2_1 _11909_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .Y(_05073_));
 sky130_fd_sc_hd__nor2_1 _11910_ (.A(_05072_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__o21a_1 _11911_ (.A1(_04985_),
    .A2(_04986_),
    .B1(_04983_),
    .X(_05075_));
 sky130_fd_sc_hd__xnor2_1 _11912_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__or2_1 _11913_ (.A(net260),
    .B(_03517_),
    .X(_05077_));
 sky130_fd_sc_hd__o211a_1 _11914_ (.A1(net229),
    .A2(_05076_),
    .B1(_05077_),
    .C1(net210),
    .X(_05079_));
 sky130_fd_sc_hd__o21a_1 _11915_ (.A1(\div_shifter[54] ),
    .A2(_04989_),
    .B1(net232),
    .X(_05080_));
 sky130_fd_sc_hd__o21ai_1 _11916_ (.A1(\div_shifter[55] ),
    .A2(_05080_),
    .B1(_02332_),
    .Y(_05081_));
 sky130_fd_sc_hd__a21oi_1 _11917_ (.A1(\div_shifter[55] ),
    .A2(_05080_),
    .B1(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__or2_1 _11918_ (.A(\div_res[22] ),
    .B(_04993_),
    .X(_05083_));
 sky130_fd_sc_hd__a21oi_1 _11919_ (.A1(net154),
    .A2(_05083_),
    .B1(\div_res[23] ),
    .Y(_05084_));
 sky130_fd_sc_hd__a311o_1 _11920_ (.A1(\div_res[23] ),
    .A2(net154),
    .A3(_05083_),
    .B1(_05084_),
    .C1(net199),
    .X(_05085_));
 sky130_fd_sc_hd__o21a_1 _11921_ (.A1(_05544_),
    .A2(_02327_),
    .B1(_02323_),
    .X(_05086_));
 sky130_fd_sc_hd__nand2_1 _11922_ (.A(_05544_),
    .B(net201),
    .Y(_05087_));
 sky130_fd_sc_hd__o221a_1 _11923_ (.A1(_05522_),
    .A2(net252),
    .B1(net237),
    .B2(reg1_val[23]),
    .C1(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__o21ai_1 _11924_ (.A1(_05554_),
    .A2(_05086_),
    .B1(_05088_),
    .Y(_05090_));
 sky130_fd_sc_hd__a221o_1 _11925_ (.A1(net246),
    .A2(_03510_),
    .B1(_03517_),
    .B2(_02315_),
    .C1(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__or4b_1 _11926_ (.A(_05079_),
    .B(_05082_),
    .C(_05091_),
    .D_N(_05085_),
    .X(_05092_));
 sky130_fd_sc_hd__o41a_1 _11927_ (.A1(_05063_),
    .A2(_05065_),
    .A3(_05071_),
    .A4(_05092_),
    .B1(net255),
    .X(_05093_));
 sky130_fd_sc_hd__a31o_1 _11928_ (.A1(curr_PC[21]),
    .A2(curr_PC[22]),
    .A3(_04814_),
    .B1(curr_PC[23]),
    .X(_05094_));
 sky130_fd_sc_hd__and3_2 _11929_ (.A(curr_PC[22]),
    .B(curr_PC[23]),
    .C(_04916_),
    .X(_05095_));
 sky130_fd_sc_hd__inv_2 _11930_ (.A(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__a31o_4 _11931_ (.A1(net258),
    .A2(_05094_),
    .A3(_05096_),
    .B1(_05093_),
    .X(dest_val[23]));
 sky130_fd_sc_hd__nor2_1 _11932_ (.A(_05038_),
    .B(_05041_),
    .Y(_05097_));
 sky130_fd_sc_hd__nand2_1 _11933_ (.A(_06526_),
    .B(net10),
    .Y(_05098_));
 sky130_fd_sc_hd__a2bb2o_2 _11934_ (.A1_N(_00137_),
    .A2_N(net8),
    .B1(_05098_),
    .B2(net117),
    .X(_05100_));
 sky130_fd_sc_hd__nor2_1 _11935_ (.A(net64),
    .B(net39),
    .Y(_05101_));
 sky130_fd_sc_hd__xnor2_1 _11936_ (.A(_05100_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__o21ai_1 _11937_ (.A1(_05010_),
    .A2(_05016_),
    .B1(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__or3_1 _11938_ (.A(_05010_),
    .B(_05016_),
    .C(_05102_),
    .X(_05104_));
 sky130_fd_sc_hd__and2_1 _11939_ (.A(_05103_),
    .B(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__o22a_1 _11940_ (.A1(net27),
    .A2(net23),
    .B1(net21),
    .B2(net25),
    .X(_05106_));
 sky130_fd_sc_hd__xnor2_1 _11941_ (.A(net66),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__o22a_1 _11942_ (.A1(net60),
    .A2(net15),
    .B1(net6),
    .B2(net59),
    .X(_05108_));
 sky130_fd_sc_hd__xnor2_1 _11943_ (.A(net41),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__o22a_1 _11944_ (.A1(net35),
    .A2(net19),
    .B1(net17),
    .B2(net37),
    .X(_05111_));
 sky130_fd_sc_hd__xnor2_1 _11945_ (.A(net120),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_05109_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__or2_1 _11947_ (.A(_05109_),
    .B(_05112_),
    .X(_05114_));
 sky130_fd_sc_hd__and2_1 _11948_ (.A(_05113_),
    .B(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__nand2b_1 _11949_ (.A_N(_05107_),
    .B(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__xnor2_1 _11950_ (.A(_05107_),
    .B(_05115_),
    .Y(_05117_));
 sky130_fd_sc_hd__o21ai_1 _11951_ (.A1(_05031_),
    .A2(_05035_),
    .B1(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__or3_1 _11952_ (.A(_05031_),
    .B(_05035_),
    .C(_05117_),
    .X(_05119_));
 sky130_fd_sc_hd__and2_1 _11953_ (.A(_05118_),
    .B(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__o21ai_1 _11954_ (.A1(_05019_),
    .A2(_05022_),
    .B1(_05120_),
    .Y(_05122_));
 sky130_fd_sc_hd__or3_1 _11955_ (.A(_05019_),
    .B(_05022_),
    .C(_05120_),
    .X(_05123_));
 sky130_fd_sc_hd__and2_1 _11956_ (.A(_05122_),
    .B(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__nand2_1 _11957_ (.A(_05105_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__or2_1 _11958_ (.A(_05105_),
    .B(_05124_),
    .X(_05126_));
 sky130_fd_sc_hd__nand2_1 _11959_ (.A(_05125_),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__or2_1 _11960_ (.A(_05097_),
    .B(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(_05097_),
    .B(_05127_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _11962_ (.A(_05128_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__a21o_1 _11963_ (.A1(_05043_),
    .A2(_05047_),
    .B1(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__nand3_1 _11964_ (.A(_05043_),
    .B(_05047_),
    .C(_05130_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand2_2 _11965_ (.A(_05131_),
    .B(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__a21oi_1 _11966_ (.A1(_04962_),
    .A2(_05049_),
    .B1(_05050_),
    .Y(_05135_));
 sky130_fd_sc_hd__nand2_1 _11967_ (.A(_04965_),
    .B(_05053_),
    .Y(_05136_));
 sky130_fd_sc_hd__o21bai_1 _11968_ (.A1(_04966_),
    .A2(_05136_),
    .B1_N(_05135_),
    .Y(_05137_));
 sky130_fd_sc_hd__or2_1 _11969_ (.A(_04967_),
    .B(_05136_),
    .X(_05138_));
 sky130_fd_sc_hd__o21ba_1 _11970_ (.A1(_04781_),
    .A2(_05138_),
    .B1_N(_05137_),
    .X(_05139_));
 sky130_fd_sc_hd__xnor2_2 _11971_ (.A(_05134_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__and4_2 _11972_ (.A(_04726_),
    .B(_04918_),
    .C(_04972_),
    .D(_05061_),
    .X(_05141_));
 sky130_fd_sc_hd__or2_1 _11973_ (.A(net149),
    .B(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__nand2_1 _11974_ (.A(_05140_),
    .B(_05142_),
    .Y(_05144_));
 sky130_fd_sc_hd__or2_1 _11975_ (.A(_05140_),
    .B(_05142_),
    .X(_05145_));
 sky130_fd_sc_hd__a21o_1 _11976_ (.A1(_02207_),
    .A2(_02208_),
    .B1(net150),
    .X(_05146_));
 sky130_fd_sc_hd__nand2_1 _11977_ (.A(_02209_),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__o211a_1 _11978_ (.A1(_02209_),
    .A2(_05146_),
    .B1(_05147_),
    .C1(_02317_),
    .X(_05148_));
 sky130_fd_sc_hd__a21oi_1 _11979_ (.A1(_05565_),
    .A2(_05068_),
    .B1(_05544_),
    .Y(_05149_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(_06380_),
    .A1(_05149_),
    .S(net298),
    .X(_05150_));
 sky130_fd_sc_hd__a21oi_1 _11981_ (.A1(_05186_),
    .A2(_05150_),
    .B1(net241),
    .Y(_05151_));
 sky130_fd_sc_hd__o21a_1 _11982_ (.A1(_05186_),
    .A2(_05150_),
    .B1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__o21ba_1 _11983_ (.A1(_05073_),
    .A2(_05075_),
    .B1_N(_05072_),
    .X(_05153_));
 sky130_fd_sc_hd__nor2_1 _11984_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05156_));
 sky130_fd_sc_hd__and2b_1 _11986_ (.A_N(_05155_),
    .B(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__xnor2_1 _11987_ (.A(_05153_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(_03370_),
    .A1(_05158_),
    .S(net260),
    .X(_05159_));
 sky130_fd_sc_hd__or3_1 _11989_ (.A(\div_shifter[55] ),
    .B(\div_shifter[54] ),
    .C(_04989_),
    .X(_05160_));
 sky130_fd_sc_hd__a21oi_1 _11990_ (.A1(net232),
    .A2(_05160_),
    .B1(\div_shifter[56] ),
    .Y(_05161_));
 sky130_fd_sc_hd__a311o_1 _11991_ (.A1(\div_shifter[56] ),
    .A2(net232),
    .A3(_05160_),
    .B1(_05161_),
    .C1(net238),
    .X(_05162_));
 sky130_fd_sc_hd__or2_1 _11992_ (.A(\div_res[23] ),
    .B(_05083_),
    .X(_05163_));
 sky130_fd_sc_hd__a21oi_1 _11993_ (.A1(net152),
    .A2(_05163_),
    .B1(\div_res[24] ),
    .Y(_05164_));
 sky130_fd_sc_hd__a31o_1 _11994_ (.A1(\div_res[24] ),
    .A2(net152),
    .A3(_05163_),
    .B1(net198),
    .X(_05166_));
 sky130_fd_sc_hd__nor2_1 _11995_ (.A(_05164_),
    .B(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__a21oi_1 _11996_ (.A1(_05165_),
    .A2(_02326_),
    .B1(net273),
    .Y(_05168_));
 sky130_fd_sc_hd__o22a_1 _11997_ (.A1(_05154_),
    .A2(net251),
    .B1(net237),
    .B2(reg1_val[24]),
    .X(_05169_));
 sky130_fd_sc_hd__o221ai_4 _11998_ (.A1(_05165_),
    .A2(net200),
    .B1(_05168_),
    .B2(_05176_),
    .C1(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__a221o_1 _11999_ (.A1(_02315_),
    .A2(_03370_),
    .B1(_03376_),
    .B2(net244),
    .C1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__or3b_1 _12000_ (.A(_05171_),
    .B(_05167_),
    .C_N(_05162_),
    .X(_05172_));
 sky130_fd_sc_hd__a211o_1 _12001_ (.A1(net210),
    .A2(_05159_),
    .B1(_05172_),
    .C1(_05152_),
    .X(_05173_));
 sky130_fd_sc_hd__a311o_1 _12002_ (.A1(net202),
    .A2(_05144_),
    .A3(_05145_),
    .B1(_05148_),
    .C1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__or2_1 _12003_ (.A(curr_PC[24]),
    .B(_05095_),
    .X(_05175_));
 sky130_fd_sc_hd__and2_1 _12004_ (.A(curr_PC[24]),
    .B(_05095_),
    .X(_05177_));
 sky130_fd_sc_hd__nor2_1 _12005_ (.A(net253),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a22o_4 _12006_ (.A1(net253),
    .A2(_05174_),
    .B1(_05175_),
    .B2(_05178_),
    .X(dest_val[24]));
 sky130_fd_sc_hd__a21o_1 _12007_ (.A1(_05140_),
    .A2(_05141_),
    .B1(net149),
    .X(_05179_));
 sky130_fd_sc_hd__o22a_1 _12008_ (.A1(net21),
    .A2(net15),
    .B1(net6),
    .B2(net60),
    .X(_05180_));
 sky130_fd_sc_hd__xnor2_1 _12009_ (.A(net41),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _12010_ (.A(_05100_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__or2_1 _12011_ (.A(_05100_),
    .B(_05181_),
    .X(_05183_));
 sky130_fd_sc_hd__nand2_1 _12012_ (.A(_05182_),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__or2_1 _12013_ (.A(net59),
    .B(net39),
    .X(_05185_));
 sky130_fd_sc_hd__xor2_1 _12014_ (.A(_05184_),
    .B(_05185_),
    .X(_05187_));
 sky130_fd_sc_hd__o31ai_2 _12015_ (.A1(net64),
    .A2(net39),
    .A3(_05100_),
    .B1(_05103_),
    .Y(_05188_));
 sky130_fd_sc_hd__o22a_1 _12016_ (.A1(net25),
    .A2(net23),
    .B1(net19),
    .B2(net27),
    .X(_05189_));
 sky130_fd_sc_hd__xnor2_1 _12017_ (.A(net66),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_1 _12018_ (.A(net116),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__and2_1 _12019_ (.A(net116),
    .B(_05190_),
    .X(_05192_));
 sky130_fd_sc_hd__nor2_1 _12020_ (.A(_05191_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__o22a_1 _12021_ (.A1(net35),
    .A2(net17),
    .B1(net8),
    .B2(net37),
    .X(_05194_));
 sky130_fd_sc_hd__xnor2_1 _12022_ (.A(net120),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__xnor2_1 _12023_ (.A(_05193_),
    .B(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_1 _12024_ (.A1(_05113_),
    .A2(_05116_),
    .B1(_05196_),
    .Y(_05198_));
 sky130_fd_sc_hd__and3_1 _12025_ (.A(_05113_),
    .B(_05116_),
    .C(_05196_),
    .X(_05199_));
 sky130_fd_sc_hd__nor2_1 _12026_ (.A(_05198_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__xor2_1 _12027_ (.A(_05188_),
    .B(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__nand2_1 _12028_ (.A(_05187_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__or2_1 _12029_ (.A(_05187_),
    .B(_05201_),
    .X(_05203_));
 sky130_fd_sc_hd__nand2_1 _12030_ (.A(_05202_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__a21o_1 _12031_ (.A1(_05118_),
    .A2(_05122_),
    .B1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__nand3_1 _12032_ (.A(_05118_),
    .B(_05122_),
    .C(_05204_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05205_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21o_1 _12034_ (.A1(_05125_),
    .A2(_05128_),
    .B1(_05207_),
    .X(_05209_));
 sky130_fd_sc_hd__inv_2 _12035_ (.A(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__and3_1 _12036_ (.A(_05125_),
    .B(_05128_),
    .C(_05207_),
    .X(_05211_));
 sky130_fd_sc_hd__nor2_1 _12037_ (.A(_05210_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__a21bo_1 _12038_ (.A1(_05049_),
    .A2(_05131_),
    .B1_N(_05133_),
    .X(_05213_));
 sky130_fd_sc_hd__o31a_1 _12039_ (.A1(_05052_),
    .A2(_05060_),
    .A3(_05134_),
    .B1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__xor2_2 _12040_ (.A(_05212_),
    .B(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__o21ai_1 _12041_ (.A1(_05179_),
    .A2(_05215_),
    .B1(net202),
    .Y(_05216_));
 sky130_fd_sc_hd__a21o_1 _12042_ (.A1(_05179_),
    .A2(_05215_),
    .B1(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__o21a_1 _12043_ (.A1(_05186_),
    .A2(_05149_),
    .B1(_05165_),
    .X(_05218_));
 sky130_fd_sc_hd__mux2_1 _12044_ (.A0(_06398_),
    .A1(_05218_),
    .S(net298),
    .X(_05220_));
 sky130_fd_sc_hd__nor2_1 _12045_ (.A(_05121_),
    .B(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__a211o_1 _12046_ (.A1(_05121_),
    .A2(_05220_),
    .B1(_05221_),
    .C1(net241),
    .X(_05222_));
 sky130_fd_sc_hd__a21oi_1 _12047_ (.A1(net153),
    .A2(_02210_),
    .B1(_02164_),
    .Y(_05223_));
 sky130_fd_sc_hd__a311o_1 _12048_ (.A1(net153),
    .A2(_02164_),
    .A3(_02210_),
    .B1(_02318_),
    .C1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__o21a_1 _12049_ (.A1(_05153_),
    .A2(_05155_),
    .B1(_05156_),
    .X(_05225_));
 sky130_fd_sc_hd__nor2_1 _12050_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_1 _12051_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05227_));
 sky130_fd_sc_hd__and2b_1 _12052_ (.A_N(_05226_),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__or2_1 _12053_ (.A(_05225_),
    .B(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__a21oi_1 _12054_ (.A1(_05225_),
    .A2(_05228_),
    .B1(net229),
    .Y(_05231_));
 sky130_fd_sc_hd__a22o_1 _12055_ (.A1(net229),
    .A2(_03237_),
    .B1(_05229_),
    .B2(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__or2_1 _12056_ (.A(\div_shifter[56] ),
    .B(_05160_),
    .X(_05233_));
 sky130_fd_sc_hd__a21oi_1 _12057_ (.A1(net232),
    .A2(_05233_),
    .B1(\div_shifter[57] ),
    .Y(_05234_));
 sky130_fd_sc_hd__a311o_1 _12058_ (.A1(\div_shifter[57] ),
    .A2(net232),
    .A3(_05233_),
    .B1(_05234_),
    .C1(net238),
    .X(_05235_));
 sky130_fd_sc_hd__or2_1 _12059_ (.A(\div_res[24] ),
    .B(_05163_),
    .X(_05236_));
 sky130_fd_sc_hd__a21oi_1 _12060_ (.A1(net152),
    .A2(_05236_),
    .B1(\div_res[25] ),
    .Y(_05237_));
 sky130_fd_sc_hd__a31o_1 _12061_ (.A1(\div_res[25] ),
    .A2(net152),
    .A3(_05236_),
    .B1(net198),
    .X(_05238_));
 sky130_fd_sc_hd__a21oi_1 _12062_ (.A1(_05099_),
    .A2(_02326_),
    .B1(net273),
    .Y(_05239_));
 sky130_fd_sc_hd__o22a_1 _12063_ (.A1(_05089_),
    .A2(net251),
    .B1(net237),
    .B2(reg1_val[25]),
    .X(_05240_));
 sky130_fd_sc_hd__o221a_1 _12064_ (.A1(_05099_),
    .A2(net200),
    .B1(_05239_),
    .B2(_05110_),
    .C1(_05240_),
    .X(_05242_));
 sky130_fd_sc_hd__o221a_1 _12065_ (.A1(_02316_),
    .A2(_03237_),
    .B1(_03244_),
    .B2(_02247_),
    .C1(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__o211a_1 _12066_ (.A1(_05237_),
    .A2(_05238_),
    .B1(_05243_),
    .C1(_05235_),
    .X(_05244_));
 sky130_fd_sc_hd__o211a_1 _12067_ (.A1(net209),
    .A2(_05232_),
    .B1(_05244_),
    .C1(_05224_),
    .X(_05245_));
 sky130_fd_sc_hd__a31o_1 _12068_ (.A1(_05217_),
    .A2(_05222_),
    .A3(_05245_),
    .B1(net259),
    .X(_05246_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(curr_PC[25]),
    .B(_05177_),
    .Y(_05247_));
 sky130_fd_sc_hd__and3_1 _12070_ (.A(curr_PC[24]),
    .B(curr_PC[25]),
    .C(_05095_),
    .X(_05248_));
 sky130_fd_sc_hd__o31ai_4 _12071_ (.A1(net253),
    .A2(_05247_),
    .A3(_05248_),
    .B1(_05246_),
    .Y(dest_val[25]));
 sky130_fd_sc_hd__and2_1 _12072_ (.A(_05140_),
    .B(_05215_),
    .X(_05249_));
 sky130_fd_sc_hd__a21o_1 _12073_ (.A1(_05141_),
    .A2(_05249_),
    .B1(net149),
    .X(_05250_));
 sky130_fd_sc_hd__o21ai_1 _12074_ (.A1(_05184_),
    .A2(_05185_),
    .B1(_05182_),
    .Y(_05252_));
 sky130_fd_sc_hd__a21o_1 _12075_ (.A1(_05193_),
    .A2(_05195_),
    .B1(_05191_),
    .X(_05253_));
 sky130_fd_sc_hd__o22a_1 _12076_ (.A1(net25),
    .A2(net19),
    .B1(net17),
    .B2(net28),
    .X(_05254_));
 sky130_fd_sc_hd__xor2_1 _12077_ (.A(net66),
    .B(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__nand2_1 _12078_ (.A(_06485_),
    .B(net10),
    .Y(_05256_));
 sky130_fd_sc_hd__a22o_1 _12079_ (.A1(_06492_),
    .A2(net10),
    .B1(_05256_),
    .B2(net121),
    .X(_05257_));
 sky130_fd_sc_hd__or2_1 _12080_ (.A(_05255_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_05255_),
    .B(_05257_),
    .Y(_05259_));
 sky130_fd_sc_hd__nand2_1 _12082_ (.A(_05258_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__xnor2_1 _12083_ (.A(_05253_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__and2b_1 _12084_ (.A_N(_05261_),
    .B(_05252_),
    .X(_05263_));
 sky130_fd_sc_hd__xnor2_1 _12085_ (.A(_05252_),
    .B(_05261_),
    .Y(_05264_));
 sky130_fd_sc_hd__o22a_1 _12086_ (.A1(net23),
    .A2(net15),
    .B1(net6),
    .B2(net21),
    .X(_05265_));
 sky130_fd_sc_hd__nor2_1 _12087_ (.A(_00284_),
    .B(net39),
    .Y(_05266_));
 sky130_fd_sc_hd__xnor2_1 _12088_ (.A(_05265_),
    .B(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_05264_),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__or2_1 _12090_ (.A(_05264_),
    .B(_05267_),
    .X(_05269_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_05268_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__a21oi_1 _12092_ (.A1(_05188_),
    .A2(_05200_),
    .B1(_05198_),
    .Y(_05271_));
 sky130_fd_sc_hd__or2_1 _12093_ (.A(_05270_),
    .B(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__nand2_1 _12094_ (.A(_05270_),
    .B(_05271_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(_05272_),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__a21o_1 _12096_ (.A1(_05202_),
    .A2(_05205_),
    .B1(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__inv_2 _12097_ (.A(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__and3_1 _12098_ (.A(_05202_),
    .B(_05205_),
    .C(_05275_),
    .X(_05278_));
 sky130_fd_sc_hd__nor2_2 _12099_ (.A(_05277_),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__a21oi_1 _12100_ (.A1(_05131_),
    .A2(_05209_),
    .B1(_05211_),
    .Y(_05280_));
 sky130_fd_sc_hd__and3_1 _12101_ (.A(_05131_),
    .B(_05133_),
    .C(_05212_),
    .X(_05281_));
 sky130_fd_sc_hd__or3_1 _12102_ (.A(_05134_),
    .B(_05210_),
    .C(_05211_),
    .X(_05282_));
 sky130_fd_sc_hd__a21o_1 _12103_ (.A1(_05135_),
    .A2(_05281_),
    .B1(_05280_),
    .X(_05283_));
 sky130_fd_sc_hd__a41o_1 _12104_ (.A1(_04965_),
    .A2(_04971_),
    .A3(_05053_),
    .A4(_05281_),
    .B1(_05283_),
    .X(_05285_));
 sky130_fd_sc_hd__xnor2_2 _12105_ (.A(_05279_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__or2_1 _12106_ (.A(_05250_),
    .B(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _12107_ (.A(_05250_),
    .B(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__o21a_1 _12108_ (.A1(_05121_),
    .A2(_05218_),
    .B1(_05099_),
    .X(_05289_));
 sky130_fd_sc_hd__mux2_1 _12109_ (.A0(_06399_),
    .A1(_05289_),
    .S(net298),
    .X(_05290_));
 sky130_fd_sc_hd__a21oi_1 _12110_ (.A1(_05349_),
    .A2(_05290_),
    .B1(net241),
    .Y(_05291_));
 sky130_fd_sc_hd__o21a_1 _12111_ (.A1(_05349_),
    .A2(_05290_),
    .B1(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__o21a_1 _12112_ (.A1(_05225_),
    .A2(_05226_),
    .B1(_05227_),
    .X(_05293_));
 sky130_fd_sc_hd__nor2_1 _12113_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05294_));
 sky130_fd_sc_hd__or2_1 _12114_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .X(_05296_));
 sky130_fd_sc_hd__nand2_1 _12115_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05297_));
 sky130_fd_sc_hd__a21oi_1 _12116_ (.A1(_05296_),
    .A2(_05297_),
    .B1(_05293_),
    .Y(_05298_));
 sky130_fd_sc_hd__a31o_1 _12117_ (.A1(_05293_),
    .A2(_05296_),
    .A3(_05297_),
    .B1(net229),
    .X(_05299_));
 sky130_fd_sc_hd__o22a_1 _12118_ (.A1(net260),
    .A2(_03099_),
    .B1(_05298_),
    .B2(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__o21a_1 _12119_ (.A1(\div_shifter[57] ),
    .A2(_05233_),
    .B1(net232),
    .X(_05301_));
 sky130_fd_sc_hd__o21ai_1 _12120_ (.A1(\div_shifter[58] ),
    .A2(_05301_),
    .B1(_02332_),
    .Y(_05302_));
 sky130_fd_sc_hd__a21oi_1 _12121_ (.A1(\div_shifter[58] ),
    .A2(_05301_),
    .B1(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__or2_1 _12122_ (.A(\div_res[25] ),
    .B(_05236_),
    .X(_05304_));
 sky130_fd_sc_hd__a21o_1 _12123_ (.A1(net152),
    .A2(_05304_),
    .B1(\div_res[26] ),
    .X(_05305_));
 sky130_fd_sc_hd__nand3_1 _12124_ (.A(\div_res[26] ),
    .B(net152),
    .C(_05304_),
    .Y(_05307_));
 sky130_fd_sc_hd__a21o_1 _12125_ (.A1(_05317_),
    .A2(_02326_),
    .B1(net273),
    .X(_05308_));
 sky130_fd_sc_hd__a2bb2o_1 _12126_ (.A1_N(reg1_val[26]),
    .A2_N(net237),
    .B1(_05306_),
    .B2(_06455_),
    .X(_05309_));
 sky130_fd_sc_hd__a221o_1 _12127_ (.A1(_05327_),
    .A2(net201),
    .B1(_05308_),
    .B2(_05338_),
    .C1(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__a221o_1 _12128_ (.A1(_02315_),
    .A2(_03099_),
    .B1(_03105_),
    .B2(net246),
    .C1(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__a31o_1 _12129_ (.A1(_02330_),
    .A2(_05305_),
    .A3(_05307_),
    .B1(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__a211o_1 _12130_ (.A1(net210),
    .A2(_05300_),
    .B1(_05303_),
    .C1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__or2_1 _12131_ (.A(net150),
    .B(_02211_),
    .X(_05314_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(_02213_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__or2_1 _12133_ (.A(_02213_),
    .B(_05314_),
    .X(_05316_));
 sky130_fd_sc_hd__a31o_1 _12134_ (.A1(_02317_),
    .A2(_05315_),
    .A3(_05316_),
    .B1(_05313_),
    .X(_05318_));
 sky130_fd_sc_hd__a311o_1 _12135_ (.A1(net202),
    .A2(_05287_),
    .A3(_05288_),
    .B1(_05292_),
    .C1(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__nand2_1 _12136_ (.A(curr_PC[26]),
    .B(_05248_),
    .Y(_05320_));
 sky130_fd_sc_hd__o21a_1 _12137_ (.A1(curr_PC[26]),
    .A2(_05248_),
    .B1(net258),
    .X(_05321_));
 sky130_fd_sc_hd__a22o_4 _12138_ (.A1(net254),
    .A2(_05319_),
    .B1(_05320_),
    .B2(_05321_),
    .X(dest_val[26]));
 sky130_fd_sc_hd__xnor2_1 _12139_ (.A(curr_PC[27]),
    .B(_05320_),
    .Y(_05322_));
 sky130_fd_sc_hd__o22a_1 _12140_ (.A1(net19),
    .A2(net15),
    .B1(net6),
    .B2(net23),
    .X(_05323_));
 sky130_fd_sc_hd__xnor2_1 _12141_ (.A(net41),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nand2_1 _12142_ (.A(_06472_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__or2_1 _12143_ (.A(_06472_),
    .B(_05324_),
    .X(_05326_));
 sky130_fd_sc_hd__and2_1 _12144_ (.A(_05325_),
    .B(_05326_),
    .X(_05328_));
 sky130_fd_sc_hd__inv_2 _12145_ (.A(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__o22a_1 _12146_ (.A1(net25),
    .A2(net17),
    .B1(net8),
    .B2(net27),
    .X(_05330_));
 sky130_fd_sc_hd__xnor2_1 _12147_ (.A(net66),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__xor2_1 _12148_ (.A(_05328_),
    .B(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__a21o_1 _12149_ (.A1(_00284_),
    .A2(_05265_),
    .B1(_00271_),
    .X(_05333_));
 sky130_fd_sc_hd__or4b_1 _12150_ (.A(net21),
    .B(net60),
    .C(net39),
    .D_N(_05265_),
    .X(_05334_));
 sky130_fd_sc_hd__and3_1 _12151_ (.A(net41),
    .B(_05333_),
    .C(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__xor2_1 _12152_ (.A(_05258_),
    .B(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__and2b_1 _12153_ (.A_N(_05332_),
    .B(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__xnor2_1 _12154_ (.A(_05332_),
    .B(_05336_),
    .Y(_05339_));
 sky130_fd_sc_hd__a21o_1 _12155_ (.A1(_05253_),
    .A2(_05260_),
    .B1(_05263_),
    .X(_05340_));
 sky130_fd_sc_hd__and2_1 _12156_ (.A(_05339_),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__xnor2_1 _12157_ (.A(_05339_),
    .B(_05340_),
    .Y(_05342_));
 sky130_fd_sc_hd__a21o_1 _12158_ (.A1(_05268_),
    .A2(_05272_),
    .B1(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__inv_2 _12159_ (.A(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__and3_1 _12160_ (.A(_05268_),
    .B(_05272_),
    .C(_05342_),
    .X(_05345_));
 sky130_fd_sc_hd__nor2_1 _12161_ (.A(_05344_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__a21o_1 _12162_ (.A1(_05209_),
    .A2(_05276_),
    .B1(_05278_),
    .X(_05347_));
 sky130_fd_sc_hd__nand2_1 _12163_ (.A(_05212_),
    .B(_05279_),
    .Y(_05348_));
 sky130_fd_sc_hd__o21ai_1 _12164_ (.A1(_05214_),
    .A2(_05348_),
    .B1(_05347_),
    .Y(_05350_));
 sky130_fd_sc_hd__xnor2_1 _12165_ (.A(_05346_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__a31o_1 _12166_ (.A1(_05141_),
    .A2(_05249_),
    .A3(_05286_),
    .B1(net149),
    .X(_05352_));
 sky130_fd_sc_hd__a21oi_1 _12167_ (.A1(_05351_),
    .A2(_05352_),
    .B1(_02242_),
    .Y(_05353_));
 sky130_fd_sc_hd__o21a_1 _12168_ (.A1(_05351_),
    .A2(_05352_),
    .B1(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__o21a_1 _12169_ (.A1(_05349_),
    .A2(_05289_),
    .B1(_05317_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _12170_ (.A0(_06400_),
    .A1(_05355_),
    .S(net298),
    .X(_05356_));
 sky130_fd_sc_hd__a21oi_1 _12171_ (.A1(_05273_),
    .A2(_05356_),
    .B1(net241),
    .Y(_05357_));
 sky130_fd_sc_hd__o21a_1 _12172_ (.A1(_05273_),
    .A2(_05356_),
    .B1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__a21oi_1 _12173_ (.A1(_02211_),
    .A2(_02213_),
    .B1(net150),
    .Y(_05359_));
 sky130_fd_sc_hd__xor2_1 _12174_ (.A(_02220_),
    .B(_05359_),
    .X(_05361_));
 sky130_fd_sc_hd__o21a_1 _12175_ (.A1(_05293_),
    .A2(_05294_),
    .B1(_05297_),
    .X(_05362_));
 sky130_fd_sc_hd__nor2_1 _12176_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _12177_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05364_));
 sky130_fd_sc_hd__and2b_1 _12178_ (.A_N(_05363_),
    .B(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__nor2_1 _12179_ (.A(_05362_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__a21o_1 _12180_ (.A1(_05362_),
    .A2(_05365_),
    .B1(net229),
    .X(_05367_));
 sky130_fd_sc_hd__or2_1 _12181_ (.A(net260),
    .B(_02957_),
    .X(_05368_));
 sky130_fd_sc_hd__o211a_1 _12182_ (.A1(_05366_),
    .A2(_05367_),
    .B1(_05368_),
    .C1(net210),
    .X(_05369_));
 sky130_fd_sc_hd__or3_1 _12183_ (.A(\div_shifter[58] ),
    .B(\div_shifter[57] ),
    .C(_05233_),
    .X(_05370_));
 sky130_fd_sc_hd__a21oi_1 _12184_ (.A1(net233),
    .A2(_05370_),
    .B1(\div_shifter[59] ),
    .Y(_05372_));
 sky130_fd_sc_hd__a311o_1 _12185_ (.A1(\div_shifter[59] ),
    .A2(net233),
    .A3(_05370_),
    .B1(_05372_),
    .C1(net238),
    .X(_05373_));
 sky130_fd_sc_hd__or2_1 _12186_ (.A(\div_res[26] ),
    .B(_05304_),
    .X(_05374_));
 sky130_fd_sc_hd__a21oi_1 _12187_ (.A1(net154),
    .A2(_05374_),
    .B1(\div_res[27] ),
    .Y(_05375_));
 sky130_fd_sc_hd__a31o_1 _12188_ (.A1(\div_res[27] ),
    .A2(net155),
    .A3(_05374_),
    .B1(net198),
    .X(_05376_));
 sky130_fd_sc_hd__nor2_1 _12189_ (.A(_05375_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__a21oi_1 _12190_ (.A1(_05262_),
    .A2(_02326_),
    .B1(net273),
    .Y(_05378_));
 sky130_fd_sc_hd__o221a_1 _12191_ (.A1(_05230_),
    .A2(net251),
    .B1(net237),
    .B2(reg1_val[27]),
    .C1(net255),
    .X(_05379_));
 sky130_fd_sc_hd__o221ai_4 _12192_ (.A1(_05262_),
    .A2(net200),
    .B1(_05378_),
    .B2(_05251_),
    .C1(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__a221o_1 _12193_ (.A1(_02315_),
    .A2(_02957_),
    .B1(_02963_),
    .B2(net245),
    .C1(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__or3b_1 _12194_ (.A(_05381_),
    .B(_05377_),
    .C_N(_05373_),
    .X(_05383_));
 sky130_fd_sc_hd__a211o_1 _12195_ (.A1(_02317_),
    .A2(_05361_),
    .B1(_05369_),
    .C1(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__o32a_4 _12196_ (.A1(_05354_),
    .A2(_05358_),
    .A3(_05384_),
    .B1(_05322_),
    .B2(net255),
    .X(dest_val[27]));
 sky130_fd_sc_hd__a21boi_1 _12197_ (.A1(_05258_),
    .A2(_05335_),
    .B1_N(_05334_),
    .Y(_05385_));
 sky130_fd_sc_hd__o21ai_1 _12198_ (.A1(_05329_),
    .A2(_05331_),
    .B1(_05325_),
    .Y(_05386_));
 sky130_fd_sc_hd__o22a_1 _12199_ (.A1(net17),
    .A2(net15),
    .B1(net6),
    .B2(net19),
    .X(_05387_));
 sky130_fd_sc_hd__xnor2_1 _12200_ (.A(net41),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _12201_ (.A(_05386_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__xnor2_1 _12202_ (.A(_05386_),
    .B(_05388_),
    .Y(_05390_));
 sky130_fd_sc_hd__or2_1 _12203_ (.A(net23),
    .B(net39),
    .X(_05391_));
 sky130_fd_sc_hd__xnor2_1 _12204_ (.A(_05390_),
    .B(_05391_),
    .Y(_05393_));
 sky130_fd_sc_hd__nor2_1 _12205_ (.A(net25),
    .B(net8),
    .Y(_05394_));
 sky130_fd_sc_hd__xnor2_1 _12206_ (.A(net66),
    .B(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__nor2_1 _12207_ (.A(_05393_),
    .B(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__and2_1 _12208_ (.A(_05393_),
    .B(_05395_),
    .X(_05397_));
 sky130_fd_sc_hd__nor3_1 _12209_ (.A(_05385_),
    .B(_05396_),
    .C(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__o21a_1 _12210_ (.A1(_05396_),
    .A2(_05397_),
    .B1(_05385_),
    .X(_05399_));
 sky130_fd_sc_hd__nor2_1 _12211_ (.A(_05398_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21ai_2 _12212_ (.A1(_05337_),
    .A2(_05341_),
    .B1(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__or3_1 _12213_ (.A(_05337_),
    .B(_05341_),
    .C(_05400_),
    .X(_05402_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_05401_),
    .B(_05402_),
    .Y(_05404_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_05279_),
    .B(_05346_),
    .Y(_05405_));
 sky130_fd_sc_hd__or4_1 _12216_ (.A(_04781_),
    .B(_05138_),
    .C(_05282_),
    .D(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__a21o_1 _12217_ (.A1(_05276_),
    .A2(_05343_),
    .B1(_05345_),
    .X(_05407_));
 sky130_fd_sc_hd__a21oi_1 _12218_ (.A1(_05137_),
    .A2(_05281_),
    .B1(_05280_),
    .Y(_05408_));
 sky130_fd_sc_hd__o211a_1 _12219_ (.A1(_05405_),
    .A2(_05408_),
    .B1(_05407_),
    .C1(_05406_),
    .X(_05409_));
 sky130_fd_sc_hd__xnor2_2 _12220_ (.A(_05404_),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__and3_1 _12221_ (.A(_05249_),
    .B(_05286_),
    .C(_05351_),
    .X(_05411_));
 sky130_fd_sc_hd__a21o_1 _12222_ (.A1(_05141_),
    .A2(_05411_),
    .B1(net149),
    .X(_05412_));
 sky130_fd_sc_hd__o21ai_1 _12223_ (.A1(_05410_),
    .A2(_05412_),
    .B1(net202),
    .Y(_05413_));
 sky130_fd_sc_hd__a21o_1 _12224_ (.A1(_05410_),
    .A2(_05412_),
    .B1(_05413_),
    .X(_05415_));
 sky130_fd_sc_hd__nor2_1 _12225_ (.A(net298),
    .B(_06401_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21oi_1 _12226_ (.A1(_05262_),
    .A2(_05355_),
    .B1(_05251_),
    .Y(_05417_));
 sky130_fd_sc_hd__a21o_1 _12227_ (.A1(net298),
    .A2(_05417_),
    .B1(_05416_),
    .X(_05418_));
 sky130_fd_sc_hd__o21ai_1 _12228_ (.A1(_05045_),
    .A2(_05418_),
    .B1(net242),
    .Y(_05419_));
 sky130_fd_sc_hd__a21o_1 _12229_ (.A1(_05045_),
    .A2(_05418_),
    .B1(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__nand2_1 _12230_ (.A(net157),
    .B(_02221_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21oi_1 _12231_ (.A1(_02224_),
    .A2(_05421_),
    .B1(_02318_),
    .Y(_05422_));
 sky130_fd_sc_hd__o21ai_1 _12232_ (.A1(_02224_),
    .A2(_05421_),
    .B1(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__o21ai_2 _12233_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05364_),
    .Y(_05424_));
 sky130_fd_sc_hd__xnor2_1 _12234_ (.A(reg1_val[28]),
    .B(_05424_),
    .Y(_05426_));
 sky130_fd_sc_hd__nor2_1 _12235_ (.A(net260),
    .B(_02821_),
    .Y(_05427_));
 sky130_fd_sc_hd__a211o_1 _12236_ (.A1(net260),
    .A2(_05426_),
    .B1(_05427_),
    .C1(net209),
    .X(_05428_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(\div_res[27] ),
    .B(_05374_),
    .X(_05429_));
 sky130_fd_sc_hd__a21oi_1 _12238_ (.A1(net155),
    .A2(_05429_),
    .B1(\div_res[28] ),
    .Y(_05430_));
 sky130_fd_sc_hd__a31o_1 _12239_ (.A1(\div_res[28] ),
    .A2(net155),
    .A3(_05429_),
    .B1(net198),
    .X(_05431_));
 sky130_fd_sc_hd__or2_1 _12240_ (.A(\div_shifter[59] ),
    .B(_05370_),
    .X(_05432_));
 sky130_fd_sc_hd__a21oi_1 _12241_ (.A1(net233),
    .A2(_05432_),
    .B1(\div_shifter[60] ),
    .Y(_05433_));
 sky130_fd_sc_hd__a31o_1 _12242_ (.A1(\div_shifter[60] ),
    .A2(net233),
    .A3(_05432_),
    .B1(net238),
    .X(_05434_));
 sky130_fd_sc_hd__o22ai_1 _12243_ (.A1(reg1_val[28]),
    .A2(_06432_),
    .B1(net200),
    .B2(_05023_),
    .Y(_05435_));
 sky130_fd_sc_hd__a21o_1 _12244_ (.A1(_05023_),
    .A2(_02326_),
    .B1(net273),
    .X(_05437_));
 sky130_fd_sc_hd__a221o_1 _12245_ (.A1(_02315_),
    .A2(_02821_),
    .B1(_05437_),
    .B2(_05034_),
    .C1(_05435_),
    .X(_05438_));
 sky130_fd_sc_hd__a21oi_2 _12246_ (.A1(net245),
    .A2(_02811_),
    .B1(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__o21a_1 _12247_ (.A1(_05433_),
    .A2(_05434_),
    .B1(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__o211a_1 _12248_ (.A1(_05430_),
    .A2(_05431_),
    .B1(_05440_),
    .C1(_05428_),
    .X(_05441_));
 sky130_fd_sc_hd__a41o_1 _12249_ (.A1(_05415_),
    .A2(_05420_),
    .A3(_05423_),
    .A4(_05441_),
    .B1(_06457_),
    .X(_05442_));
 sky130_fd_sc_hd__or2_1 _12250_ (.A(_05012_),
    .B(net251),
    .X(_05443_));
 sky130_fd_sc_hd__a21oi_4 _12251_ (.A1(_05442_),
    .A2(_05443_),
    .B1(net259),
    .Y(dest_val[28]));
 sky130_fd_sc_hd__o22a_1 _12252_ (.A1(net16),
    .A2(net8),
    .B1(net7),
    .B2(net17),
    .X(_05444_));
 sky130_fd_sc_hd__xnor2_1 _12253_ (.A(net42),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21bai_1 _12254_ (.A1(net19),
    .A2(net39),
    .B1_N(net67),
    .Y(_05447_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(net67),
    .B(net42),
    .Y(_05448_));
 sky130_fd_sc_hd__o21a_1 _12256_ (.A1(net19),
    .A2(_05448_),
    .B1(_05447_),
    .X(_05449_));
 sky130_fd_sc_hd__xnor2_1 _12257_ (.A(_05445_),
    .B(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__and2b_1 _12258_ (.A_N(_05450_),
    .B(_05395_),
    .X(_05451_));
 sky130_fd_sc_hd__and2b_1 _12259_ (.A_N(_05395_),
    .B(_05450_),
    .X(_05452_));
 sky130_fd_sc_hd__or2_1 _12260_ (.A(_05451_),
    .B(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__o21ai_1 _12261_ (.A1(_05390_),
    .A2(_05391_),
    .B1(_05389_),
    .Y(_05454_));
 sky130_fd_sc_hd__and2b_1 _12262_ (.A_N(_05453_),
    .B(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__xnor2_1 _12263_ (.A(_05453_),
    .B(_05454_),
    .Y(_05456_));
 sky130_fd_sc_hd__nor3_1 _12264_ (.A(_05396_),
    .B(_05398_),
    .C(_05456_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21a_1 _12265_ (.A1(_05396_),
    .A2(_05398_),
    .B1(_05456_),
    .X(_05459_));
 sky130_fd_sc_hd__or2_1 _12266_ (.A(_05458_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__a21boi_1 _12267_ (.A1(_05343_),
    .A2(_05401_),
    .B1_N(_05402_),
    .Y(_05461_));
 sky130_fd_sc_hd__a41o_1 _12268_ (.A1(_05346_),
    .A2(_05350_),
    .A3(_05401_),
    .A4(_05402_),
    .B1(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__and2b_1 _12269_ (.A_N(_05460_),
    .B(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__xor2_2 _12270_ (.A(_05460_),
    .B(_05462_),
    .X(_05464_));
 sky130_fd_sc_hd__a31o_1 _12271_ (.A1(_05141_),
    .A2(_05410_),
    .A3(_05411_),
    .B1(net149),
    .X(_05465_));
 sky130_fd_sc_hd__nor2_1 _12272_ (.A(_05464_),
    .B(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21o_1 _12273_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_02242_),
    .X(_05467_));
 sky130_fd_sc_hd__a21bo_1 _12274_ (.A1(_05034_),
    .A2(_05417_),
    .B1_N(_05023_),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_1 _12275_ (.A0(_06402_),
    .A1(_05469_),
    .S(net298),
    .X(_05470_));
 sky130_fd_sc_hd__nor2_1 _12276_ (.A(_04980_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__a21o_1 _12277_ (.A1(_04980_),
    .A2(_05470_),
    .B1(net241),
    .X(_05472_));
 sky130_fd_sc_hd__and2_1 _12278_ (.A(net151),
    .B(_02225_),
    .X(_05473_));
 sky130_fd_sc_hd__nor2_1 _12279_ (.A(_02229_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a211o_1 _12280_ (.A1(_02229_),
    .A2(_05473_),
    .B1(_05474_),
    .C1(_02318_),
    .X(_05475_));
 sky130_fd_sc_hd__and3_1 _12281_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_05424_),
    .X(_05476_));
 sky130_fd_sc_hd__a21oi_1 _12282_ (.A1(reg1_val[28]),
    .A2(_05424_),
    .B1(reg1_val[29]),
    .Y(_05477_));
 sky130_fd_sc_hd__o21a_1 _12283_ (.A1(_05476_),
    .A2(_05477_),
    .B1(net260),
    .X(_05478_));
 sky130_fd_sc_hd__nor2_1 _12284_ (.A(_06299_),
    .B(_02649_),
    .Y(_05480_));
 sky130_fd_sc_hd__or2_1 _12285_ (.A(\div_shifter[60] ),
    .B(_05432_),
    .X(_05481_));
 sky130_fd_sc_hd__a21oi_1 _12286_ (.A1(net234),
    .A2(_05481_),
    .B1(\div_shifter[61] ),
    .Y(_05482_));
 sky130_fd_sc_hd__a311o_2 _12287_ (.A1(\div_shifter[61] ),
    .A2(net234),
    .A3(_05481_),
    .B1(_05482_),
    .C1(net239),
    .X(_05483_));
 sky130_fd_sc_hd__or2_1 _12288_ (.A(\div_res[28] ),
    .B(_05429_),
    .X(_05484_));
 sky130_fd_sc_hd__a21oi_1 _12289_ (.A1(net155),
    .A2(_05484_),
    .B1(\div_res[29] ),
    .Y(_05485_));
 sky130_fd_sc_hd__a311o_1 _12290_ (.A1(\div_res[29] ),
    .A2(net155),
    .A3(_05484_),
    .B1(_05485_),
    .C1(net198),
    .X(_05486_));
 sky130_fd_sc_hd__a2bb2o_1 _12291_ (.A1_N(reg1_val[29]),
    .A2_N(_06432_),
    .B1(_02319_),
    .B2(_04958_),
    .X(_05487_));
 sky130_fd_sc_hd__o21ai_1 _12292_ (.A1(_04958_),
    .A2(_02327_),
    .B1(_02323_),
    .Y(_05488_));
 sky130_fd_sc_hd__a221o_1 _12293_ (.A1(_02315_),
    .A2(_02649_),
    .B1(_05488_),
    .B2(_04969_),
    .C1(_05487_),
    .X(_05489_));
 sky130_fd_sc_hd__a21oi_1 _12294_ (.A1(net245),
    .A2(_02663_),
    .B1(_05489_),
    .Y(_05491_));
 sky130_fd_sc_hd__and3_1 _12295_ (.A(_05483_),
    .B(_05486_),
    .C(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__o311a_1 _12296_ (.A1(net209),
    .A2(_05478_),
    .A3(_05480_),
    .B1(_05492_),
    .C1(_05475_),
    .X(_05493_));
 sky130_fd_sc_hd__o221a_1 _12297_ (.A1(_05466_),
    .A2(_05467_),
    .B1(_05471_),
    .B2(_05472_),
    .C1(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__o22a_2 _12298_ (.A1(_04947_),
    .A2(net251),
    .B1(_06457_),
    .B2(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__nor2_8 _12299_ (.A(net259),
    .B(_05495_),
    .Y(dest_val[29]));
 sky130_fd_sc_hd__o2bb2a_1 _12300_ (.A1_N(_05445_),
    .A2_N(_05449_),
    .B1(_05448_),
    .B2(net19),
    .X(_05496_));
 sky130_fd_sc_hd__or3_1 _12301_ (.A(net17),
    .B(net8),
    .C(_00665_),
    .X(_05497_));
 sky130_fd_sc_hd__o31ai_1 _12302_ (.A1(net66),
    .A2(_00408_),
    .A3(net8),
    .B1(net40),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_2 _12303_ (.A1(net8),
    .A2(_00665_),
    .B1(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__nor2_1 _12304_ (.A(_00377_),
    .B(net39),
    .Y(_05501_));
 sky130_fd_sc_hd__nor2_1 _12305_ (.A(_05499_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21a_1 _12306_ (.A1(_05499_),
    .A2(_05501_),
    .B1(_05497_),
    .X(_05503_));
 sky130_fd_sc_hd__xnor2_1 _12307_ (.A(_05496_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__or3_1 _12308_ (.A(_05451_),
    .B(_05455_),
    .C(_05504_),
    .X(_05505_));
 sky130_fd_sc_hd__o21a_1 _12309_ (.A1(_05451_),
    .A2(_05455_),
    .B1(_05504_),
    .X(_05506_));
 sky130_fd_sc_hd__o21ai_1 _12310_ (.A1(_05451_),
    .A2(_05455_),
    .B1(_05504_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _12311_ (.A(_05505_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__or2_1 _12312_ (.A(_05404_),
    .B(_05460_),
    .X(_05509_));
 sky130_fd_sc_hd__nor2_1 _12313_ (.A(_05405_),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__o22ai_1 _12314_ (.A1(_05401_),
    .A2(_05458_),
    .B1(_05509_),
    .B2(_05407_),
    .Y(_05512_));
 sky130_fd_sc_hd__a211o_1 _12315_ (.A1(_05285_),
    .A2(_05510_),
    .B1(_05512_),
    .C1(_05459_),
    .X(_05513_));
 sky130_fd_sc_hd__xor2_2 _12316_ (.A(_05508_),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__and2_1 _12317_ (.A(_05410_),
    .B(_05464_),
    .X(_05515_));
 sky130_fd_sc_hd__a41o_1 _12318_ (.A1(_05141_),
    .A2(_05410_),
    .A3(_05411_),
    .A4(_05464_),
    .B1(net149),
    .X(_05516_));
 sky130_fd_sc_hd__nor2_1 _12319_ (.A(_05514_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__a21o_1 _12320_ (.A1(_05514_),
    .A2(_05516_),
    .B1(_02242_),
    .X(_05518_));
 sky130_fd_sc_hd__a21o_1 _12321_ (.A1(_04969_),
    .A2(_05469_),
    .B1(_04958_),
    .X(_05519_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(_06403_),
    .A1(_05519_),
    .S(net298),
    .X(_05520_));
 sky130_fd_sc_hd__o21ai_1 _12323_ (.A1(_05479_),
    .A2(_05520_),
    .B1(_02324_),
    .Y(_05521_));
 sky130_fd_sc_hd__a21o_1 _12324_ (.A1(_05479_),
    .A2(_05520_),
    .B1(_05521_),
    .X(_05523_));
 sky130_fd_sc_hd__o21a_1 _12325_ (.A1(_02225_),
    .A2(_02229_),
    .B1(net151),
    .X(_05524_));
 sky130_fd_sc_hd__nor2_1 _12326_ (.A(_02232_),
    .B(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__a211o_1 _12327_ (.A1(_02232_),
    .A2(_05524_),
    .B1(_05525_),
    .C1(_02318_),
    .X(_05526_));
 sky130_fd_sc_hd__xor2_1 _12328_ (.A(reg1_val[30]),
    .B(_05476_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _12329_ (.A0(_02527_),
    .A1(_05527_),
    .S(net260),
    .X(_05528_));
 sky130_fd_sc_hd__or2_1 _12330_ (.A(\div_res[29] ),
    .B(_05484_),
    .X(_05529_));
 sky130_fd_sc_hd__a21o_1 _12331_ (.A1(net155),
    .A2(_05529_),
    .B1(\div_res[30] ),
    .X(_05530_));
 sky130_fd_sc_hd__nand3_1 _12332_ (.A(\div_res[30] ),
    .B(net155),
    .C(_05529_),
    .Y(_05531_));
 sky130_fd_sc_hd__o21a_1 _12333_ (.A1(_05457_),
    .A2(_02327_),
    .B1(_02323_),
    .X(_05532_));
 sky130_fd_sc_hd__o2bb2a_1 _12334_ (.A1_N(_05457_),
    .A2_N(net201),
    .B1(_06432_),
    .B2(reg1_val[30]),
    .X(_05534_));
 sky130_fd_sc_hd__o21ai_1 _12335_ (.A1(_05468_),
    .A2(_05532_),
    .B1(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__a221o_1 _12336_ (.A1(net246),
    .A2(_02501_),
    .B1(_02527_),
    .B2(_02315_),
    .C1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__or2_1 _12337_ (.A(\div_shifter[61] ),
    .B(_05481_),
    .X(_05537_));
 sky130_fd_sc_hd__a21oi_1 _12338_ (.A1(net234),
    .A2(_05537_),
    .B1(\div_shifter[62] ),
    .Y(_05538_));
 sky130_fd_sc_hd__a31o_1 _12339_ (.A1(\div_shifter[62] ),
    .A2(net234),
    .A3(_05537_),
    .B1(net239),
    .X(_05539_));
 sky130_fd_sc_hd__o21ai_1 _12340_ (.A1(_05538_),
    .A2(_05539_),
    .B1(_05526_),
    .Y(_05540_));
 sky130_fd_sc_hd__a311o_1 _12341_ (.A1(_02330_),
    .A2(_05530_),
    .A3(_05531_),
    .B1(_05536_),
    .C1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__a21oi_1 _12342_ (.A1(net210),
    .A2(_05528_),
    .B1(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__o211a_1 _12343_ (.A1(_05517_),
    .A2(_05518_),
    .B1(_05523_),
    .C1(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__o22a_2 _12344_ (.A1(_05436_),
    .A2(net251),
    .B1(_06457_),
    .B2(_05543_),
    .X(_05545_));
 sky130_fd_sc_hd__nor2_8 _12345_ (.A(net259),
    .B(_05545_),
    .Y(dest_val[30]));
 sky130_fd_sc_hd__a41oi_2 _12346_ (.A1(_05141_),
    .A2(_05411_),
    .A3(_05514_),
    .A4(_05515_),
    .B1(net149),
    .Y(_05546_));
 sky130_fd_sc_hd__o21a_1 _12347_ (.A1(_05496_),
    .A2(_05502_),
    .B1(_05497_),
    .X(_05547_));
 sky130_fd_sc_hd__xnor2_1 _12348_ (.A(_05499_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__nor2_1 _12349_ (.A(net10),
    .B(net40),
    .Y(_05549_));
 sky130_fd_sc_hd__xnor2_1 _12350_ (.A(_05548_),
    .B(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__o31a_1 _12351_ (.A1(_05459_),
    .A2(_05463_),
    .A3(_05506_),
    .B1(_05505_),
    .X(_05551_));
 sky130_fd_sc_hd__xnor2_1 _12352_ (.A(_05550_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand2_1 _12353_ (.A(_05546_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21a_1 _12354_ (.A1(_05546_),
    .A2(_05552_),
    .B1(_02241_),
    .X(_05555_));
 sky130_fd_sc_hd__a211o_1 _12355_ (.A1(_05479_),
    .A2(_05519_),
    .B1(net303),
    .C1(_05457_),
    .X(_05556_));
 sky130_fd_sc_hd__o21ai_1 _12356_ (.A1(net298),
    .A2(_06405_),
    .B1(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__xnor2_1 _12357_ (.A(_05403_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__o31a_1 _12358_ (.A1(_02225_),
    .A2(_02229_),
    .A3(_02232_),
    .B1(net151),
    .X(_05559_));
 sky130_fd_sc_hd__or2_1 _12359_ (.A(_02237_),
    .B(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__nand2_1 _12360_ (.A(_02237_),
    .B(_05559_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand3_1 _12361_ (.A(reg1_val[30]),
    .B(net260),
    .C(_05476_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _12362_ (.A(_02346_),
    .B(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__o211a_1 _12363_ (.A1(_02346_),
    .A2(_05562_),
    .B1(_05563_),
    .C1(net210),
    .X(_05564_));
 sky130_fd_sc_hd__o21a_1 _12364_ (.A1(\div_res[30] ),
    .A2(_05529_),
    .B1(net155),
    .X(_05566_));
 sky130_fd_sc_hd__o21ai_1 _12365_ (.A1(\div_res[31] ),
    .A2(_05566_),
    .B1(_02330_),
    .Y(_05567_));
 sky130_fd_sc_hd__a21oi_1 _12366_ (.A1(\div_res[31] ),
    .A2(_05566_),
    .B1(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__o21ai_1 _12367_ (.A1(\div_shifter[62] ),
    .A2(_05537_),
    .B1(net234),
    .Y(_05569_));
 sky130_fd_sc_hd__xnor2_1 _12368_ (.A(\div_shifter[63] ),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21ai_1 _12369_ (.A1(reg1_val[31]),
    .A2(net237),
    .B1(net251),
    .Y(_05571_));
 sky130_fd_sc_hd__or2_1 _12370_ (.A(reg1_val[31]),
    .B(_05392_),
    .X(_05572_));
 sky130_fd_sc_hd__a31o_1 _12371_ (.A1(reg1_val[31]),
    .A2(_05392_),
    .A3(net201),
    .B1(_05571_),
    .X(_05573_));
 sky130_fd_sc_hd__a221o_1 _12372_ (.A1(_05403_),
    .A2(_02326_),
    .B1(_05572_),
    .B2(net273),
    .C1(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__a221o_1 _12373_ (.A1(net246),
    .A2(_02310_),
    .B1(_02315_),
    .B2(_02347_),
    .C1(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__a211o_1 _12374_ (.A1(_02332_),
    .A2(_05570_),
    .B1(_05575_),
    .C1(_05568_),
    .X(_05577_));
 sky130_fd_sc_hd__a311o_1 _12375_ (.A1(_02317_),
    .A2(_05560_),
    .A3(_05561_),
    .B1(_05564_),
    .C1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__a221o_1 _12376_ (.A1(_05553_),
    .A2(_05555_),
    .B1(_05558_),
    .B2(_02324_),
    .C1(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__o211a_4 _12377_ (.A1(_05392_),
    .A2(net251),
    .B1(_05579_),
    .C1(net255),
    .X(dest_val[31]));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(net302),
    .A1(curr_PC[0]),
    .S(net254),
    .X(_05580_));
 sky130_fd_sc_hd__nand2_1 _12379_ (.A(_04849_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__or2_1 _12380_ (.A(_04849_),
    .B(_05580_),
    .X(_05582_));
 sky130_fd_sc_hd__and2_4 _12381_ (.A(_05581_),
    .B(_05582_),
    .X(new_PC[0]));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(net301),
    .A1(curr_PC[1]),
    .S(net255),
    .X(_05583_));
 sky130_fd_sc_hd__nand2_1 _12383_ (.A(_05987_),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__or2_1 _12384_ (.A(_05987_),
    .B(_05583_),
    .X(_05586_));
 sky130_fd_sc_hd__nand2_1 _12385_ (.A(_05584_),
    .B(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__or2_1 _12386_ (.A(_05581_),
    .B(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__nand2_1 _12387_ (.A(_05581_),
    .B(_05587_),
    .Y(_05589_));
 sky130_fd_sc_hd__and2_4 _12388_ (.A(_05588_),
    .B(_05589_),
    .X(new_PC[1]));
 sky130_fd_sc_hd__mux2_1 _12389_ (.A0(reg1_val[2]),
    .A1(curr_PC[2]),
    .S(net254),
    .X(_05590_));
 sky130_fd_sc_hd__nand2_1 _12390_ (.A(_05917_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__or2_1 _12391_ (.A(_05917_),
    .B(_05590_),
    .X(_05592_));
 sky130_fd_sc_hd__nand2_1 _12392_ (.A(_05591_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__a21o_1 _12393_ (.A1(_05584_),
    .A2(_05588_),
    .B1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__nand3_1 _12394_ (.A(_05584_),
    .B(_05588_),
    .C(_05593_),
    .Y(_05596_));
 sky130_fd_sc_hd__and2_4 _12395_ (.A(_05594_),
    .B(_05596_),
    .X(new_PC[2]));
 sky130_fd_sc_hd__mux2_1 _12396_ (.A0(reg1_val[3]),
    .A1(curr_PC[3]),
    .S(net254),
    .X(_05597_));
 sky130_fd_sc_hd__nand2_1 _12397_ (.A(_05845_),
    .B(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__or2_1 _12398_ (.A(_05845_),
    .B(_05597_),
    .X(_05599_));
 sky130_fd_sc_hd__nand2_1 _12399_ (.A(_05598_),
    .B(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__a21o_1 _12400_ (.A1(_05591_),
    .A2(_05594_),
    .B1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__nand3_1 _12401_ (.A(_05591_),
    .B(_05594_),
    .C(_05600_),
    .Y(_05602_));
 sky130_fd_sc_hd__and2_4 _12402_ (.A(_05601_),
    .B(_05602_),
    .X(new_PC[3]));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(reg1_val[4]),
    .A1(curr_PC[4]),
    .S(net256),
    .X(_05603_));
 sky130_fd_sc_hd__nand2_1 _12404_ (.A(_05782_),
    .B(_05603_),
    .Y(_05605_));
 sky130_fd_sc_hd__or2_1 _12405_ (.A(_05782_),
    .B(_05603_),
    .X(_05606_));
 sky130_fd_sc_hd__nand2_1 _12406_ (.A(_05605_),
    .B(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__a21o_1 _12407_ (.A1(_05598_),
    .A2(_05601_),
    .B1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__nand3_1 _12408_ (.A(_05598_),
    .B(_05601_),
    .C(_05607_),
    .Y(_05609_));
 sky130_fd_sc_hd__and2_4 _12409_ (.A(_05608_),
    .B(_05609_),
    .X(new_PC[4]));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(reg1_val[5]),
    .A1(curr_PC[5]),
    .S(net256),
    .X(_05610_));
 sky130_fd_sc_hd__nand2_1 _12411_ (.A(_05652_),
    .B(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__or2_1 _12412_ (.A(_05652_),
    .B(_05610_),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_05611_),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__a21o_1 _12414_ (.A1(_05605_),
    .A2(_05608_),
    .B1(_05613_),
    .X(_05615_));
 sky130_fd_sc_hd__nand3_1 _12415_ (.A(_05605_),
    .B(_05608_),
    .C(_05613_),
    .Y(_05616_));
 sky130_fd_sc_hd__and2_4 _12416_ (.A(_05615_),
    .B(_05616_),
    .X(new_PC[5]));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(reg1_val[6]),
    .A1(curr_PC[6]),
    .S(net256),
    .X(_05617_));
 sky130_fd_sc_hd__nand2_1 _12418_ (.A(_05718_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__or2_1 _12419_ (.A(_05718_),
    .B(_05617_),
    .X(_05619_));
 sky130_fd_sc_hd__nand2_1 _12420_ (.A(_05618_),
    .B(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__a21o_1 _12421_ (.A1(_05611_),
    .A2(_05615_),
    .B1(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__nand3_1 _12422_ (.A(_05611_),
    .B(_05615_),
    .C(_05620_),
    .Y(_05622_));
 sky130_fd_sc_hd__and2_4 _12423_ (.A(_05621_),
    .B(_05622_),
    .X(new_PC[6]));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(reg1_val[7]),
    .A1(curr_PC[7]),
    .S(net254),
    .X(_05624_));
 sky130_fd_sc_hd__nand2_1 _12425_ (.A(_05576_),
    .B(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hd__or2_1 _12426_ (.A(_05576_),
    .B(_05624_),
    .X(_05626_));
 sky130_fd_sc_hd__nand2_1 _12427_ (.A(_05625_),
    .B(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__a21o_1 _12428_ (.A1(_05618_),
    .A2(_05621_),
    .B1(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__nand3_1 _12429_ (.A(_05618_),
    .B(_05621_),
    .C(_05627_),
    .Y(_05629_));
 sky130_fd_sc_hd__and2_4 _12430_ (.A(_05628_),
    .B(_05629_),
    .X(new_PC[7]));
 sky130_fd_sc_hd__mux2_1 _12431_ (.A0(reg1_val[8]),
    .A1(curr_PC[8]),
    .S(net256),
    .X(_05630_));
 sky130_fd_sc_hd__nand2_1 _12432_ (.A(_05500_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__or2_1 _12433_ (.A(_05500_),
    .B(_05630_),
    .X(_05632_));
 sky130_fd_sc_hd__nand2_1 _12434_ (.A(_05631_),
    .B(_05632_),
    .Y(_05634_));
 sky130_fd_sc_hd__a21o_1 _12435_ (.A1(_05625_),
    .A2(_05628_),
    .B1(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__nand3_1 _12436_ (.A(_05625_),
    .B(_05628_),
    .C(_05634_),
    .Y(_05636_));
 sky130_fd_sc_hd__and2_4 _12437_ (.A(_05635_),
    .B(_05636_),
    .X(new_PC[8]));
 sky130_fd_sc_hd__mux2_1 _12438_ (.A0(reg1_val[9]),
    .A1(curr_PC[9]),
    .S(net256),
    .X(_05637_));
 sky130_fd_sc_hd__nand2_1 _12439_ (.A(_05132_),
    .B(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__or2_1 _12440_ (.A(_05132_),
    .B(_05637_),
    .X(_05639_));
 sky130_fd_sc_hd__nand2_1 _12441_ (.A(_05638_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__a21o_1 _12442_ (.A1(_05631_),
    .A2(_05635_),
    .B1(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__nand3_1 _12443_ (.A(_05631_),
    .B(_05635_),
    .C(_05640_),
    .Y(_05642_));
 sky130_fd_sc_hd__and2_4 _12444_ (.A(_05641_),
    .B(_05642_),
    .X(new_PC[9]));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(reg1_val[10]),
    .A1(curr_PC[10]),
    .S(net256),
    .X(_05644_));
 sky130_fd_sc_hd__nand2_1 _12446_ (.A(_05067_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__or2_1 _12447_ (.A(_05067_),
    .B(_05644_),
    .X(_05646_));
 sky130_fd_sc_hd__nand2_1 _12448_ (.A(_05645_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__a21o_1 _12449_ (.A1(_05638_),
    .A2(_05641_),
    .B1(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__nand3_1 _12450_ (.A(_05638_),
    .B(_05641_),
    .C(_05647_),
    .Y(_05649_));
 sky130_fd_sc_hd__and2_4 _12451_ (.A(_05648_),
    .B(_05649_),
    .X(new_PC[10]));
 sky130_fd_sc_hd__mux2_1 _12452_ (.A0(reg1_val[11]),
    .A1(curr_PC[11]),
    .S(net256),
    .X(_05650_));
 sky130_fd_sc_hd__nand2_1 _12453_ (.A(_05284_),
    .B(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__or2_1 _12454_ (.A(_05284_),
    .B(_05650_),
    .X(_05653_));
 sky130_fd_sc_hd__nand2_1 _12455_ (.A(_05651_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__a21o_1 _12456_ (.A1(_05645_),
    .A2(_05648_),
    .B1(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__nand3_1 _12457_ (.A(_05645_),
    .B(_05648_),
    .C(_05654_),
    .Y(_05656_));
 sky130_fd_sc_hd__and2_4 _12458_ (.A(_05655_),
    .B(_05656_),
    .X(new_PC[11]));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(reg1_val[12]),
    .A1(curr_PC[12]),
    .S(net257),
    .X(_05657_));
 sky130_fd_sc_hd__nand2_1 _12460_ (.A(_05208_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__or2_1 _12461_ (.A(_05208_),
    .B(_05657_),
    .X(_05659_));
 sky130_fd_sc_hd__nand2_1 _12462_ (.A(_05658_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__a21o_1 _12463_ (.A1(_05651_),
    .A2(_05655_),
    .B1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__nand3_1 _12464_ (.A(_05651_),
    .B(_05655_),
    .C(_05660_),
    .Y(_05663_));
 sky130_fd_sc_hd__and2_4 _12465_ (.A(_05661_),
    .B(_05663_),
    .X(new_PC[12]));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(reg1_val[13]),
    .A1(curr_PC[13]),
    .S(net256),
    .X(_05664_));
 sky130_fd_sc_hd__nand2_1 _12467_ (.A(_04991_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__or2_1 _12468_ (.A(_04991_),
    .B(_05664_),
    .X(_05666_));
 sky130_fd_sc_hd__nand2_1 _12469_ (.A(_05665_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__a21o_1 _12470_ (.A1(_05658_),
    .A2(_05661_),
    .B1(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__nand3_1 _12471_ (.A(_05658_),
    .B(_05661_),
    .C(_05667_),
    .Y(_05669_));
 sky130_fd_sc_hd__and2_4 _12472_ (.A(_05668_),
    .B(_05669_),
    .X(new_PC[13]));
 sky130_fd_sc_hd__mux2_1 _12473_ (.A0(reg1_val[14]),
    .A1(curr_PC[14]),
    .S(net256),
    .X(_05670_));
 sky130_fd_sc_hd__nand2_1 _12474_ (.A(_04925_),
    .B(_05670_),
    .Y(_05672_));
 sky130_fd_sc_hd__or2_1 _12475_ (.A(_04925_),
    .B(_05670_),
    .X(_05673_));
 sky130_fd_sc_hd__nand2_1 _12476_ (.A(_05672_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__a21o_1 _12477_ (.A1(_05665_),
    .A2(_05668_),
    .B1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__nand3_1 _12478_ (.A(_05665_),
    .B(_05668_),
    .C(_05674_),
    .Y(_05676_));
 sky130_fd_sc_hd__and2_4 _12479_ (.A(_05675_),
    .B(_05676_),
    .X(new_PC[14]));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(reg1_val[15]),
    .A1(curr_PC[15]),
    .S(net256),
    .X(_05677_));
 sky130_fd_sc_hd__nand2_1 _12481_ (.A(_05414_),
    .B(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__or2_1 _12482_ (.A(_05414_),
    .B(_05677_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _12483_ (.A(_05678_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__a21o_1 _12484_ (.A1(_05672_),
    .A2(_05675_),
    .B1(_05680_),
    .X(_05682_));
 sky130_fd_sc_hd__nand3_1 _12485_ (.A(_05672_),
    .B(_05675_),
    .C(_05680_),
    .Y(_05683_));
 sky130_fd_sc_hd__and2_4 _12486_ (.A(_05682_),
    .B(_05683_),
    .X(new_PC[15]));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(reg1_val[16]),
    .A1(curr_PC[16]),
    .S(net257),
    .X(_05684_));
 sky130_fd_sc_hd__xnor2_1 _12488_ (.A(net276),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__a21o_1 _12489_ (.A1(_05678_),
    .A2(_05682_),
    .B1(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__nand3_1 _12490_ (.A(_05678_),
    .B(_05682_),
    .C(_05685_),
    .Y(_05687_));
 sky130_fd_sc_hd__and2_4 _12491_ (.A(_05686_),
    .B(_05687_),
    .X(new_PC[16]));
 sky130_fd_sc_hd__mux2_2 _12492_ (.A0(reg1_val[17]),
    .A1(curr_PC[17]),
    .S(net256),
    .X(_05688_));
 sky130_fd_sc_hd__xnor2_4 _12493_ (.A(net276),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__a21bo_1 _12494_ (.A1(net276),
    .A2(_05684_),
    .B1_N(_05686_),
    .X(_05691_));
 sky130_fd_sc_hd__xnor2_4 _12495_ (.A(_05689_),
    .B(_05691_),
    .Y(new_PC[17]));
 sky130_fd_sc_hd__mux2_1 _12496_ (.A0(reg1_val[18]),
    .A1(curr_PC[18]),
    .S(net256),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _12497_ (.A(net276),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__or2_1 _12498_ (.A(net276),
    .B(_05692_),
    .X(_05694_));
 sky130_fd_sc_hd__nand2_1 _12499_ (.A(_05693_),
    .B(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__or2_1 _12500_ (.A(_05686_),
    .B(_05689_),
    .X(_05696_));
 sky130_fd_sc_hd__o21ai_1 _12501_ (.A1(_05684_),
    .A2(_05688_),
    .B1(net276),
    .Y(_05697_));
 sky130_fd_sc_hd__a21o_1 _12502_ (.A1(_05696_),
    .A2(_05697_),
    .B1(_05695_),
    .X(_05698_));
 sky130_fd_sc_hd__nand3_1 _12503_ (.A(_05695_),
    .B(_05696_),
    .C(_05697_),
    .Y(_05699_));
 sky130_fd_sc_hd__and2_4 _12504_ (.A(_05698_),
    .B(_05699_),
    .X(new_PC[18]));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(reg1_val[19]),
    .A1(curr_PC[19]),
    .S(net256),
    .X(_05701_));
 sky130_fd_sc_hd__nand2_1 _12506_ (.A(net276),
    .B(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__or2_1 _12507_ (.A(net276),
    .B(_05701_),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_2 _12508_ (.A(_05702_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_2 _12509_ (.A(_05693_),
    .B(_05698_),
    .Y(_05705_));
 sky130_fd_sc_hd__xnor2_4 _12510_ (.A(_05704_),
    .B(_05705_),
    .Y(new_PC[19]));
 sky130_fd_sc_hd__mux2_2 _12511_ (.A0(reg1_val[20]),
    .A1(curr_PC[20]),
    .S(net256),
    .X(_05706_));
 sky130_fd_sc_hd__nand2_1 _12512_ (.A(net277),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__or2_1 _12513_ (.A(net277),
    .B(_05706_),
    .X(_05708_));
 sky130_fd_sc_hd__nand2_2 _12514_ (.A(_05707_),
    .B(_05708_),
    .Y(_05710_));
 sky130_fd_sc_hd__or3_1 _12515_ (.A(_05695_),
    .B(_05696_),
    .C(_05704_),
    .X(_05711_));
 sky130_fd_sc_hd__and3_1 _12516_ (.A(_05693_),
    .B(_05697_),
    .C(_05702_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_2 _12517_ (.A(_05711_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__inv_2 _12518_ (.A(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__xnor2_4 _12519_ (.A(_05710_),
    .B(_05713_),
    .Y(new_PC[20]));
 sky130_fd_sc_hd__mux2_4 _12520_ (.A0(reg1_val[21]),
    .A1(curr_PC[21]),
    .S(net256),
    .X(_05715_));
 sky130_fd_sc_hd__xnor2_4 _12521_ (.A(net277),
    .B(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_2 _12522_ (.A1(_05710_),
    .A2(_05714_),
    .B1(_05707_),
    .Y(_05717_));
 sky130_fd_sc_hd__xnor2_4 _12523_ (.A(_05716_),
    .B(_05717_),
    .Y(new_PC[21]));
 sky130_fd_sc_hd__mux2_1 _12524_ (.A0(reg1_val[22]),
    .A1(curr_PC[22]),
    .S(net256),
    .X(_05719_));
 sky130_fd_sc_hd__and2_1 _12525_ (.A(net277),
    .B(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__or2_1 _12526_ (.A(net276),
    .B(_05719_),
    .X(_05721_));
 sky130_fd_sc_hd__nand2b_2 _12527_ (.A_N(_05720_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__o21ai_2 _12528_ (.A1(_05706_),
    .A2(_05715_),
    .B1(net276),
    .Y(_05723_));
 sky130_fd_sc_hd__nor2_1 _12529_ (.A(_05710_),
    .B(_05716_),
    .Y(_05724_));
 sky130_fd_sc_hd__inv_2 _12530_ (.A(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_4 _12531_ (.A1(_05714_),
    .A2(_05725_),
    .B1(_05723_),
    .Y(_05726_));
 sky130_fd_sc_hd__xnor2_4 _12532_ (.A(_05722_),
    .B(_05726_),
    .Y(new_PC[22]));
 sky130_fd_sc_hd__mux2_4 _12533_ (.A0(reg1_val[23]),
    .A1(curr_PC[23]),
    .S(net254),
    .X(_05727_));
 sky130_fd_sc_hd__xnor2_4 _12534_ (.A(net276),
    .B(_05727_),
    .Y(_05729_));
 sky130_fd_sc_hd__a21o_1 _12535_ (.A1(_05721_),
    .A2(_05726_),
    .B1(_05720_),
    .X(_05730_));
 sky130_fd_sc_hd__xnor2_4 _12536_ (.A(_05729_),
    .B(_05730_),
    .Y(new_PC[23]));
 sky130_fd_sc_hd__mux2_4 _12537_ (.A0(reg1_val[24]),
    .A1(curr_PC[24]),
    .S(net254),
    .X(_05731_));
 sky130_fd_sc_hd__xnor2_4 _12538_ (.A(net277),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__or4_1 _12539_ (.A(_05711_),
    .B(_05722_),
    .C(_05725_),
    .D(_05729_),
    .X(_05733_));
 sky130_fd_sc_hd__o21ai_1 _12540_ (.A1(_05719_),
    .A2(_05727_),
    .B1(net276),
    .Y(_05734_));
 sky130_fd_sc_hd__and4_2 _12541_ (.A(_05712_),
    .B(_05723_),
    .C(_05733_),
    .D(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__xor2_4 _12542_ (.A(_05732_),
    .B(_05735_),
    .X(new_PC[24]));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(reg1_val[25]),
    .A1(curr_PC[25]),
    .S(net254),
    .X(_05736_));
 sky130_fd_sc_hd__and2_1 _12544_ (.A(net276),
    .B(_05736_),
    .X(_05738_));
 sky130_fd_sc_hd__nor2_1 _12545_ (.A(net276),
    .B(_05736_),
    .Y(_05739_));
 sky130_fd_sc_hd__nor2_2 _12546_ (.A(_05738_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__o2bb2a_2 _12547_ (.A1_N(net277),
    .A2_N(_05731_),
    .B1(_05732_),
    .B2(_05735_),
    .X(_05741_));
 sky130_fd_sc_hd__xnor2_4 _12548_ (.A(_05740_),
    .B(_05741_),
    .Y(new_PC[25]));
 sky130_fd_sc_hd__mux2_2 _12549_ (.A0(reg1_val[26]),
    .A1(curr_PC[26]),
    .S(net254),
    .X(_05742_));
 sky130_fd_sc_hd__and2_1 _12550_ (.A(net276),
    .B(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__nor2_1 _12551_ (.A(net276),
    .B(_05742_),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_2 _12552_ (.A(_05743_),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ba_2 _12553_ (.A1(_05739_),
    .A2(_05741_),
    .B1_N(_05738_),
    .X(_05746_));
 sky130_fd_sc_hd__xnor2_4 _12554_ (.A(_05745_),
    .B(_05746_),
    .Y(new_PC[26]));
 sky130_fd_sc_hd__o21ba_1 _12555_ (.A1(_05744_),
    .A2(_05746_),
    .B1_N(_05743_),
    .X(_05748_));
 sky130_fd_sc_hd__mux2_2 _12556_ (.A0(reg1_val[27]),
    .A1(curr_PC[27]),
    .S(net254),
    .X(_05749_));
 sky130_fd_sc_hd__xor2_2 _12557_ (.A(net277),
    .B(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__xnor2_4 _12558_ (.A(_05748_),
    .B(_05750_),
    .Y(new_PC[27]));
 sky130_fd_sc_hd__nand2_2 _12559_ (.A(reg1_val[0]),
    .B(_04849_),
    .Y(_05751_));
 sky130_fd_sc_hd__or2_1 _12560_ (.A(reg1_val[0]),
    .B(_04849_),
    .X(_05752_));
 sky130_fd_sc_hd__and2_4 _12561_ (.A(_05751_),
    .B(_05752_),
    .X(loadstore_address[0]));
 sky130_fd_sc_hd__or2_1 _12562_ (.A(reg1_val[1]),
    .B(_05987_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(net301),
    .B(_05987_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_2 _12564_ (.A(_05753_),
    .B(_05754_),
    .Y(_05756_));
 sky130_fd_sc_hd__xor2_4 _12565_ (.A(_05751_),
    .B(_05756_),
    .X(loadstore_address[1]));
 sky130_fd_sc_hd__o21a_2 _12566_ (.A1(_05751_),
    .A2(_05756_),
    .B1(_05754_),
    .X(_05757_));
 sky130_fd_sc_hd__nor2_1 _12567_ (.A(reg1_val[2]),
    .B(_05917_),
    .Y(_05758_));
 sky130_fd_sc_hd__nand2_1 _12568_ (.A(reg1_val[2]),
    .B(_05917_),
    .Y(_05759_));
 sky130_fd_sc_hd__and2b_1 _12569_ (.A_N(_05758_),
    .B(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__xnor2_4 _12570_ (.A(_05757_),
    .B(_05760_),
    .Y(loadstore_address[2]));
 sky130_fd_sc_hd__o21a_2 _12571_ (.A1(_05757_),
    .A2(_05758_),
    .B1(_05759_),
    .X(_05761_));
 sky130_fd_sc_hd__nor2_1 _12572_ (.A(reg1_val[3]),
    .B(_05845_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _12573_ (.A(reg1_val[3]),
    .B(_05845_),
    .Y(_05763_));
 sky130_fd_sc_hd__and2b_1 _12574_ (.A_N(_05762_),
    .B(_05763_),
    .X(_05765_));
 sky130_fd_sc_hd__xnor2_4 _12575_ (.A(_05761_),
    .B(_05765_),
    .Y(loadstore_address[3]));
 sky130_fd_sc_hd__o21a_2 _12576_ (.A1(_05761_),
    .A2(_05762_),
    .B1(_05763_),
    .X(_05766_));
 sky130_fd_sc_hd__nor2_1 _12577_ (.A(reg1_val[4]),
    .B(_05782_),
    .Y(_05767_));
 sky130_fd_sc_hd__nand2_1 _12578_ (.A(reg1_val[4]),
    .B(_05782_),
    .Y(_05768_));
 sky130_fd_sc_hd__and2b_1 _12579_ (.A_N(_05767_),
    .B(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__xnor2_4 _12580_ (.A(_05766_),
    .B(_05769_),
    .Y(loadstore_address[4]));
 sky130_fd_sc_hd__o21a_2 _12581_ (.A1(_05766_),
    .A2(_05767_),
    .B1(_05768_),
    .X(_05770_));
 sky130_fd_sc_hd__nor2_1 _12582_ (.A(reg1_val[5]),
    .B(_05652_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _12583_ (.A(reg1_val[5]),
    .B(_05652_),
    .Y(_05772_));
 sky130_fd_sc_hd__nand2b_2 _12584_ (.A_N(_05771_),
    .B(_05772_),
    .Y(_05774_));
 sky130_fd_sc_hd__xor2_4 _12585_ (.A(_05770_),
    .B(_05774_),
    .X(loadstore_address[5]));
 sky130_fd_sc_hd__o21a_2 _12586_ (.A1(_05770_),
    .A2(_05771_),
    .B1(_05772_),
    .X(_05775_));
 sky130_fd_sc_hd__nor2_1 _12587_ (.A(reg1_val[6]),
    .B(_05718_),
    .Y(_05776_));
 sky130_fd_sc_hd__and2_1 _12588_ (.A(reg1_val[6]),
    .B(_05718_),
    .X(_05777_));
 sky130_fd_sc_hd__or2_2 _12589_ (.A(_05776_),
    .B(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__xor2_4 _12590_ (.A(_05775_),
    .B(_05778_),
    .X(loadstore_address[6]));
 sky130_fd_sc_hd__o21ba_2 _12591_ (.A1(_05775_),
    .A2(_05776_),
    .B1_N(_05777_),
    .X(_05779_));
 sky130_fd_sc_hd__nor2_1 _12592_ (.A(reg1_val[7]),
    .B(_05576_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand2_1 _12593_ (.A(reg1_val[7]),
    .B(_05576_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2b_2 _12594_ (.A_N(_05780_),
    .B(_05781_),
    .Y(_05783_));
 sky130_fd_sc_hd__xor2_4 _12595_ (.A(_05779_),
    .B(_05783_),
    .X(loadstore_address[7]));
 sky130_fd_sc_hd__o21a_2 _12596_ (.A1(_05779_),
    .A2(_05780_),
    .B1(_05781_),
    .X(_05784_));
 sky130_fd_sc_hd__nor2_1 _12597_ (.A(reg1_val[8]),
    .B(_05500_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_1 _12598_ (.A(reg1_val[8]),
    .B(_05500_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2b_2 _12599_ (.A_N(_05785_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__xor2_4 _12600_ (.A(_05784_),
    .B(_05787_),
    .X(loadstore_address[8]));
 sky130_fd_sc_hd__o21a_2 _12601_ (.A1(_05784_),
    .A2(_05785_),
    .B1(_05786_),
    .X(_05788_));
 sky130_fd_sc_hd__or2_1 _12602_ (.A(reg1_val[9]),
    .B(_05132_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _12603_ (.A(reg1_val[9]),
    .B(_05132_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_2 _12604_ (.A(_05789_),
    .B(_05790_),
    .Y(_05792_));
 sky130_fd_sc_hd__xor2_4 _12605_ (.A(_05788_),
    .B(_05792_),
    .X(loadstore_address[9]));
 sky130_fd_sc_hd__nand2_1 _12606_ (.A(reg1_val[10]),
    .B(_05067_),
    .Y(_05793_));
 sky130_fd_sc_hd__or2_1 _12607_ (.A(reg1_val[10]),
    .B(_05067_),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_1 _12608_ (.A(_05793_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2b_1 _12609_ (.A_N(_05788_),
    .B(_05789_),
    .Y(_05796_));
 sky130_fd_sc_hd__a21o_1 _12610_ (.A1(_05790_),
    .A2(_05796_),
    .B1(_05795_),
    .X(_05797_));
 sky130_fd_sc_hd__nand3_1 _12611_ (.A(_05790_),
    .B(_05795_),
    .C(_05796_),
    .Y(_05798_));
 sky130_fd_sc_hd__and2_4 _12612_ (.A(_05797_),
    .B(_05798_),
    .X(loadstore_address[10]));
 sky130_fd_sc_hd__nand2_1 _12613_ (.A(reg1_val[11]),
    .B(_05284_),
    .Y(_05799_));
 sky130_fd_sc_hd__or2_1 _12614_ (.A(reg1_val[11]),
    .B(_05284_),
    .X(_05801_));
 sky130_fd_sc_hd__nand2_1 _12615_ (.A(_05799_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__a21o_1 _12616_ (.A1(_05793_),
    .A2(_05797_),
    .B1(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__nand3_1 _12617_ (.A(_05793_),
    .B(_05797_),
    .C(_05802_),
    .Y(_05804_));
 sky130_fd_sc_hd__and2_4 _12618_ (.A(_05803_),
    .B(_05804_),
    .X(loadstore_address[11]));
 sky130_fd_sc_hd__nand2_1 _12619_ (.A(reg1_val[12]),
    .B(_05208_),
    .Y(_05805_));
 sky130_fd_sc_hd__or2_1 _12620_ (.A(reg1_val[12]),
    .B(_05208_),
    .X(_05806_));
 sky130_fd_sc_hd__nand2_1 _12621_ (.A(_05805_),
    .B(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__a21o_1 _12622_ (.A1(_05799_),
    .A2(_05803_),
    .B1(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__nand3_1 _12623_ (.A(_05799_),
    .B(_05803_),
    .C(_05807_),
    .Y(_05809_));
 sky130_fd_sc_hd__and2_4 _12624_ (.A(_05808_),
    .B(_05809_),
    .X(loadstore_address[12]));
 sky130_fd_sc_hd__nand2_1 _12625_ (.A(reg1_val[13]),
    .B(_04991_),
    .Y(_05811_));
 sky130_fd_sc_hd__or2_1 _12626_ (.A(reg1_val[13]),
    .B(_04991_),
    .X(_05812_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(_05811_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__a21o_1 _12628_ (.A1(_05805_),
    .A2(_05808_),
    .B1(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__nand3_1 _12629_ (.A(_05805_),
    .B(_05808_),
    .C(_05813_),
    .Y(_05815_));
 sky130_fd_sc_hd__and2_4 _12630_ (.A(_05814_),
    .B(_05815_),
    .X(loadstore_address[13]));
 sky130_fd_sc_hd__nand2_1 _12631_ (.A(reg1_val[14]),
    .B(_04925_),
    .Y(_05816_));
 sky130_fd_sc_hd__or2_1 _12632_ (.A(reg1_val[14]),
    .B(_04925_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_1 _12633_ (.A(_05816_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__a21o_1 _12634_ (.A1(_05811_),
    .A2(_05814_),
    .B1(_05818_),
    .X(_05820_));
 sky130_fd_sc_hd__nand3_1 _12635_ (.A(_05811_),
    .B(_05814_),
    .C(_05818_),
    .Y(_05821_));
 sky130_fd_sc_hd__and2_4 _12636_ (.A(_05820_),
    .B(_05821_),
    .X(loadstore_address[14]));
 sky130_fd_sc_hd__xnor2_2 _12637_ (.A(reg1_val[15]),
    .B(_05414_),
    .Y(_05822_));
 sky130_fd_sc_hd__a21oi_4 _12638_ (.A1(_05816_),
    .A2(_05820_),
    .B1(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__and3_2 _12639_ (.A(_05816_),
    .B(_05820_),
    .C(_05822_),
    .X(_05824_));
 sky130_fd_sc_hd__nor2_8 _12640_ (.A(_05823_),
    .B(_05824_),
    .Y(loadstore_address[15]));
 sky130_fd_sc_hd__xnor2_4 _12641_ (.A(_04531_),
    .B(_04817_),
    .Y(_05825_));
 sky130_fd_sc_hd__a21o_1 _12642_ (.A1(reg1_val[15]),
    .A2(_05414_),
    .B1(_05823_),
    .X(_05826_));
 sky130_fd_sc_hd__nand2_1 _12643_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__xor2_4 _12644_ (.A(_05825_),
    .B(_05826_),
    .X(loadstore_address[16]));
 sky130_fd_sc_hd__a21bo_1 _12645_ (.A1(reg1_val[16]),
    .A2(net278),
    .B1_N(_05827_),
    .X(_05829_));
 sky130_fd_sc_hd__xnor2_4 _12646_ (.A(reg1_val[17]),
    .B(net278),
    .Y(_05830_));
 sky130_fd_sc_hd__xnor2_4 _12647_ (.A(_05829_),
    .B(_05830_),
    .Y(loadstore_address[17]));
 sky130_fd_sc_hd__and2_1 _12648_ (.A(reg1_val[18]),
    .B(net278),
    .X(_05831_));
 sky130_fd_sc_hd__or2_1 _12649_ (.A(reg1_val[18]),
    .B(net278),
    .X(_05832_));
 sky130_fd_sc_hd__nand2b_2 _12650_ (.A_N(_05831_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__a2bb2o_2 _12651_ (.A1_N(_05827_),
    .A2_N(_05830_),
    .B1(net278),
    .B2(_06465_),
    .X(_05834_));
 sky130_fd_sc_hd__xnor2_4 _12652_ (.A(_05833_),
    .B(_05834_),
    .Y(loadstore_address[18]));
 sky130_fd_sc_hd__a21o_1 _12653_ (.A1(_05832_),
    .A2(_05834_),
    .B1(_05831_),
    .X(_05835_));
 sky130_fd_sc_hd__xnor2_4 _12654_ (.A(reg1_val[19]),
    .B(net278),
    .Y(_05837_));
 sky130_fd_sc_hd__xnor2_4 _12655_ (.A(_05835_),
    .B(_05837_),
    .Y(loadstore_address[19]));
 sky130_fd_sc_hd__xnor2_2 _12656_ (.A(reg1_val[20]),
    .B(net278),
    .Y(_05838_));
 sky130_fd_sc_hd__or4_2 _12657_ (.A(_05827_),
    .B(_05830_),
    .C(_05833_),
    .D(_05837_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_2 _12658_ (.A(_04817_),
    .B(_06466_),
    .Y(_05840_));
 sky130_fd_sc_hd__a21oi_4 _12659_ (.A1(_05839_),
    .A2(_05840_),
    .B1(_05838_),
    .Y(_05841_));
 sky130_fd_sc_hd__and3_2 _12660_ (.A(_05838_),
    .B(_05839_),
    .C(_05840_),
    .X(_05842_));
 sky130_fd_sc_hd__nor2_8 _12661_ (.A(_05841_),
    .B(_05842_),
    .Y(loadstore_address[20]));
 sky130_fd_sc_hd__nor2_1 _12662_ (.A(reg1_val[21]),
    .B(net278),
    .Y(_05843_));
 sky130_fd_sc_hd__nand2_2 _12663_ (.A(reg1_val[21]),
    .B(net278),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2b_2 _12664_ (.A_N(_05843_),
    .B(_05844_),
    .Y(_05846_));
 sky130_fd_sc_hd__a21oi_4 _12665_ (.A1(reg1_val[20]),
    .A2(net278),
    .B1(_05841_),
    .Y(_05847_));
 sky130_fd_sc_hd__xor2_4 _12666_ (.A(_05846_),
    .B(_05847_),
    .X(loadstore_address[21]));
 sky130_fd_sc_hd__and2_1 _12667_ (.A(reg1_val[22]),
    .B(net278),
    .X(_05848_));
 sky130_fd_sc_hd__or2_1 _12668_ (.A(reg1_val[22]),
    .B(net278),
    .X(_05849_));
 sky130_fd_sc_hd__nand2b_2 _12669_ (.A_N(_05848_),
    .B(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__o21ai_4 _12670_ (.A1(_05843_),
    .A2(_05847_),
    .B1(_05844_),
    .Y(_05851_));
 sky130_fd_sc_hd__xnor2_4 _12671_ (.A(_05850_),
    .B(_05851_),
    .Y(loadstore_address[22]));
 sky130_fd_sc_hd__a21o_1 _12672_ (.A1(_05849_),
    .A2(_05851_),
    .B1(_05848_),
    .X(_05852_));
 sky130_fd_sc_hd__xnor2_4 _12673_ (.A(reg1_val[23]),
    .B(net278),
    .Y(_05853_));
 sky130_fd_sc_hd__xnor2_4 _12674_ (.A(_05852_),
    .B(_05853_),
    .Y(loadstore_address[23]));
 sky130_fd_sc_hd__nand2_1 _12675_ (.A(reg1_val[24]),
    .B(net278),
    .Y(_05855_));
 sky130_fd_sc_hd__or2_1 _12676_ (.A(reg1_val[24]),
    .B(net279),
    .X(_05856_));
 sky130_fd_sc_hd__nand2_2 _12677_ (.A(_05855_),
    .B(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__or4_1 _12678_ (.A(_05838_),
    .B(_05846_),
    .C(_05850_),
    .D(_05853_),
    .X(_05858_));
 sky130_fd_sc_hd__a2bb2o_2 _12679_ (.A1_N(_05839_),
    .A2_N(_05858_),
    .B1(net278),
    .B2(_06467_),
    .X(_05859_));
 sky130_fd_sc_hd__nand2b_1 _12680_ (.A_N(_05857_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__xnor2_4 _12681_ (.A(_05857_),
    .B(_05859_),
    .Y(loadstore_address[24]));
 sky130_fd_sc_hd__nand2_2 _12682_ (.A(_05855_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__xnor2_4 _12683_ (.A(reg1_val[25]),
    .B(net279),
    .Y(_05862_));
 sky130_fd_sc_hd__xnor2_4 _12684_ (.A(_05861_),
    .B(_05862_),
    .Y(loadstore_address[25]));
 sky130_fd_sc_hd__and2_1 _12685_ (.A(reg1_val[26]),
    .B(net279),
    .X(_05864_));
 sky130_fd_sc_hd__or2_1 _12686_ (.A(reg1_val[26]),
    .B(net279),
    .X(_05865_));
 sky130_fd_sc_hd__nand2b_2 _12687_ (.A_N(_05864_),
    .B(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__or2_1 _12688_ (.A(_05860_),
    .B(_05862_),
    .X(_05867_));
 sky130_fd_sc_hd__a21bo_2 _12689_ (.A1(net279),
    .A2(_06468_),
    .B1_N(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__xnor2_4 _12690_ (.A(_05866_),
    .B(_05868_),
    .Y(loadstore_address[26]));
 sky130_fd_sc_hd__a21o_1 _12691_ (.A1(_05865_),
    .A2(_05868_),
    .B1(_05864_),
    .X(_05869_));
 sky130_fd_sc_hd__xnor2_2 _12692_ (.A(reg1_val[27]),
    .B(net279),
    .Y(_05870_));
 sky130_fd_sc_hd__xnor2_4 _12693_ (.A(_05869_),
    .B(_05870_),
    .Y(loadstore_address[27]));
 sky130_fd_sc_hd__and2_1 _12694_ (.A(reg1_val[28]),
    .B(net279),
    .X(_05872_));
 sky130_fd_sc_hd__nor2_1 _12695_ (.A(reg1_val[28]),
    .B(net279),
    .Y(_05873_));
 sky130_fd_sc_hd__or2_1 _12696_ (.A(_05872_),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_1 _12697_ (.A(net279),
    .B(_00218_),
    .Y(_05875_));
 sky130_fd_sc_hd__or3_1 _12698_ (.A(_05866_),
    .B(_05867_),
    .C(_05870_),
    .X(_05876_));
 sky130_fd_sc_hd__a21oi_2 _12699_ (.A1(_05875_),
    .A2(_05876_),
    .B1(_05874_),
    .Y(_05877_));
 sky130_fd_sc_hd__and3_2 _12700_ (.A(_05874_),
    .B(_05875_),
    .C(_05876_),
    .X(_05878_));
 sky130_fd_sc_hd__nor2_8 _12701_ (.A(_05877_),
    .B(_05878_),
    .Y(loadstore_address[28]));
 sky130_fd_sc_hd__or2_1 _12702_ (.A(reg1_val[29]),
    .B(net279),
    .X(_05879_));
 sky130_fd_sc_hd__nand2_1 _12703_ (.A(reg1_val[29]),
    .B(net279),
    .Y(_05880_));
 sky130_fd_sc_hd__nand2_2 _12704_ (.A(_05879_),
    .B(_05880_),
    .Y(_05882_));
 sky130_fd_sc_hd__or2_2 _12705_ (.A(_05872_),
    .B(_05877_),
    .X(_05883_));
 sky130_fd_sc_hd__xnor2_4 _12706_ (.A(_05882_),
    .B(_05883_),
    .Y(loadstore_address[29]));
 sky130_fd_sc_hd__and2_1 _12707_ (.A(reg1_val[30]),
    .B(net279),
    .X(_05884_));
 sky130_fd_sc_hd__or2_1 _12708_ (.A(reg1_val[30]),
    .B(net279),
    .X(_05885_));
 sky130_fd_sc_hd__nand2b_2 _12709_ (.A_N(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__a21bo_2 _12710_ (.A1(_05879_),
    .A2(_05883_),
    .B1_N(_05880_),
    .X(_05887_));
 sky130_fd_sc_hd__xnor2_4 _12711_ (.A(_05886_),
    .B(_05887_),
    .Y(loadstore_address[30]));
 sky130_fd_sc_hd__a21oi_1 _12712_ (.A1(_05885_),
    .A2(_05887_),
    .B1(_05884_),
    .Y(_05888_));
 sky130_fd_sc_hd__xnor2_2 _12713_ (.A(_04552_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__xnor2_4 _12714_ (.A(net278),
    .B(_05889_),
    .Y(loadstore_address[31]));
 sky130_fd_sc_hd__nand2_1 _12715_ (.A(net477),
    .B(net443),
    .Y(_05891_));
 sky130_fd_sc_hd__nand3_1 _12716_ (.A(net482),
    .B(net477),
    .C(net443),
    .Y(_05892_));
 sky130_fd_sc_hd__and4_1 _12717_ (.A(net460),
    .B(net482),
    .C(net477),
    .D(net443),
    .X(_05893_));
 sky130_fd_sc_hd__inv_2 _12718_ (.A(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__nand2_1 _12719_ (.A(net337),
    .B(_05893_),
    .Y(_05895_));
 sky130_fd_sc_hd__nor2_1 _12720_ (.A(net266),
    .B(net483),
    .Y(_05896_));
 sky130_fd_sc_hd__nor3_1 _12721_ (.A(rst),
    .B(net196),
    .C(_05896_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_4 _12722_ (.A(net271),
    .B(_06435_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_1 _12723_ (.A(net266),
    .B(_06434_),
    .Y(_05898_));
 sky130_fd_sc_hd__or2_1 _12724_ (.A(net339),
    .B(net179),
    .X(_05900_));
 sky130_fd_sc_hd__o211a_1 _12725_ (.A1(net45),
    .A2(net178),
    .B1(net340),
    .C1(net287),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _12726_ (.A(net216),
    .B(net182),
    .Y(_05901_));
 sky130_fd_sc_hd__o211a_1 _12727_ (.A1(net342),
    .A2(net181),
    .B1(_05901_),
    .C1(net292),
    .X(_00002_));
 sky130_fd_sc_hd__or2_1 _12728_ (.A(net351),
    .B(net181),
    .X(_05902_));
 sky130_fd_sc_hd__o211a_1 _12729_ (.A1(_00224_),
    .A2(net176),
    .B1(net352),
    .C1(net294),
    .X(_00003_));
 sky130_fd_sc_hd__nand2_1 _12730_ (.A(net158),
    .B(net181),
    .Y(_05903_));
 sky130_fd_sc_hd__o211a_1 _12731_ (.A1(net335),
    .A2(net181),
    .B1(_05903_),
    .C1(net294),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _12732_ (.A(net411),
    .B(net181),
    .X(_05904_));
 sky130_fd_sc_hd__o211a_1 _12733_ (.A1(_06491_),
    .A2(net177),
    .B1(net412),
    .C1(net294),
    .X(_00005_));
 sky130_fd_sc_hd__nand2_1 _12734_ (.A(net146),
    .B(net182),
    .Y(_05906_));
 sky130_fd_sc_hd__o211a_1 _12735_ (.A1(net333),
    .A2(net182),
    .B1(_05906_),
    .C1(net293),
    .X(_00006_));
 sky130_fd_sc_hd__nand2_1 _12736_ (.A(net139),
    .B(net182),
    .Y(_05907_));
 sky130_fd_sc_hd__o211a_1 _12737_ (.A1(net319),
    .A2(net182),
    .B1(_05907_),
    .C1(net293),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _12738_ (.A(net383),
    .B(net182),
    .X(_05908_));
 sky130_fd_sc_hd__o211a_1 _12739_ (.A1(_06522_),
    .A2(net177),
    .B1(net384),
    .C1(net296),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _12740_ (.A(net362),
    .B(net182),
    .X(_05909_));
 sky130_fd_sc_hd__o211a_1 _12741_ (.A1(_06513_),
    .A2(net177),
    .B1(net363),
    .C1(net293),
    .X(_00009_));
 sky130_fd_sc_hd__or2_1 _12742_ (.A(net379),
    .B(_05897_),
    .X(_05910_));
 sky130_fd_sc_hd__o211a_1 _12743_ (.A1(_06502_),
    .A2(net177),
    .B1(net380),
    .C1(net294),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _12744_ (.A(net369),
    .B(net181),
    .X(_05912_));
 sky130_fd_sc_hd__o211a_1 _12745_ (.A1(_00457_),
    .A2(net177),
    .B1(net370),
    .C1(net295),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _12746_ (.A(net360),
    .B(net182),
    .X(_05913_));
 sky130_fd_sc_hd__o211a_1 _12747_ (.A1(_00450_),
    .A2(net177),
    .B1(net361),
    .C1(net295),
    .X(_00012_));
 sky130_fd_sc_hd__or2_1 _12748_ (.A(net387),
    .B(net182),
    .X(_05914_));
 sky130_fd_sc_hd__o211a_1 _12749_ (.A1(_00445_),
    .A2(net177),
    .B1(net388),
    .C1(net293),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _12750_ (.A(net367),
    .B(net182),
    .X(_05915_));
 sky130_fd_sc_hd__o211a_1 _12751_ (.A1(_00436_),
    .A2(net177),
    .B1(net368),
    .C1(net293),
    .X(_00014_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(net92),
    .B(net182),
    .Y(_05916_));
 sky130_fd_sc_hd__o211a_1 _12753_ (.A1(net315),
    .A2(net182),
    .B1(_05916_),
    .C1(net293),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _12754_ (.A(net376),
    .B(net180),
    .X(_05918_));
 sky130_fd_sc_hd__o211a_1 _12755_ (.A1(_00323_),
    .A2(net178),
    .B1(net377),
    .C1(net290),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _12756_ (.A(net371),
    .B(net180),
    .X(_05919_));
 sky130_fd_sc_hd__o211a_1 _12757_ (.A1(_00310_),
    .A2(net178),
    .B1(net372),
    .C1(net290),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _12758_ (.A(net364),
    .B(net180),
    .X(_05920_));
 sky130_fd_sc_hd__o211a_1 _12759_ (.A1(_00300_),
    .A2(net178),
    .B1(net365),
    .C1(net290),
    .X(_00018_));
 sky130_fd_sc_hd__nand2_1 _12760_ (.A(net105),
    .B(net180),
    .Y(_05921_));
 sky130_fd_sc_hd__o211a_1 _12761_ (.A1(net317),
    .A2(net180),
    .B1(_05921_),
    .C1(net290),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_1 _12762_ (.A(net109),
    .B(net179),
    .Y(_05922_));
 sky130_fd_sc_hd__o211a_1 _12763_ (.A1(net331),
    .A2(net179),
    .B1(_05922_),
    .C1(net289),
    .X(_00020_));
 sky130_fd_sc_hd__or2_1 _12764_ (.A(net394),
    .B(net179),
    .X(_05924_));
 sky130_fd_sc_hd__o211a_1 _12765_ (.A1(_00211_),
    .A2(net178),
    .B1(net395),
    .C1(net291),
    .X(_00021_));
 sky130_fd_sc_hd__nand2_1 _12766_ (.A(net73),
    .B(net179),
    .Y(_05925_));
 sky130_fd_sc_hd__o211a_1 _12767_ (.A1(net329),
    .A2(net179),
    .B1(_05925_),
    .C1(net289),
    .X(_00022_));
 sky130_fd_sc_hd__nand2_1 _12768_ (.A(net76),
    .B(net179),
    .Y(_05926_));
 sky130_fd_sc_hd__o211a_1 _12769_ (.A1(net311),
    .A2(net179),
    .B1(_05926_),
    .C1(net289),
    .X(_00023_));
 sky130_fd_sc_hd__or2_1 _12770_ (.A(net392),
    .B(net179),
    .X(_05927_));
 sky130_fd_sc_hd__o211a_1 _12771_ (.A1(_00186_),
    .A2(net178),
    .B1(net393),
    .C1(net289),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _12772_ (.A(net63),
    .B(net179),
    .Y(_05928_));
 sky130_fd_sc_hd__o211a_1 _12773_ (.A1(net321),
    .A2(net179),
    .B1(_05928_),
    .C1(net289),
    .X(_00025_));
 sky130_fd_sc_hd__nand2_1 _12774_ (.A(_00246_),
    .B(net179),
    .Y(_05930_));
 sky130_fd_sc_hd__o211a_1 _12775_ (.A1(net325),
    .A2(net179),
    .B1(_05930_),
    .C1(net289),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _12776_ (.A(net59),
    .B(net179),
    .Y(_05931_));
 sky130_fd_sc_hd__o211a_1 _12777_ (.A1(net323),
    .A2(net179),
    .B1(_05931_),
    .C1(net289),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _12778_ (.A(net385),
    .B(net179),
    .X(_05932_));
 sky130_fd_sc_hd__o211a_1 _12779_ (.A1(_00284_),
    .A2(net178),
    .B1(net386),
    .C1(net289),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _12780_ (.A(net374),
    .B(net180),
    .X(_05933_));
 sky130_fd_sc_hd__o211a_1 _12781_ (.A1(_00271_),
    .A2(net178),
    .B1(net375),
    .C1(net290),
    .X(_00029_));
 sky130_fd_sc_hd__nand2_1 _12782_ (.A(net24),
    .B(net180),
    .Y(_05934_));
 sky130_fd_sc_hd__o211a_1 _12783_ (.A1(net313),
    .A2(net180),
    .B1(_05934_),
    .C1(net290),
    .X(_00030_));
 sky130_fd_sc_hd__nand2_1 _12784_ (.A(_00349_),
    .B(net180),
    .Y(_05936_));
 sky130_fd_sc_hd__o211a_1 _12785_ (.A1(net327),
    .A2(net180),
    .B1(_05936_),
    .C1(net290),
    .X(_00031_));
 sky130_fd_sc_hd__nand2_1 _12786_ (.A(_00377_),
    .B(net180),
    .Y(_05937_));
 sky130_fd_sc_hd__o211a_1 _12787_ (.A1(net309),
    .A2(net180),
    .B1(_05937_),
    .C1(net290),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _12788_ (.A(net381),
    .B(net182),
    .X(_05938_));
 sky130_fd_sc_hd__o211a_1 _12789_ (.A1(_00567_),
    .A2(net176),
    .B1(net382),
    .C1(net293),
    .X(_00033_));
 sky130_fd_sc_hd__or2_1 _12790_ (.A(_04411_),
    .B(net309),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_1 _12791_ (.A(_04411_),
    .B(net309),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_1 _12792_ (.A(_05939_),
    .B(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__nand2b_1 _12793_ (.A_N(net576),
    .B(net327),
    .Y(_05942_));
 sky130_fd_sc_hd__and2b_1 _12794_ (.A_N(net313),
    .B(net560),
    .X(_05944_));
 sky130_fd_sc_hd__nand2b_1 _12795_ (.A_N(net570),
    .B(net374),
    .Y(_05945_));
 sky130_fd_sc_hd__and2b_1 _12796_ (.A_N(net385),
    .B(\div_shifter[57] ),
    .X(_05946_));
 sky130_fd_sc_hd__nand2b_1 _12797_ (.A_N(\div_shifter[57] ),
    .B(net385),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2b_1 _12798_ (.A_N(_05946_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__nand2b_1 _12799_ (.A_N(net568),
    .B(net323),
    .Y(_05949_));
 sky130_fd_sc_hd__and2b_1 _12800_ (.A_N(net325),
    .B(net562),
    .X(_05950_));
 sky130_fd_sc_hd__nand2b_1 _12801_ (.A_N(\div_shifter[54] ),
    .B(net321),
    .Y(_05951_));
 sky130_fd_sc_hd__and2b_1 _12802_ (.A_N(net392),
    .B(net558),
    .X(_05952_));
 sky130_fd_sc_hd__nand2b_1 _12803_ (.A_N(net583),
    .B(net311),
    .Y(_05953_));
 sky130_fd_sc_hd__and2b_1 _12804_ (.A_N(net329),
    .B(\div_shifter[51] ),
    .X(_05955_));
 sky130_fd_sc_hd__nand2b_1 _12805_ (.A_N(\div_shifter[50] ),
    .B(net394),
    .Y(_05956_));
 sky130_fd_sc_hd__and2b_1 _12806_ (.A_N(net331),
    .B(net566),
    .X(_05957_));
 sky130_fd_sc_hd__nand2b_1 _12807_ (.A_N(net566),
    .B(net331),
    .Y(_05958_));
 sky130_fd_sc_hd__nand2b_1 _12808_ (.A_N(\div_shifter[48] ),
    .B(net317),
    .Y(_05959_));
 sky130_fd_sc_hd__nand2b_1 _12809_ (.A_N(net564),
    .B(net364),
    .Y(_05960_));
 sky130_fd_sc_hd__nand2b_1 _12810_ (.A_N(net588),
    .B(net371),
    .Y(_05961_));
 sky130_fd_sc_hd__nand2b_1 _12811_ (.A_N(\div_shifter[45] ),
    .B(net376),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2b_1 _12812_ (.A_N(net580),
    .B(net315),
    .Y(_05963_));
 sky130_fd_sc_hd__nand2b_1 _12813_ (.A_N(net597),
    .B(net367),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2b_1 _12814_ (.A_N(net582),
    .B(net387),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2b_1 _12815_ (.A_N(net578),
    .B(net360),
    .Y(_05967_));
 sky130_fd_sc_hd__nand2b_1 _12816_ (.A_N(net574),
    .B(net369),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2b_1 _12817_ (.A_N(\div_shifter[39] ),
    .B(net379),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2b_1 _12818_ (.A_N(net572),
    .B(net362),
    .Y(_05970_));
 sky130_fd_sc_hd__nand2b_1 _12819_ (.A_N(net590),
    .B(net383),
    .Y(_05971_));
 sky130_fd_sc_hd__and2b_1 _12820_ (.A_N(net319),
    .B(\div_shifter[36] ),
    .X(_05972_));
 sky130_fd_sc_hd__nand2b_1 _12821_ (.A_N(\div_shifter[36] ),
    .B(net319),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2b_1 _12822_ (.A_N(_05972_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__and2b_1 _12823_ (.A_N(net333),
    .B(net552),
    .X(_05975_));
 sky130_fd_sc_hd__nand2b_1 _12824_ (.A_N(net552),
    .B(net333),
    .Y(_05977_));
 sky130_fd_sc_hd__nand2b_1 _12825_ (.A_N(_05975_),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__nand2b_1 _12826_ (.A_N(net556),
    .B(net411),
    .Y(_05979_));
 sky130_fd_sc_hd__nand2b_1 _12827_ (.A_N(\div_shifter[33] ),
    .B(net335),
    .Y(_05980_));
 sky130_fd_sc_hd__and2b_1 _12828_ (.A_N(net351),
    .B(net546),
    .X(_05981_));
 sky130_fd_sc_hd__and2b_1 _12829_ (.A_N(net546),
    .B(net351),
    .X(_05982_));
 sky130_fd_sc_hd__nor2_1 _12830_ (.A(_05981_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__nand2b_1 _12831_ (.A_N(net344),
    .B(net342),
    .Y(_05984_));
 sky130_fd_sc_hd__a21o_1 _12832_ (.A1(_05983_),
    .A2(_05984_),
    .B1(_05981_),
    .X(_05985_));
 sky130_fd_sc_hd__nand2b_1 _12833_ (.A_N(net335),
    .B(\div_shifter[33] ),
    .Y(_05986_));
 sky130_fd_sc_hd__a21bo_1 _12834_ (.A1(_05980_),
    .A2(_05985_),
    .B1_N(_05986_),
    .X(_05988_));
 sky130_fd_sc_hd__nand2b_1 _12835_ (.A_N(net411),
    .B(net556),
    .Y(_05989_));
 sky130_fd_sc_hd__a21bo_1 _12836_ (.A1(_05979_),
    .A2(_05988_),
    .B1_N(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__a21o_1 _12837_ (.A1(_05977_),
    .A2(_05990_),
    .B1(_05975_),
    .X(_05991_));
 sky130_fd_sc_hd__a21o_1 _12838_ (.A1(_05973_),
    .A2(_05991_),
    .B1(_05972_),
    .X(_05992_));
 sky130_fd_sc_hd__nand2b_1 _12839_ (.A_N(net383),
    .B(net590),
    .Y(_05993_));
 sky130_fd_sc_hd__a21bo_1 _12840_ (.A1(_05971_),
    .A2(_05992_),
    .B1_N(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__nand2b_1 _12841_ (.A_N(net362),
    .B(net572),
    .Y(_05995_));
 sky130_fd_sc_hd__a21bo_1 _12842_ (.A1(_05970_),
    .A2(_05994_),
    .B1_N(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__nand2b_1 _12843_ (.A_N(net379),
    .B(\div_shifter[39] ),
    .Y(_05997_));
 sky130_fd_sc_hd__a21bo_1 _12844_ (.A1(_05969_),
    .A2(_05996_),
    .B1_N(_05997_),
    .X(_05999_));
 sky130_fd_sc_hd__nand2b_1 _12845_ (.A_N(net369),
    .B(net574),
    .Y(_06000_));
 sky130_fd_sc_hd__a21bo_1 _12846_ (.A1(_05968_),
    .A2(_05999_),
    .B1_N(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__nand2b_1 _12847_ (.A_N(net360),
    .B(net578),
    .Y(_06002_));
 sky130_fd_sc_hd__a21bo_1 _12848_ (.A1(_05967_),
    .A2(_06001_),
    .B1_N(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2b_1 _12849_ (.A_N(net387),
    .B(net582),
    .Y(_06004_));
 sky130_fd_sc_hd__a21bo_1 _12850_ (.A1(_05966_),
    .A2(_06003_),
    .B1_N(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__nand2b_1 _12851_ (.A_N(net367),
    .B(net597),
    .Y(_06006_));
 sky130_fd_sc_hd__a21bo_1 _12852_ (.A1(_05964_),
    .A2(_06005_),
    .B1_N(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__nand2b_1 _12853_ (.A_N(net315),
    .B(net580),
    .Y(_06008_));
 sky130_fd_sc_hd__a21bo_1 _12854_ (.A1(_05963_),
    .A2(_06007_),
    .B1_N(_06008_),
    .X(_06010_));
 sky130_fd_sc_hd__nand2b_1 _12855_ (.A_N(net376),
    .B(\div_shifter[45] ),
    .Y(_06011_));
 sky130_fd_sc_hd__a21bo_1 _12856_ (.A1(_05962_),
    .A2(_06010_),
    .B1_N(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__nand2b_1 _12857_ (.A_N(net371),
    .B(net588),
    .Y(_06013_));
 sky130_fd_sc_hd__a21bo_1 _12858_ (.A1(_05961_),
    .A2(_06012_),
    .B1_N(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__nand2b_1 _12859_ (.A_N(net364),
    .B(net564),
    .Y(_06015_));
 sky130_fd_sc_hd__a21bo_1 _12860_ (.A1(_05960_),
    .A2(_06014_),
    .B1_N(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__nand2b_1 _12861_ (.A_N(net317),
    .B(\div_shifter[48] ),
    .Y(_06017_));
 sky130_fd_sc_hd__a21bo_1 _12862_ (.A1(_05959_),
    .A2(_06016_),
    .B1_N(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__a21o_1 _12863_ (.A1(_05958_),
    .A2(_06018_),
    .B1(_05957_),
    .X(_06019_));
 sky130_fd_sc_hd__nand2b_1 _12864_ (.A_N(net394),
    .B(\div_shifter[50] ),
    .Y(_06021_));
 sky130_fd_sc_hd__a21bo_1 _12865_ (.A1(_05956_),
    .A2(_06019_),
    .B1_N(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2b_1 _12866_ (.A_N(\div_shifter[51] ),
    .B(net329),
    .Y(_06023_));
 sky130_fd_sc_hd__nand2b_1 _12867_ (.A_N(_05955_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__a21o_1 _12868_ (.A1(_06022_),
    .A2(_06023_),
    .B1(_05955_),
    .X(_06025_));
 sky130_fd_sc_hd__nand2b_1 _12869_ (.A_N(net311),
    .B(net583),
    .Y(_06026_));
 sky130_fd_sc_hd__a21bo_1 _12870_ (.A1(_05953_),
    .A2(_06025_),
    .B1_N(_06026_),
    .X(_06027_));
 sky130_fd_sc_hd__nand2b_1 _12871_ (.A_N(net558),
    .B(net392),
    .Y(_06028_));
 sky130_fd_sc_hd__nand2b_1 _12872_ (.A_N(_05952_),
    .B(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__a21o_1 _12873_ (.A1(_06027_),
    .A2(_06028_),
    .B1(_05952_),
    .X(_06030_));
 sky130_fd_sc_hd__nand2b_1 _12874_ (.A_N(net321),
    .B(\div_shifter[54] ),
    .Y(_06032_));
 sky130_fd_sc_hd__a21bo_1 _12875_ (.A1(_05951_),
    .A2(_06030_),
    .B1_N(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__nand2b_1 _12876_ (.A_N(net562),
    .B(net325),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2b_1 _12877_ (.A_N(_05950_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__a21o_1 _12878_ (.A1(_06033_),
    .A2(_06034_),
    .B1(_05950_),
    .X(_06036_));
 sky130_fd_sc_hd__nand2b_1 _12879_ (.A_N(net323),
    .B(net568),
    .Y(_06037_));
 sky130_fd_sc_hd__a21bo_1 _12880_ (.A1(_05949_),
    .A2(_06036_),
    .B1_N(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__a21o_1 _12881_ (.A1(_05947_),
    .A2(_06038_),
    .B1(_05946_),
    .X(_06039_));
 sky130_fd_sc_hd__nand2b_1 _12882_ (.A_N(net374),
    .B(net570),
    .Y(_06040_));
 sky130_fd_sc_hd__a21boi_1 _12883_ (.A1(_05945_),
    .A2(_06039_),
    .B1_N(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__and2b_1 _12884_ (.A_N(net560),
    .B(net313),
    .X(_06043_));
 sky130_fd_sc_hd__nor2_1 _12885_ (.A(_05944_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__o21bai_1 _12886_ (.A1(_06041_),
    .A2(_06043_),
    .B1_N(_05944_),
    .Y(_06045_));
 sky130_fd_sc_hd__nand2b_1 _12887_ (.A_N(net327),
    .B(net576),
    .Y(_06046_));
 sky130_fd_sc_hd__a21boi_1 _12888_ (.A1(_05942_),
    .A2(_06045_),
    .B1_N(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__or2_1 _12889_ (.A(_05941_),
    .B(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__a21oi_1 _12890_ (.A1(_05939_),
    .A2(_06048_),
    .B1(net381),
    .Y(_06049_));
 sky130_fd_sc_hd__and3_1 _12891_ (.A(net381),
    .B(_05939_),
    .C(_06048_),
    .X(_06050_));
 sky130_fd_sc_hd__o21bai_2 _12892_ (.A1(_04400_),
    .A2(_06050_),
    .B1_N(_06049_),
    .Y(_06051_));
 sky130_fd_sc_hd__a22o_1 _12893_ (.A1(net517),
    .A2(net194),
    .B1(net2),
    .B2(net268),
    .X(_06052_));
 sky130_fd_sc_hd__and2_1 _12894_ (.A(net288),
    .B(_06052_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _12895_ (.A1(net517),
    .A2(net268),
    .B1(net194),
    .B2(\div_res[1] ),
    .X(_06054_));
 sky130_fd_sc_hd__and2_1 _12896_ (.A(net288),
    .B(net518),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _12897_ (.A1(\div_res[1] ),
    .A2(net268),
    .B1(net194),
    .B2(net554),
    .X(_06055_));
 sky130_fd_sc_hd__and2_1 _12898_ (.A(net288),
    .B(net555),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _12899_ (.A1(net603),
    .A2(net268),
    .B1(net194),
    .B2(net523),
    .X(_06056_));
 sky130_fd_sc_hd__and2_1 _12900_ (.A(net288),
    .B(net524),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _12901_ (.A1(net523),
    .A2(net268),
    .B1(net194),
    .B2(net530),
    .X(_06057_));
 sky130_fd_sc_hd__and2_1 _12902_ (.A(net288),
    .B(net544),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _12903_ (.A1(net530),
    .A2(net267),
    .B1(net193),
    .B2(net495),
    .X(_06058_));
 sky130_fd_sc_hd__and2_1 _12904_ (.A(net288),
    .B(net531),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _12905_ (.A1(net495),
    .A2(net267),
    .B1(net193),
    .B2(\div_res[6] ),
    .X(_06060_));
 sky130_fd_sc_hd__and2_1 _12906_ (.A(net287),
    .B(net496),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _12907_ (.A1(net534),
    .A2(net267),
    .B1(net193),
    .B2(\div_res[7] ),
    .X(_06061_));
 sky130_fd_sc_hd__and2_1 _12908_ (.A(net287),
    .B(net535),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _12909_ (.A1(\div_res[7] ),
    .A2(net267),
    .B1(net193),
    .B2(net493),
    .X(_06062_));
 sky130_fd_sc_hd__and2_1 _12910_ (.A(net287),
    .B(net494),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _12911_ (.A1(net493),
    .A2(net267),
    .B1(net193),
    .B2(net504),
    .X(_06063_));
 sky130_fd_sc_hd__and2_1 _12912_ (.A(net287),
    .B(net505),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _12913_ (.A1(net504),
    .A2(net267),
    .B1(net193),
    .B2(net511),
    .X(_06064_));
 sky130_fd_sc_hd__and2_1 _12914_ (.A(net287),
    .B(net512),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _12915_ (.A1(net511),
    .A2(net267),
    .B1(net193),
    .B2(net525),
    .X(_06066_));
 sky130_fd_sc_hd__and2_1 _12916_ (.A(net287),
    .B(net526),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _12917_ (.A1(\div_res[11] ),
    .A2(net267),
    .B1(net193),
    .B2(net501),
    .X(_06067_));
 sky130_fd_sc_hd__and2_1 _12918_ (.A(net287),
    .B(net502),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _12919_ (.A1(net501),
    .A2(net267),
    .B1(net193),
    .B2(net521),
    .X(_06068_));
 sky130_fd_sc_hd__and2_1 _12920_ (.A(net287),
    .B(net522),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _12921_ (.A1(\div_res[13] ),
    .A2(net267),
    .B1(net193),
    .B2(net486),
    .X(_06069_));
 sky130_fd_sc_hd__and2_1 _12922_ (.A(net291),
    .B(net487),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _12923_ (.A1(net486),
    .A2(net268),
    .B1(net197),
    .B2(net509),
    .X(_06070_));
 sky130_fd_sc_hd__and2_1 _12924_ (.A(net288),
    .B(net510),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _12925_ (.A1(net509),
    .A2(net268),
    .B1(net194),
    .B2(net513),
    .X(_06072_));
 sky130_fd_sc_hd__and2_1 _12926_ (.A(net288),
    .B(_06072_),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _12927_ (.A1(net513),
    .A2(net269),
    .B1(net195),
    .B2(net484),
    .X(_06073_));
 sky130_fd_sc_hd__and2_1 _12928_ (.A(net290),
    .B(net514),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _12929_ (.A1(net484),
    .A2(net269),
    .B1(net193),
    .B2(net474),
    .X(_06074_));
 sky130_fd_sc_hd__and2_1 _12930_ (.A(net289),
    .B(net485),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _12931_ (.A1(net474),
    .A2(net269),
    .B1(net193),
    .B2(\div_res[19] ),
    .X(_06075_));
 sky130_fd_sc_hd__and2_1 _12932_ (.A(net287),
    .B(net475),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _12933_ (.A1(\div_res[19] ),
    .A2(net269),
    .B1(net194),
    .B2(net540),
    .X(_06076_));
 sky130_fd_sc_hd__and2_1 _12934_ (.A(net287),
    .B(net541),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _12935_ (.A1(\div_res[20] ),
    .A2(net267),
    .B1(net194),
    .B2(net527),
    .X(_06078_));
 sky130_fd_sc_hd__and2_1 _12936_ (.A(net287),
    .B(net528),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _12937_ (.A1(\div_res[21] ),
    .A2(net267),
    .B1(net194),
    .B2(net506),
    .X(_06079_));
 sky130_fd_sc_hd__and2_1 _12938_ (.A(net287),
    .B(net507),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _12939_ (.A1(\div_res[22] ),
    .A2(net267),
    .B1(net193),
    .B2(net498),
    .X(_06080_));
 sky130_fd_sc_hd__and2_1 _12940_ (.A(net287),
    .B(net499),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _12941_ (.A1(net498),
    .A2(net268),
    .B1(net194),
    .B2(net479),
    .X(_06081_));
 sky130_fd_sc_hd__and2_1 _12942_ (.A(net288),
    .B(net533),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _12943_ (.A1(net479),
    .A2(net267),
    .B1(net193),
    .B2(\div_res[25] ),
    .X(_06082_));
 sky130_fd_sc_hd__and2_1 _12944_ (.A(net287),
    .B(net480),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _12945_ (.A1(net515),
    .A2(net267),
    .B1(net193),
    .B2(net489),
    .X(_06084_));
 sky130_fd_sc_hd__and2_1 _12946_ (.A(net287),
    .B(net516),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _12947_ (.A1(net489),
    .A2(net267),
    .B1(net193),
    .B2(\div_res[27] ),
    .X(_06085_));
 sky130_fd_sc_hd__and2_1 _12948_ (.A(net288),
    .B(net490),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _12949_ (.A1(net519),
    .A2(net268),
    .B1(net194),
    .B2(net471),
    .X(_06086_));
 sky130_fd_sc_hd__and2_1 _12950_ (.A(net288),
    .B(net520),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _12951_ (.A1(net471),
    .A2(net268),
    .B1(net194),
    .B2(\div_res[29] ),
    .X(_06087_));
 sky130_fd_sc_hd__and2_1 _12952_ (.A(net288),
    .B(net472),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _12953_ (.A1(\div_res[29] ),
    .A2(net268),
    .B1(net194),
    .B2(net537),
    .X(_06088_));
 sky130_fd_sc_hd__and2_1 _12954_ (.A(net288),
    .B(net538),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _12955_ (.A1(\div_res[30] ),
    .A2(net268),
    .B1(net194),
    .B2(net455),
    .X(_06090_));
 sky130_fd_sc_hd__and2_1 _12956_ (.A(net288),
    .B(net456),
    .X(_00065_));
 sky130_fd_sc_hd__o22a_1 _12957_ (.A1(net347),
    .A2(net192),
    .B1(net177),
    .B2(net300),
    .X(_06091_));
 sky130_fd_sc_hd__nor2_1 _12958_ (.A(rst),
    .B(_06091_),
    .Y(_00066_));
 sky130_fd_sc_hd__a21oi_1 _12959_ (.A1(_04454_),
    .A2(net272),
    .B1(rst),
    .Y(_06092_));
 sky130_fd_sc_hd__o221a_1 _12960_ (.A1(net307),
    .A2(net192),
    .B1(net250),
    .B2(net177),
    .C1(_06092_),
    .X(_00067_));
 sky130_fd_sc_hd__o221a_1 _12961_ (.A1(net307),
    .A2(net266),
    .B1(net192),
    .B2(net389),
    .C1(net295),
    .X(_06093_));
 sky130_fd_sc_hd__a21boi_1 _12962_ (.A1(_00276_),
    .A2(_05897_),
    .B1_N(net390),
    .Y(_00068_));
 sky130_fd_sc_hd__o221a_1 _12963_ (.A1(net389),
    .A2(net266),
    .B1(net192),
    .B2(net463),
    .C1(net295),
    .X(_06094_));
 sky130_fd_sc_hd__a21boi_1 _12964_ (.A1(net205),
    .A2(net181),
    .B1_N(net464),
    .Y(_00069_));
 sky130_fd_sc_hd__o221a_1 _12965_ (.A1(net463),
    .A2(net266),
    .B1(net192),
    .B2(net465),
    .C1(net294),
    .X(_06096_));
 sky130_fd_sc_hd__a21boi_1 _12966_ (.A1(_00238_),
    .A2(_05897_),
    .B1_N(net466),
    .Y(_00070_));
 sky130_fd_sc_hd__o221a_1 _12967_ (.A1(\div_shifter[4] ),
    .A2(net266),
    .B1(net192),
    .B2(net452),
    .C1(net294),
    .X(_06097_));
 sky130_fd_sc_hd__a21boi_1 _12968_ (.A1(net208),
    .A2(net182),
    .B1_N(net453),
    .Y(_00071_));
 sky130_fd_sc_hd__o221a_1 _12969_ (.A1(net452),
    .A2(net266),
    .B1(net192),
    .B2(net427),
    .C1(net294),
    .X(_06098_));
 sky130_fd_sc_hd__a21boi_1 _12970_ (.A1(_00175_),
    .A2(net182),
    .B1_N(net459),
    .Y(_00072_));
 sky130_fd_sc_hd__o221a_1 _12971_ (.A1(net427),
    .A2(net266),
    .B1(net192),
    .B2(\div_shifter[7] ),
    .C1(net294),
    .X(_06099_));
 sky130_fd_sc_hd__a21boi_1 _12972_ (.A1(net185),
    .A2(_05897_),
    .B1_N(net428),
    .Y(_00073_));
 sky130_fd_sc_hd__o221a_1 _12973_ (.A1(\div_shifter[7] ),
    .A2(net266),
    .B1(net192),
    .B2(net440),
    .C1(net294),
    .X(_06100_));
 sky130_fd_sc_hd__a21boi_1 _12974_ (.A1(_00202_),
    .A2(net181),
    .B1_N(net441),
    .Y(_00074_));
 sky130_fd_sc_hd__o221a_1 _12975_ (.A1(net440),
    .A2(net266),
    .B1(net192),
    .B2(net446),
    .C1(net294),
    .X(_06102_));
 sky130_fd_sc_hd__a21boi_1 _12976_ (.A1(net187),
    .A2(net181),
    .B1_N(net447),
    .Y(_00075_));
 sky130_fd_sc_hd__o221a_1 _12977_ (.A1(net446),
    .A2(net266),
    .B1(net192),
    .B2(net450),
    .C1(net294),
    .X(_06103_));
 sky130_fd_sc_hd__a21boi_1 _12978_ (.A1(_00160_),
    .A2(net181),
    .B1_N(net451),
    .Y(_00076_));
 sky130_fd_sc_hd__o221a_1 _12979_ (.A1(\div_shifter[10] ),
    .A2(net265),
    .B1(net192),
    .B2(net401),
    .C1(net294),
    .X(_06104_));
 sky130_fd_sc_hd__o21a_1 _12980_ (.A1(_00146_),
    .A2(net177),
    .B1(net402),
    .X(_00077_));
 sky130_fd_sc_hd__o221a_1 _12981_ (.A1(net401),
    .A2(net265),
    .B1(net191),
    .B2(net438),
    .C1(net292),
    .X(_06105_));
 sky130_fd_sc_hd__a21boi_1 _12982_ (.A1(_00302_),
    .A2(net181),
    .B1_N(net468),
    .Y(_00078_));
 sky130_fd_sc_hd__o221a_1 _12983_ (.A1(net438),
    .A2(net266),
    .B1(net191),
    .B2(net404),
    .C1(net294),
    .X(_06106_));
 sky130_fd_sc_hd__a21boi_1 _12984_ (.A1(net130),
    .A2(net181),
    .B1_N(net439),
    .Y(_00079_));
 sky130_fd_sc_hd__o221a_1 _12985_ (.A1(net404),
    .A2(net265),
    .B1(net192),
    .B2(net396),
    .C1(net292),
    .X(_06108_));
 sky130_fd_sc_hd__a21boi_1 _12986_ (.A1(_00321_),
    .A2(net181),
    .B1_N(net405),
    .Y(_00080_));
 sky130_fd_sc_hd__o221a_1 _12987_ (.A1(net396),
    .A2(net265),
    .B1(net191),
    .B2(net348),
    .C1(net292),
    .X(_06109_));
 sky130_fd_sc_hd__o21a_1 _12988_ (.A1(_00319_),
    .A2(net176),
    .B1(net397),
    .X(_00081_));
 sky130_fd_sc_hd__o221a_1 _12989_ (.A1(net348),
    .A2(net265),
    .B1(net191),
    .B2(\div_shifter[16] ),
    .C1(net292),
    .X(_06110_));
 sky130_fd_sc_hd__a21boi_1 _12990_ (.A1(_00389_),
    .A2(net181),
    .B1_N(net349),
    .Y(_00082_));
 sky130_fd_sc_hd__o221a_1 _12991_ (.A1(\div_shifter[16] ),
    .A2(net266),
    .B1(net192),
    .B2(net419),
    .C1(net292),
    .X(_06111_));
 sky130_fd_sc_hd__o21a_1 _12992_ (.A1(net90),
    .A2(net176),
    .B1(net420),
    .X(_00083_));
 sky130_fd_sc_hd__o221a_1 _12993_ (.A1(net419),
    .A2(net265),
    .B1(net191),
    .B2(net422),
    .C1(net292),
    .X(_06112_));
 sky130_fd_sc_hd__o21a_1 _12994_ (.A1(_00432_),
    .A2(net176),
    .B1(net423),
    .X(_00084_));
 sky130_fd_sc_hd__o221a_1 _12995_ (.A1(\div_shifter[18] ),
    .A2(net265),
    .B1(net191),
    .B2(net416),
    .C1(net292),
    .X(_06114_));
 sky130_fd_sc_hd__o21a_1 _12996_ (.A1(net87),
    .A2(net176),
    .B1(net417),
    .X(_00085_));
 sky130_fd_sc_hd__o221a_1 _12997_ (.A1(net416),
    .A2(net265),
    .B1(net191),
    .B2(net434),
    .C1(net292),
    .X(_06115_));
 sky130_fd_sc_hd__o21a_1 _12998_ (.A1(_00448_),
    .A2(net176),
    .B1(net435),
    .X(_00086_));
 sky130_fd_sc_hd__o221a_1 _12999_ (.A1(\div_shifter[20] ),
    .A2(net265),
    .B1(net191),
    .B2(net413),
    .C1(net292),
    .X(_06116_));
 sky130_fd_sc_hd__o21a_1 _13000_ (.A1(net112),
    .A2(net176),
    .B1(net414),
    .X(_00087_));
 sky130_fd_sc_hd__o221a_1 _13001_ (.A1(net413),
    .A2(net265),
    .B1(net191),
    .B2(net432),
    .C1(net292),
    .X(_06117_));
 sky130_fd_sc_hd__o21a_1 _13002_ (.A1(_06507_),
    .A2(net176),
    .B1(net433),
    .X(_00088_));
 sky130_fd_sc_hd__o221a_1 _13003_ (.A1(\div_shifter[22] ),
    .A2(net265),
    .B1(net191),
    .B2(net406),
    .C1(net292),
    .X(_06118_));
 sky130_fd_sc_hd__o21a_1 _13004_ (.A1(net115),
    .A2(net176),
    .B1(net407),
    .X(_00089_));
 sky130_fd_sc_hd__o221a_1 _13005_ (.A1(net406),
    .A2(net265),
    .B1(net191),
    .B2(net436),
    .C1(net292),
    .X(_06120_));
 sky130_fd_sc_hd__o21a_1 _13006_ (.A1(_06524_),
    .A2(net176),
    .B1(net437),
    .X(_00090_));
 sky130_fd_sc_hd__o221a_1 _13007_ (.A1(\div_shifter[24] ),
    .A2(net265),
    .B1(net191),
    .B2(net424),
    .C1(net292),
    .X(_06121_));
 sky130_fd_sc_hd__o21a_1 _13008_ (.A1(net117),
    .A2(net176),
    .B1(net425),
    .X(_00091_));
 sky130_fd_sc_hd__o221a_1 _13009_ (.A1(net424),
    .A2(net265),
    .B1(net191),
    .B2(net430),
    .C1(net292),
    .X(_06122_));
 sky130_fd_sc_hd__o21a_1 _13010_ (.A1(_06483_),
    .A2(net176),
    .B1(net431),
    .X(_00092_));
 sky130_fd_sc_hd__o221a_1 _13011_ (.A1(\div_shifter[26] ),
    .A2(net265),
    .B1(net191),
    .B2(net398),
    .C1(net296),
    .X(_06123_));
 sky130_fd_sc_hd__o21a_1 _13012_ (.A1(net121),
    .A2(net176),
    .B1(net399),
    .X(_00093_));
 sky130_fd_sc_hd__o221a_1 _13013_ (.A1(net398),
    .A2(net265),
    .B1(net191),
    .B2(net357),
    .C1(net292),
    .X(_06124_));
 sky130_fd_sc_hd__o21a_1 _13014_ (.A1(_00227_),
    .A2(net176),
    .B1(net449),
    .X(_00094_));
 sky130_fd_sc_hd__a221o_1 _13015_ (.A1(net358),
    .A2(net272),
    .B1(net197),
    .B2(net354),
    .C1(rst),
    .X(_06126_));
 sky130_fd_sc_hd__a21oi_1 _13016_ (.A1(_00222_),
    .A2(net181),
    .B1(net359),
    .Y(_00095_));
 sky130_fd_sc_hd__a221o_1 _13017_ (.A1(net354),
    .A2(net272),
    .B1(net197),
    .B2(_04422_),
    .C1(rst),
    .X(_06127_));
 sky130_fd_sc_hd__a21oi_1 _13018_ (.A1(_00408_),
    .A2(net181),
    .B1(net355),
    .Y(_00096_));
 sky130_fd_sc_hd__a21oi_1 _13019_ (.A1(_04422_),
    .A2(net272),
    .B1(rst),
    .Y(_06128_));
 sky130_fd_sc_hd__o221a_1 _13020_ (.A1(net344),
    .A2(net191),
    .B1(net45),
    .B2(net176),
    .C1(_06128_),
    .X(_00097_));
 sky130_fd_sc_hd__nand3_1 _13021_ (.A(net344),
    .B(net342),
    .C(net1),
    .Y(_06129_));
 sky130_fd_sc_hd__a21o_1 _13022_ (.A1(net342),
    .A2(net1),
    .B1(net344),
    .X(_06130_));
 sky130_fd_sc_hd__a32o_1 _13023_ (.A1(net272),
    .A2(_06129_),
    .A3(_06130_),
    .B1(net197),
    .B2(net546),
    .X(_06131_));
 sky130_fd_sc_hd__and2_1 _13024_ (.A(net296),
    .B(net547),
    .X(_00098_));
 sky130_fd_sc_hd__xor2_1 _13025_ (.A(_05983_),
    .B(_05984_),
    .X(_06133_));
 sky130_fd_sc_hd__mux2_1 _13026_ (.A0(net546),
    .A1(_06133_),
    .S(net1),
    .X(_06134_));
 sky130_fd_sc_hd__a22o_1 _13027_ (.A1(net585),
    .A2(net197),
    .B1(_06134_),
    .B2(net272),
    .X(_06135_));
 sky130_fd_sc_hd__and2_1 _13028_ (.A(net296),
    .B(_06135_),
    .X(_00099_));
 sky130_fd_sc_hd__nand2_1 _13029_ (.A(_05980_),
    .B(_05986_),
    .Y(_06136_));
 sky130_fd_sc_hd__xnor2_1 _13030_ (.A(_05985_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(\div_shifter[33] ),
    .A1(_06137_),
    .S(net1),
    .X(_06138_));
 sky130_fd_sc_hd__a22o_1 _13032_ (.A1(net556),
    .A2(net196),
    .B1(_06138_),
    .B2(net271),
    .X(_06139_));
 sky130_fd_sc_hd__and2_1 _13033_ (.A(net293),
    .B(net557),
    .X(_00100_));
 sky130_fd_sc_hd__nand2_1 _13034_ (.A(_05979_),
    .B(_05989_),
    .Y(_06141_));
 sky130_fd_sc_hd__xnor2_1 _13035_ (.A(_05988_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__mux2_1 _13036_ (.A0(\div_shifter[34] ),
    .A1(_06142_),
    .S(net1),
    .X(_06143_));
 sky130_fd_sc_hd__a22o_1 _13037_ (.A1(net552),
    .A2(net196),
    .B1(_06143_),
    .B2(net271),
    .X(_06144_));
 sky130_fd_sc_hd__and2_1 _13038_ (.A(net293),
    .B(net553),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _13039_ (.A(_05978_),
    .B(_05990_),
    .Y(_06145_));
 sky130_fd_sc_hd__mux2_1 _13040_ (.A0(net552),
    .A1(_06145_),
    .S(net1),
    .X(_06146_));
 sky130_fd_sc_hd__a22o_1 _13041_ (.A1(net594),
    .A2(net196),
    .B1(_06146_),
    .B2(net271),
    .X(_06147_));
 sky130_fd_sc_hd__and2_1 _13042_ (.A(net293),
    .B(_06147_),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _13043_ (.A(_05974_),
    .B(_05991_),
    .Y(_06148_));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(\div_shifter[36] ),
    .A1(_06148_),
    .S(net549),
    .X(_06150_));
 sky130_fd_sc_hd__a22o_1 _13045_ (.A1(net590),
    .A2(net196),
    .B1(_06150_),
    .B2(net271),
    .X(_06151_));
 sky130_fd_sc_hd__and2_1 _13046_ (.A(net293),
    .B(net591),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _13047_ (.A(_05971_),
    .B(_05993_),
    .Y(_06152_));
 sky130_fd_sc_hd__xnor2_1 _13048_ (.A(_05992_),
    .B(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__mux2_1 _13049_ (.A0(\div_shifter[37] ),
    .A1(_06153_),
    .S(net1),
    .X(_06154_));
 sky130_fd_sc_hd__a22o_1 _13050_ (.A1(net572),
    .A2(net196),
    .B1(_06154_),
    .B2(net271),
    .X(_06155_));
 sky130_fd_sc_hd__and2_1 _13051_ (.A(net293),
    .B(net573),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_1 _13052_ (.A(_05970_),
    .B(_05995_),
    .Y(_06156_));
 sky130_fd_sc_hd__xnor2_1 _13053_ (.A(_05994_),
    .B(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__mux2_1 _13054_ (.A0(net572),
    .A1(_06157_),
    .S(net1),
    .X(_06159_));
 sky130_fd_sc_hd__a22o_1 _13055_ (.A1(net598),
    .A2(net196),
    .B1(_06159_),
    .B2(net271),
    .X(_06160_));
 sky130_fd_sc_hd__and2_1 _13056_ (.A(net294),
    .B(_06160_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(_05969_),
    .B(_05997_),
    .Y(_06161_));
 sky130_fd_sc_hd__xnor2_1 _13058_ (.A(_05996_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__mux2_1 _13059_ (.A0(\div_shifter[39] ),
    .A1(_06162_),
    .S(net1),
    .X(_06163_));
 sky130_fd_sc_hd__a22o_1 _13060_ (.A1(net574),
    .A2(net196),
    .B1(_06163_),
    .B2(net271),
    .X(_06164_));
 sky130_fd_sc_hd__and2_1 _13061_ (.A(net294),
    .B(net575),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_1 _13062_ (.A(_05968_),
    .B(_06000_),
    .Y(_06165_));
 sky130_fd_sc_hd__xnor2_1 _13063_ (.A(_05999_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__mux2_1 _13064_ (.A0(net574),
    .A1(_06166_),
    .S(net1),
    .X(_06168_));
 sky130_fd_sc_hd__a22o_1 _13065_ (.A1(net578),
    .A2(net197),
    .B1(_06168_),
    .B2(net271),
    .X(_06169_));
 sky130_fd_sc_hd__and2_1 _13066_ (.A(net294),
    .B(net579),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _13067_ (.A(_05967_),
    .B(_06002_),
    .Y(_06170_));
 sky130_fd_sc_hd__xnor2_1 _13068_ (.A(_06001_),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__mux2_1 _13069_ (.A0(net578),
    .A1(_06171_),
    .S(net1),
    .X(_06172_));
 sky130_fd_sc_hd__a22o_1 _13070_ (.A1(net582),
    .A2(net196),
    .B1(_06172_),
    .B2(net271),
    .X(_06173_));
 sky130_fd_sc_hd__and2_1 _13071_ (.A(net293),
    .B(_06173_),
    .X(_00108_));
 sky130_fd_sc_hd__nand2_1 _13072_ (.A(_05966_),
    .B(_06004_),
    .Y(_06174_));
 sky130_fd_sc_hd__xnor2_1 _13073_ (.A(_06003_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__mux2_1 _13074_ (.A0(net582),
    .A1(_06175_),
    .S(net549),
    .X(_06177_));
 sky130_fd_sc_hd__a22o_1 _13075_ (.A1(net597),
    .A2(net196),
    .B1(_06177_),
    .B2(net271),
    .X(_06178_));
 sky130_fd_sc_hd__and2_1 _13076_ (.A(net293),
    .B(_06178_),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _13077_ (.A(_05964_),
    .B(_06006_),
    .Y(_06179_));
 sky130_fd_sc_hd__xnor2_1 _13078_ (.A(_06005_),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(\div_shifter[43] ),
    .A1(_06180_),
    .S(net1),
    .X(_06181_));
 sky130_fd_sc_hd__a22o_1 _13080_ (.A1(net580),
    .A2(net196),
    .B1(_06181_),
    .B2(net271),
    .X(_06182_));
 sky130_fd_sc_hd__and2_1 _13081_ (.A(net293),
    .B(net581),
    .X(_00110_));
 sky130_fd_sc_hd__nand2_1 _13082_ (.A(_05963_),
    .B(_06008_),
    .Y(_06183_));
 sky130_fd_sc_hd__xnor2_1 _13083_ (.A(_06007_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(net580),
    .A1(_06184_),
    .S(net1),
    .X(_06186_));
 sky130_fd_sc_hd__a22o_1 _13085_ (.A1(net601),
    .A2(net195),
    .B1(_06186_),
    .B2(net271),
    .X(_06187_));
 sky130_fd_sc_hd__and2_1 _13086_ (.A(net293),
    .B(_06187_),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _13087_ (.A(_05962_),
    .B(_06011_),
    .Y(_06188_));
 sky130_fd_sc_hd__xnor2_1 _13088_ (.A(_06010_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(\div_shifter[45] ),
    .A1(_06189_),
    .S(net1),
    .X(_06190_));
 sky130_fd_sc_hd__a22o_1 _13090_ (.A1(net588),
    .A2(net195),
    .B1(_06190_),
    .B2(net270),
    .X(_06191_));
 sky130_fd_sc_hd__and2_1 _13091_ (.A(net290),
    .B(net589),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_1 _13092_ (.A(_05961_),
    .B(_06013_),
    .Y(_06192_));
 sky130_fd_sc_hd__xnor2_1 _13093_ (.A(_06012_),
    .B(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(\div_shifter[46] ),
    .A1(_06193_),
    .S(net2),
    .X(_06195_));
 sky130_fd_sc_hd__a22o_1 _13095_ (.A1(net564),
    .A2(net197),
    .B1(_06195_),
    .B2(net269),
    .X(_06196_));
 sky130_fd_sc_hd__and2_1 _13096_ (.A(net290),
    .B(net565),
    .X(_00113_));
 sky130_fd_sc_hd__nand2_1 _13097_ (.A(_05960_),
    .B(_06015_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_1 _13098_ (.A(_06014_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__mux2_1 _13099_ (.A0(net564),
    .A1(_06198_),
    .S(net2),
    .X(_06199_));
 sky130_fd_sc_hd__a22o_1 _13100_ (.A1(net600),
    .A2(net197),
    .B1(_06199_),
    .B2(net269),
    .X(_06200_));
 sky130_fd_sc_hd__and2_1 _13101_ (.A(net290),
    .B(_06200_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_1 _13102_ (.A(_05959_),
    .B(_06017_),
    .Y(_06201_));
 sky130_fd_sc_hd__xnor2_1 _13103_ (.A(_06016_),
    .B(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(\div_shifter[48] ),
    .A1(_06202_),
    .S(net2),
    .X(_06204_));
 sky130_fd_sc_hd__a22o_1 _13105_ (.A1(net566),
    .A2(net195),
    .B1(_06204_),
    .B2(net269),
    .X(_06205_));
 sky130_fd_sc_hd__and2_1 _13106_ (.A(net291),
    .B(net567),
    .X(_00115_));
 sky130_fd_sc_hd__nand2b_1 _13107_ (.A_N(_05957_),
    .B(_05958_),
    .Y(_06206_));
 sky130_fd_sc_hd__xnor2_1 _13108_ (.A(_06018_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__mux2_1 _13109_ (.A0(net566),
    .A1(_06207_),
    .S(net2),
    .X(_06208_));
 sky130_fd_sc_hd__a22o_1 _13110_ (.A1(net595),
    .A2(net195),
    .B1(_06208_),
    .B2(net269),
    .X(_06209_));
 sky130_fd_sc_hd__and2_1 _13111_ (.A(net291),
    .B(net596),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(_05956_),
    .B(_06021_),
    .Y(_06210_));
 sky130_fd_sc_hd__xnor2_1 _13113_ (.A(_06019_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__mux2_1 _13114_ (.A0(\div_shifter[50] ),
    .A1(_06211_),
    .S(net2),
    .X(_06213_));
 sky130_fd_sc_hd__a22o_1 _13115_ (.A1(net586),
    .A2(net195),
    .B1(_06213_),
    .B2(net269),
    .X(_06214_));
 sky130_fd_sc_hd__and2_1 _13116_ (.A(net291),
    .B(net587),
    .X(_00117_));
 sky130_fd_sc_hd__xnor2_1 _13117_ (.A(_06022_),
    .B(_06024_),
    .Y(_06215_));
 sky130_fd_sc_hd__mux2_1 _13118_ (.A0(\div_shifter[51] ),
    .A1(_06215_),
    .S(net2),
    .X(_06216_));
 sky130_fd_sc_hd__a22o_1 _13119_ (.A1(net583),
    .A2(net195),
    .B1(_06216_),
    .B2(net269),
    .X(_06217_));
 sky130_fd_sc_hd__and2_1 _13120_ (.A(net289),
    .B(net584),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _13121_ (.A(_05953_),
    .B(_06026_),
    .Y(_06218_));
 sky130_fd_sc_hd__xnor2_1 _13122_ (.A(_06025_),
    .B(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__mux2_1 _13123_ (.A0(\div_shifter[52] ),
    .A1(_06219_),
    .S(net2),
    .X(_06220_));
 sky130_fd_sc_hd__a22o_1 _13124_ (.A1(net558),
    .A2(net195),
    .B1(_06220_),
    .B2(net269),
    .X(_06222_));
 sky130_fd_sc_hd__and2_1 _13125_ (.A(net289),
    .B(net559),
    .X(_00119_));
 sky130_fd_sc_hd__xnor2_1 _13126_ (.A(_06027_),
    .B(_06029_),
    .Y(_06223_));
 sky130_fd_sc_hd__mux2_1 _13127_ (.A0(net558),
    .A1(_06223_),
    .S(net2),
    .X(_06224_));
 sky130_fd_sc_hd__a22o_1 _13128_ (.A1(net599),
    .A2(net195),
    .B1(_06224_),
    .B2(net269),
    .X(_06225_));
 sky130_fd_sc_hd__and2_1 _13129_ (.A(net289),
    .B(_06225_),
    .X(_00120_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(_05951_),
    .B(_06032_),
    .Y(_06226_));
 sky130_fd_sc_hd__xnor2_1 _13131_ (.A(_06030_),
    .B(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__mux2_1 _13132_ (.A0(\div_shifter[54] ),
    .A1(_06227_),
    .S(net2),
    .X(_06228_));
 sky130_fd_sc_hd__a22o_1 _13133_ (.A1(net562),
    .A2(net195),
    .B1(_06228_),
    .B2(net269),
    .X(_06229_));
 sky130_fd_sc_hd__and2_1 _13134_ (.A(net289),
    .B(net563),
    .X(_00121_));
 sky130_fd_sc_hd__xnor2_1 _13135_ (.A(_06033_),
    .B(_06035_),
    .Y(_06231_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(net562),
    .A1(_06231_),
    .S(net2),
    .X(_06232_));
 sky130_fd_sc_hd__a22o_1 _13137_ (.A1(net568),
    .A2(net195),
    .B1(_06232_),
    .B2(net269),
    .X(_06233_));
 sky130_fd_sc_hd__and2_1 _13138_ (.A(net289),
    .B(net569),
    .X(_00122_));
 sky130_fd_sc_hd__nand2_1 _13139_ (.A(_05949_),
    .B(_06037_),
    .Y(_06234_));
 sky130_fd_sc_hd__xnor2_1 _13140_ (.A(_06036_),
    .B(_06234_),
    .Y(_06235_));
 sky130_fd_sc_hd__mux2_1 _13141_ (.A0(net568),
    .A1(_06235_),
    .S(net2),
    .X(_06236_));
 sky130_fd_sc_hd__a22o_1 _13142_ (.A1(net592),
    .A2(net195),
    .B1(_06236_),
    .B2(net269),
    .X(_06237_));
 sky130_fd_sc_hd__and2_1 _13143_ (.A(net289),
    .B(_06237_),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_1 _13144_ (.A(_05948_),
    .B(_06038_),
    .Y(_06239_));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(\div_shifter[57] ),
    .A1(_06239_),
    .S(net2),
    .X(_06240_));
 sky130_fd_sc_hd__a22o_1 _13146_ (.A1(net570),
    .A2(net195),
    .B1(_06240_),
    .B2(net269),
    .X(_06241_));
 sky130_fd_sc_hd__and2_1 _13147_ (.A(net289),
    .B(net571),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(_05945_),
    .B(_06040_),
    .Y(_06242_));
 sky130_fd_sc_hd__xnor2_1 _13149_ (.A(_06039_),
    .B(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__mux2_1 _13150_ (.A0(\div_shifter[58] ),
    .A1(_06243_),
    .S(net2),
    .X(_06244_));
 sky130_fd_sc_hd__a22o_1 _13151_ (.A1(net560),
    .A2(net197),
    .B1(_06244_),
    .B2(net270),
    .X(_06245_));
 sky130_fd_sc_hd__and2_1 _13152_ (.A(net290),
    .B(net561),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_1 _13153_ (.A(_06041_),
    .B(_06044_),
    .Y(_06246_));
 sky130_fd_sc_hd__mux2_1 _13154_ (.A0(net560),
    .A1(_06246_),
    .S(net2),
    .X(_06248_));
 sky130_fd_sc_hd__a22o_1 _13155_ (.A1(net576),
    .A2(net195),
    .B1(_06248_),
    .B2(net270),
    .X(_06249_));
 sky130_fd_sc_hd__and2_1 _13156_ (.A(net290),
    .B(net577),
    .X(_00126_));
 sky130_fd_sc_hd__nand2_1 _13157_ (.A(_05942_),
    .B(_06046_),
    .Y(_06250_));
 sky130_fd_sc_hd__xnor2_1 _13158_ (.A(_06045_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(\div_shifter[60] ),
    .A1(_06251_),
    .S(net2),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_1 _13160_ (.A1(net550),
    .A2(net195),
    .B1(_06252_),
    .B2(net270),
    .X(_06253_));
 sky130_fd_sc_hd__and2_1 _13161_ (.A(net290),
    .B(net551),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_1 _13162_ (.A(_05941_),
    .B(_06047_),
    .Y(_06254_));
 sky130_fd_sc_hd__nor2_1 _13163_ (.A(_04411_),
    .B(net1),
    .Y(_06255_));
 sky130_fd_sc_hd__a31o_1 _13164_ (.A1(_06048_),
    .A2(net1),
    .A3(_06254_),
    .B1(_06255_),
    .X(_06257_));
 sky130_fd_sc_hd__a22o_1 _13165_ (.A1(net548),
    .A2(net195),
    .B1(_06257_),
    .B2(net270),
    .X(_06258_));
 sky130_fd_sc_hd__and2_1 _13166_ (.A(net290),
    .B(_06258_),
    .X(_00128_));
 sky130_fd_sc_hd__or3_1 _13167_ (.A(_04400_),
    .B(_06049_),
    .C(_06050_),
    .X(_06259_));
 sky130_fd_sc_hd__a32o_1 _13168_ (.A1(net593),
    .A2(net270),
    .A3(_06259_),
    .B1(net194),
    .B2(net409),
    .X(_06260_));
 sky130_fd_sc_hd__and2_1 _13169_ (.A(net288),
    .B(net410),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _13170_ (.A(net443),
    .B(net192),
    .Y(_06261_));
 sky130_fd_sc_hd__o211a_1 _13171_ (.A1(net443),
    .A2(net272),
    .B1(net295),
    .C1(net444),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _13172_ (.A1(net477),
    .A2(net196),
    .B1(_05891_),
    .B2(net272),
    .X(_06262_));
 sky130_fd_sc_hd__o211a_1 _13173_ (.A1(net477),
    .A2(net443),
    .B1(net295),
    .C1(_06262_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _13174_ (.A1(net482),
    .A2(net196),
    .B1(_05892_),
    .B2(net271),
    .X(_06264_));
 sky130_fd_sc_hd__a21o_1 _13175_ (.A1(net477),
    .A2(net443),
    .B1(net482),
    .X(_06265_));
 sky130_fd_sc_hd__and3_1 _13176_ (.A(net295),
    .B(_06264_),
    .C(net605),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _13177_ (.A1(net460),
    .A2(net196),
    .B1(_05894_),
    .B2(net271),
    .X(_06266_));
 sky130_fd_sc_hd__a31o_1 _13178_ (.A1(\div_counter[2] ),
    .A2(\div_counter[1] ),
    .A3(net443),
    .B1(net460),
    .X(_06267_));
 sky130_fd_sc_hd__and3_1 _13179_ (.A(net295),
    .B(_06266_),
    .C(net461),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13180_ (.A1(net337),
    .A2(net196),
    .B1(_05895_),
    .B2(net272),
    .X(_06268_));
 sky130_fd_sc_hd__o211a_1 _13181_ (.A1(net337),
    .A2(_05893_),
    .B1(_06268_),
    .C1(net295),
    .X(_00134_));
 sky130_fd_sc_hd__o21a_1 _13182_ (.A1(net469),
    .A2(_05896_),
    .B1(net295),
    .X(_00135_));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00000_),
    .Q(busy_l));
 sky130_fd_sc_hd__dfxtp_1 _13184_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net341),
    .Q(divi1_sign));
 sky130_fd_sc_hd__dfxtp_1 _13185_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net343),
    .Q(\divi2_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13186_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00003_),
    .Q(\divi2_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13187_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net336),
    .Q(\divi2_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13188_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00005_),
    .Q(\divi2_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13189_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net334),
    .Q(\divi2_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13190_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net320),
    .Q(\divi2_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13191_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00008_),
    .Q(\divi2_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13192_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00009_),
    .Q(\divi2_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13193_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00010_),
    .Q(\divi2_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13194_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00011_),
    .Q(\divi2_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13195_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00012_),
    .Q(\divi2_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13196_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00013_),
    .Q(\divi2_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13197_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00014_),
    .Q(\divi2_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13198_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net316),
    .Q(\divi2_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13199_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net378),
    .Q(\divi2_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13200_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net373),
    .Q(\divi2_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13201_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net366),
    .Q(\divi2_l[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13202_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net318),
    .Q(\divi2_l[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13203_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net332),
    .Q(\divi2_l[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13204_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00021_),
    .Q(\divi2_l[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13205_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net330),
    .Q(\divi2_l[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13206_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net312),
    .Q(\divi2_l[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13207_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00024_),
    .Q(\divi2_l[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13208_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net322),
    .Q(\divi2_l[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13209_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net326),
    .Q(\divi2_l[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13210_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net324),
    .Q(\divi2_l[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13211_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00028_),
    .Q(\divi2_l[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13212_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00029_),
    .Q(\divi2_l[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13213_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net314),
    .Q(\divi2_l[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13214_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net328),
    .Q(\divi2_l[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13215_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net310),
    .Q(\divi2_l[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13216_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00033_),
    .Q(\divi2_l[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13217_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00034_),
    .Q(\div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13218_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00035_),
    .Q(\div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13219_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00036_),
    .Q(\div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13220_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00037_),
    .Q(\div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13221_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00038_),
    .Q(\div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00039_),
    .Q(\div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13223_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net497),
    .Q(\div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13224_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net536),
    .Q(\div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00042_),
    .Q(\div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00043_),
    .Q(\div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00044_),
    .Q(\div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13228_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00045_),
    .Q(\div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net503),
    .Q(\div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00047_),
    .Q(\div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net488),
    .Q(\div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00049_),
    .Q(\div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00050_),
    .Q(\div_res[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00051_),
    .Q(\div_res[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00052_),
    .Q(\div_res[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net476),
    .Q(\div_res[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net542),
    .Q(\div_res[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net529),
    .Q(\div_res[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13239_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net508),
    .Q(\div_res[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net500),
    .Q(\div_res[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00058_),
    .Q(\div_res[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net481),
    .Q(\div_res[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00060_),
    .Q(\div_res[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net491),
    .Q(\div_res[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00062_),
    .Q(\div_res[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net473),
    .Q(\div_res[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net539),
    .Q(\div_res[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net457),
    .Q(\div_res[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00066_),
    .Q(\div_shifter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net308),
    .Q(\div_shifter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net391),
    .Q(\div_shifter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00069_),
    .Q(\div_shifter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00070_),
    .Q(\div_shifter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net454),
    .Q(\div_shifter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00072_),
    .Q(\div_shifter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net429),
    .Q(\div_shifter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net442),
    .Q(\div_shifter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00075_),
    .Q(\div_shifter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00076_),
    .Q(\div_shifter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net403),
    .Q(\div_shifter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00078_),
    .Q(\div_shifter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00079_),
    .Q(\div_shifter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00080_),
    .Q(\div_shifter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00081_),
    .Q(\div_shifter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net350),
    .Q(\div_shifter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net421),
    .Q(\div_shifter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00084_),
    .Q(\div_shifter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net418),
    .Q(\div_shifter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00086_),
    .Q(\div_shifter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net415),
    .Q(\div_shifter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00088_),
    .Q(\div_shifter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net408),
    .Q(\div_shifter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00090_),
    .Q(\div_shifter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13274_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net426),
    .Q(\div_shifter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00092_),
    .Q(\div_shifter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net400),
    .Q(\div_shifter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00094_),
    .Q(\div_shifter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00095_),
    .Q(\div_shifter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net356),
    .Q(\div_shifter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net345),
    .Q(\div_shifter[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00098_),
    .Q(\div_shifter[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00099_),
    .Q(\div_shifter[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00100_),
    .Q(\div_shifter[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00101_),
    .Q(\div_shifter[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00102_),
    .Q(\div_shifter[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00103_),
    .Q(\div_shifter[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00104_),
    .Q(\div_shifter[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00105_),
    .Q(\div_shifter[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00106_),
    .Q(\div_shifter[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00107_),
    .Q(\div_shifter[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00108_),
    .Q(\div_shifter[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00109_),
    .Q(\div_shifter[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00110_),
    .Q(\div_shifter[44] ));
 sky130_fd_sc_hd__dfxtp_2 _13294_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00111_),
    .Q(\div_shifter[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00112_),
    .Q(\div_shifter[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00113_),
    .Q(\div_shifter[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00114_),
    .Q(\div_shifter[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00115_),
    .Q(\div_shifter[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00116_),
    .Q(\div_shifter[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00117_),
    .Q(\div_shifter[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00118_),
    .Q(\div_shifter[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00119_),
    .Q(\div_shifter[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00120_),
    .Q(\div_shifter[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00121_),
    .Q(\div_shifter[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00122_),
    .Q(\div_shifter[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00123_),
    .Q(\div_shifter[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00124_),
    .Q(\div_shifter[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00125_),
    .Q(\div_shifter[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00126_),
    .Q(\div_shifter[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00127_),
    .Q(\div_shifter[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00128_),
    .Q(\div_shifter[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00129_),
    .Q(\div_shifter[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net445),
    .Q(\div_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net478),
    .Q(\div_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net606),
    .Q(\div_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net462),
    .Q(\div_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net338),
    .Q(\div_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net470),
    .Q(div_complete));
 sky130_fd_sc_hd__buf_12 _13319_ (.A(instruction[11]),
    .X(loadstore_dest[0]));
 sky130_fd_sc_hd__buf_12 _13320_ (.A(instruction[12]),
    .X(loadstore_dest[1]));
 sky130_fd_sc_hd__buf_12 _13321_ (.A(instruction[13]),
    .X(loadstore_dest[2]));
 sky130_fd_sc_hd__buf_12 _13322_ (.A(instruction[14]),
    .X(loadstore_dest[3]));
 sky130_fd_sc_hd__buf_12 _13323_ (.A(instruction[15]),
    .X(loadstore_dest[4]));
 sky130_fd_sc_hd__buf_12 _13324_ (.A(instruction[16]),
    .X(loadstore_dest[5]));
 sky130_fd_sc_hd__buf_12 _13325_ (.A(instruction[5]),
    .X(loadstore_size[0]));
 sky130_fd_sc_hd__buf_12 _13326_ (.A(instruction[6]),
    .X(loadstore_size[1]));
 sky130_fd_sc_hd__buf_12 _13327_ (.A(instruction[8]),
    .X(pred_idx[0]));
 sky130_fd_sc_hd__buf_12 _13328_ (.A(instruction[9]),
    .X(pred_idx[1]));
 sky130_fd_sc_hd__buf_12 _13329_ (.A(instruction[10]),
    .X(pred_idx[2]));
 sky130_fd_sc_hd__buf_12 _13330_ (.A(instruction[4]),
    .X(sign_extend));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout1 (.A(_06051_),
    .X(net1));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(_00299_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_00167_),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(_00166_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_00163_),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_16 fanout109 (.A(_00155_),
    .X(net109));
 sky130_fd_sc_hd__buf_8 fanout11 (.A(_00454_),
    .X(net11));
 sky130_fd_sc_hd__buf_12 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_12 fanout112 (.A(_06504_),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_16 fanout113 (.A(_06498_),
    .X(net113));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(_06498_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_16 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(_06482_),
    .X(net117));
 sky130_fd_sc_hd__buf_12 fanout118 (.A(_06482_),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout12 (.A(_00454_),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_16 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_16 fanout121 (.A(_06471_),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(_00456_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(_00456_),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(_00451_),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(_00451_),
    .X(net125));
 sky130_fd_sc_hd__buf_12 fanout126 (.A(net128),
    .X(net126));
 sky130_fd_sc_hd__buf_12 fanout127 (.A(_00320_),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_16 fanout129 (.A(_00298_),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__buf_12 fanout130 (.A(_00298_),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(_00298_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(_00213_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(_00205_),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(_00189_),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(_00189_),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_8 fanout139 (.A(_00136_),
    .X(net139));
 sky130_fd_sc_hd__buf_6 fanout14 (.A(_00440_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_8 fanout141 (.A(_06523_),
    .X(net141));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_6 fanout143 (.A(_06512_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_6 fanout145 (.A(_06501_),
    .X(net145));
 sky130_fd_sc_hd__buf_6 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_8 fanout147 (.A(_06479_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(_02135_),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net157),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net157),
    .X(net152));
 sky130_fd_sc_hd__buf_2 fanout153 (.A(net157),
    .X(net153));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(net156),
    .X(net154));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(_02134_),
    .X(net157));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(_00411_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_8 fanout159 (.A(_00411_),
    .X(net159));
 sky130_fd_sc_hd__buf_8 fanout16 (.A(_00409_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_8 fanout160 (.A(_00286_),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(_00286_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(_00282_),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(_00248_),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(_00248_),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(_00242_),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(_00242_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(_00225_),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout17 (.A(_00377_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(_00179_),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(_00179_),
    .X(net171));
 sky130_fd_sc_hd__buf_12 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_12 fanout173 (.A(_00145_),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(_06490_),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(_06490_),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_05898_),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(_05897_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout18 (.A(_00377_),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(_05897_),
    .X(net180));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_05897_),
    .X(net182));
 sky130_fd_sc_hd__buf_8 fanout183 (.A(_00171_),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(_00171_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_16 fanout185 (.A(_00171_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_16 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__buf_8 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_16 fanout188 (.A(_00158_),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(_06474_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout19 (.A(_00349_),
    .X(net19));
 sky130_fd_sc_hd__buf_6 fanout190 (.A(_06473_),
    .X(net190));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(_06437_),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net197),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(net197),
    .X(net195));
 sky130_fd_sc_hd__buf_6 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(_06436_),
    .X(net197));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(_02331_),
    .X(net198));
 sky130_fd_sc_hd__buf_2 fanout199 (.A(_02331_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout2 (.A(_06051_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_8 fanout20 (.A(_00349_),
    .X(net20));
 sky130_fd_sc_hd__buf_6 fanout200 (.A(_02320_),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(_02241_),
    .X(net202));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(_00236_),
    .X(net203));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(_00236_),
    .X(net204));
 sky130_fd_sc_hd__buf_12 fanout205 (.A(_00236_),
    .X(net205));
 sky130_fd_sc_hd__buf_8 fanout206 (.A(_00173_),
    .X(net206));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(_00173_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_16 fanout208 (.A(_00173_),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 fanout209 (.A(_06447_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 fanout21 (.A(_00270_),
    .X(net21));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(_06446_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_6 fanout213 (.A(_06333_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(_06332_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(net219),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(_06328_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_8 fanout22 (.A(_00270_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(_06322_),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(_06315_),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(_06314_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(_06309_),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_8 fanout226 (.A(net228),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(_06308_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(_06300_),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_8 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(_04915_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(_04915_),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(_02515_),
    .X(net232));
 sky130_fd_sc_hd__buf_2 fanout233 (.A(_02515_),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(_02515_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(_02515_),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(_02334_),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(_02333_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(_02333_),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout24 (.A(_00264_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 fanout241 (.A(_02325_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_8 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net246),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_8 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(_02246_),
    .X(net246));
 sky130_fd_sc_hd__buf_6 fanout247 (.A(_00266_),
    .X(net247));
 sky130_fd_sc_hd__buf_12 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_12 fanout249 (.A(_00256_),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_8 fanout251 (.A(_06456_),
    .X(net251));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(_06456_),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__buf_6 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net257),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_6 fanout257 (.A(_06428_),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_16 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_8 fanout259 (.A(_06427_),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout26 (.A(_00231_),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(_06299_),
    .X(net261));
 sky130_fd_sc_hd__buf_6 fanout262 (.A(net264),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_4 fanout264 (.A(_04893_),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(_04465_),
    .X(net266));
 sky130_fd_sc_hd__buf_4 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(net270),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_6 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout270 (.A(net458),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_8 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net458),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(_02322_),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_8 fanout275 (.A(_06458_),
    .X(net275));
 sky130_fd_sc_hd__buf_6 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(_04817_),
    .X(net277));
 sky130_fd_sc_hd__buf_12 fanout278 (.A(_04817_),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout279 (.A(_04817_),
    .X(net279));
 sky130_fd_sc_hd__buf_8 fanout28 (.A(_00230_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(_04806_),
    .X(net280));
 sky130_fd_sc_hd__buf_2 fanout281 (.A(_04806_),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_8 fanout282 (.A(_04806_),
    .X(net282));
 sky130_fd_sc_hd__buf_6 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 fanout284 (.A(_04795_),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(_04607_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net291),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(net291),
    .X(net289));
 sky130_fd_sc_hd__buf_6 fanout29 (.A(_00138_),
    .X(net29));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_2 fanout291 (.A(_04574_),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(net296),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(net296),
    .X(net293));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net296),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(_04574_),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_8 fanout297 (.A(_04563_),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_8 fanout298 (.A(_04563_),
    .X(net298));
 sky130_fd_sc_hd__buf_6 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout30 (.A(_00138_),
    .X(net30));
 sky130_fd_sc_hd__buf_6 fanout300 (.A(_04498_),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_16 fanout301 (.A(reg1_val[1]),
    .X(net301));
 sky130_fd_sc_hd__buf_6 fanout302 (.A(reg1_val[0]),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_8 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_6 fanout304 (.A(instruction[7]),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_8 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(instruction[6]),
    .X(net306));
 sky130_fd_sc_hd__buf_6 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__buf_6 fanout32 (.A(_06527_),
    .X(net32));
 sky130_fd_sc_hd__buf_8 fanout33 (.A(_06516_),
    .X(net33));
 sky130_fd_sc_hd__buf_4 fanout34 (.A(_06516_),
    .X(net34));
 sky130_fd_sc_hd__buf_6 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(_06493_),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(_06487_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_8 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_8 fanout40 (.A(_00662_),
    .X(net40));
 sky130_fd_sc_hd__buf_8 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_8 fanout42 (.A(net45),
    .X(net42));
 sky130_fd_sc_hd__buf_12 fanout43 (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_8 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_6 fanout45 (.A(_00661_),
    .X(net45));
 sky130_fd_sc_hd__buf_6 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_8 fanout47 (.A(_00449_),
    .X(net47));
 sky130_fd_sc_hd__buf_6 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_8 fanout49 (.A(_00433_),
    .X(net49));
 sky130_fd_sc_hd__buf_6 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_8 fanout51 (.A(_00394_),
    .X(net51));
 sky130_fd_sc_hd__buf_8 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(_00392_),
    .X(net53));
 sky130_fd_sc_hd__buf_6 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_8 fanout55 (.A(_00327_),
    .X(net55));
 sky130_fd_sc_hd__buf_8 fanout56 (.A(_00313_),
    .X(net56));
 sky130_fd_sc_hd__buf_6 fanout57 (.A(_00311_),
    .X(net57));
 sky130_fd_sc_hd__buf_6 fanout58 (.A(_00289_),
    .X(net58));
 sky130_fd_sc_hd__buf_6 fanout59 (.A(_00289_),
    .X(net59));
 sky130_fd_sc_hd__buf_6 fanout6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 fanout60 (.A(_00285_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(_00285_),
    .X(net61));
 sky130_fd_sc_hd__buf_6 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_8 fanout63 (.A(_00251_),
    .X(net63));
 sky130_fd_sc_hd__buf_6 fanout64 (.A(_00246_),
    .X(net64));
 sky130_fd_sc_hd__buf_6 fanout65 (.A(_00246_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 fanout66 (.A(net68),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_12 fanout68 (.A(_00222_),
    .X(net68));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_6 fanout7 (.A(_00666_),
    .X(net7));
 sky130_fd_sc_hd__buf_8 fanout70 (.A(_00210_),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(net73),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_00201_),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(net76),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_8 fanout76 (.A(_00194_),
    .X(net76));
 sky130_fd_sc_hd__buf_8 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(_00187_),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(_06509_),
    .X(net79));
 sky130_fd_sc_hd__buf_6 fanout8 (.A(_00568_),
    .X(net8));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(_06509_),
    .X(net80));
 sky130_fd_sc_hd__buf_6 fanout81 (.A(_00444_),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(_00444_),
    .X(net82));
 sky130_fd_sc_hd__buf_8 fanout83 (.A(_00437_),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_8 fanout84 (.A(_00437_),
    .X(net84));
 sky130_fd_sc_hd__buf_6 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_12 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_12 fanout87 (.A(_00431_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_16 fanout88 (.A(net90),
    .X(net88));
 sky130_fd_sc_hd__buf_6 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout9 (.A(_00568_),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 fanout90 (.A(_00387_),
    .X(net90));
 sky130_fd_sc_hd__buf_8 fanout91 (.A(_00329_),
    .X(net91));
 sky130_fd_sc_hd__buf_6 fanout92 (.A(_00329_),
    .X(net92));
 sky130_fd_sc_hd__buf_6 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(_00324_),
    .X(net94));
 sky130_fd_sc_hd__buf_6 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_8 fanout96 (.A(_00322_),
    .X(net96));
 sky130_fd_sc_hd__buf_8 fanout98 (.A(_00306_),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\div_shifter[1] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00015_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\div_shifter[23] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_06118_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00089_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\div_shifter[63] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_06260_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\divi2_l[3] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_05904_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\div_shifter[21] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_06116_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_00087_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\divi2_l[17] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\div_shifter[19] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_06114_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_00085_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\div_shifter[17] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_06111_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00083_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\div_shifter[18] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_06112_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\div_shifter[25] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_06121_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00019_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_00091_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\div_shifter[6] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_06099_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_00073_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\div_shifter[26] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_06122_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\div_shifter[22] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_06117_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\div_shifter[20] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_06115_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\divi2_l[5] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\div_shifter[24] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_06120_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net467),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_06106_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\div_shifter[8] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_06100_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_00074_),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 hold137 (.A(\div_counter[0] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_06261_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_00130_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00007_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\div_shifter[9] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_06102_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\div_shifter[27] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_06124_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\div_shifter[10] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_06103_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\div_shifter[5] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_06097_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_00071_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\div_res[31] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\divi2_l[23] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_06090_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_00065_),
    .X(net457));
 sky130_fd_sc_hd__buf_1 hold152 (.A(busy_l),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_06098_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\div_counter[3] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_06267_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_00133_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\div_shifter[3] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_06094_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\div_shifter[4] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00025_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_06096_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\div_shifter[12] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_06105_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(div_complete),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_00135_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\div_res[28] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_06087_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_00063_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\div_res[18] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_06075_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\divi2_l[25] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_00053_),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 hold171 (.A(net604),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_00131_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\div_res[24] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_06082_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_00059_),
    .X(net481));
 sky130_fd_sc_hd__buf_1 hold176 (.A(net492),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_05895_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\div_res[17] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_06074_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_00027_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\div_res[14] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_06069_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_00048_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\div_res[26] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_06085_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_00061_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\div_counter[2] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\div_res[8] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_06062_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\div_res[5] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\divi2_l[24] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_06060_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_00040_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net532),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_06080_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_00057_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\div_res[12] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_06067_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_00046_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\div_res[9] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_06063_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00067_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00026_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\div_res[22] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_06079_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00056_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net545),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_06070_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\div_res[10] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_06064_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\div_res[16] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_06073_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\div_res[25] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\divi2_l[29] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_06084_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\div_res[0] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_06054_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\div_res[27] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_06086_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\div_res[13] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_06068_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(net543),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_06056_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\div_res[11] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_00031_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_06066_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\div_res[21] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_06078_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_00055_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\div_res[4] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_06058_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\div_res[23] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_06081_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\div_res[6] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_06061_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\divi2_l[20] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_00041_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\div_res[30] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_06088_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_00064_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\div_res[20] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_06076_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_00054_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\div_res[3] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_06057_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\div_res[15] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_00022_),
    .X(net330));
 sky130_fd_sc_hd__buf_1 hold240 (.A(\div_shifter[32] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_06131_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\div_shifter[62] ),
    .X(net548));
 sky130_fd_sc_hd__buf_1 hold243 (.A(_06051_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\div_shifter[61] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_06253_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\div_shifter[35] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_06144_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\div_res[2] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_06055_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\divi2_l[18] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\div_shifter[34] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_06139_),
    .X(net557));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold252 (.A(\div_shifter[53] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_06222_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\div_shifter[59] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_06245_),
    .X(net561));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold256 (.A(\div_shifter[55] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_06229_),
    .X(net563));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold258 (.A(\div_shifter[47] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_06196_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_00020_),
    .X(net332));
 sky130_fd_sc_hd__buf_1 hold260 (.A(\div_shifter[49] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_06205_),
    .X(net567));
 sky130_fd_sc_hd__buf_1 hold262 (.A(\div_shifter[56] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_06233_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\div_shifter[58] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_06241_),
    .X(net571));
 sky130_fd_sc_hd__buf_1 hold266 (.A(\div_shifter[38] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_06155_),
    .X(net573));
 sky130_fd_sc_hd__buf_1 hold268 (.A(\div_shifter[40] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_06164_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\divi2_l[4] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\div_shifter[60] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_06249_),
    .X(net577));
 sky130_fd_sc_hd__buf_1 hold272 (.A(\div_shifter[41] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_06169_),
    .X(net579));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold274 (.A(\div_shifter[44] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_06182_),
    .X(net581));
 sky130_fd_sc_hd__buf_1 hold276 (.A(net607),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\div_shifter[52] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_06217_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\div_shifter[33] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_00006_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\div_shifter[51] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_06214_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\div_shifter[46] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_06191_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\div_shifter[37] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_06151_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\div_shifter[57] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\div_shifter[62] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\div_shifter[36] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\div_shifter[50] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\divi2_l[2] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_06209_),
    .X(net596));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold291 (.A(\div_shifter[43] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\div_shifter[39] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\div_shifter[54] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\div_shifter[48] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\div_shifter[45] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\div_shifter[30] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\div_res[2] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\div_counter[1] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_06265_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\divi2_l[30] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00004_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_00132_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\div_shifter[42] ),
    .X(net607));
 sky130_fd_sc_hd__buf_1 hold31 (.A(\div_counter[4] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_00134_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(divi1_sign),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_05900_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_00001_),
    .X(net341));
 sky130_fd_sc_hd__buf_1 hold36 (.A(\divi2_l[0] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_00002_),
    .X(net343));
 sky130_fd_sc_hd__buf_1 hold38 (.A(\div_shifter[31] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_00097_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00032_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\div_shifter[0] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_04454_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\div_shifter[15] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_06110_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_00082_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\divi2_l[1] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_05902_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\div_shifter[29] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_04432_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_06127_),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\divi2_l[21] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_00096_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\div_shifter[28] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_04443_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_06126_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\divi2_l[10] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_05913_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\divi2_l[7] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_05909_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\divi2_l[16] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_05920_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00023_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_00018_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\divi2_l[12] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_05915_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\divi2_l[9] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_05912_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\divi2_l[15] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_05919_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_00017_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\divi2_l[27] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_05933_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\divi2_l[28] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\divi2_l[14] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_05918_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_00016_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\divi2_l[8] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_05910_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\divi2_l[31] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_05938_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\divi2_l[6] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_05908_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\divi2_l[26] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00030_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_05932_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\divi2_l[11] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_05914_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\div_shifter[2] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_06093_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_00068_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\divi2_l[22] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_05927_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\divi2_l[19] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_05924_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\divi2_l[13] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\div_shifter[14] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_06109_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net448),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_06123_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00093_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\div_shifter[11] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_06104_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_00077_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\div_shifter[13] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_06108_),
    .X(net405));
 sky130_fd_sc_hd__buf_6 max_cap10 (.A(_00567_),
    .X(net10));
 sky130_fd_sc_hd__buf_6 max_cap110 (.A(_06505_),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 max_cap119 (.A(_06472_),
    .X(net119));
 sky130_fd_sc_hd__buf_4 max_cap128 (.A(_00320_),
    .X(net128));
 sky130_fd_sc_hd__buf_4 max_cap240 (.A(_02326_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 max_cap242 (.A(_02324_),
    .X(net242));
 sky130_fd_sc_hd__buf_6 max_cap250 (.A(_00255_),
    .X(net250));
 sky130_fd_sc_hd__buf_6 max_cap97 (.A(_00310_),
    .X(net97));
 sky130_fd_sc_hd__buf_6 max_cap99 (.A(_00300_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 wire201 (.A(_02319_),
    .X(net201));
 sky130_fd_sc_hd__buf_1 wire3 (.A(_02238_),
    .X(net3));
 sky130_fd_sc_hd__buf_1 wire4 (.A(_02639_),
    .X(net4));
 sky130_fd_sc_hd__buf_1 wire5 (.A(_02637_),
    .X(net5));
endmodule

