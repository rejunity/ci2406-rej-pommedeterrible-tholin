magic
tech sky130B
magscale 1 2
timestamp 1717285392
<< obsli1 >>
rect 1104 2159 138828 167569
<< obsm1 >>
rect 1104 2128 138888 167600
<< metal2 >>
rect 14002 169200 14058 170000
rect 41970 169200 42026 170000
rect 69938 169200 69994 170000
rect 97906 169200 97962 170000
rect 125874 169200 125930 170000
rect 5722 0 5778 800
rect 6734 0 6790 800
rect 7746 0 7802 800
rect 8758 0 8814 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11794 0 11850 800
rect 12806 0 12862 800
rect 13818 0 13874 800
rect 14830 0 14886 800
rect 15842 0 15898 800
rect 16854 0 16910 800
rect 17866 0 17922 800
rect 18878 0 18934 800
rect 19890 0 19946 800
rect 20902 0 20958 800
rect 21914 0 21970 800
rect 22926 0 22982 800
rect 23938 0 23994 800
rect 24950 0 25006 800
rect 25962 0 26018 800
rect 26974 0 27030 800
rect 27986 0 28042 800
rect 28998 0 29054 800
rect 30010 0 30066 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 33046 0 33102 800
rect 34058 0 34114 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39118 0 39174 800
rect 40130 0 40186 800
rect 41142 0 41198 800
rect 42154 0 42210 800
rect 43166 0 43222 800
rect 44178 0 44234 800
rect 45190 0 45246 800
rect 46202 0 46258 800
rect 47214 0 47270 800
rect 48226 0 48282 800
rect 49238 0 49294 800
rect 50250 0 50306 800
rect 51262 0 51318 800
rect 52274 0 52330 800
rect 53286 0 53342 800
rect 54298 0 54354 800
rect 55310 0 55366 800
rect 56322 0 56378 800
rect 57334 0 57390 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60370 0 60426 800
rect 61382 0 61438 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70490 0 70546 800
rect 71502 0 71558 800
rect 72514 0 72570 800
rect 73526 0 73582 800
rect 74538 0 74594 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77574 0 77630 800
rect 78586 0 78642 800
rect 79598 0 79654 800
rect 80610 0 80666 800
rect 81622 0 81678 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84658 0 84714 800
rect 85670 0 85726 800
rect 86682 0 86738 800
rect 87694 0 87750 800
rect 88706 0 88762 800
rect 89718 0 89774 800
rect 90730 0 90786 800
rect 91742 0 91798 800
rect 92754 0 92810 800
rect 93766 0 93822 800
rect 94778 0 94834 800
rect 95790 0 95846 800
rect 96802 0 96858 800
rect 97814 0 97870 800
rect 98826 0 98882 800
rect 99838 0 99894 800
rect 100850 0 100906 800
rect 101862 0 101918 800
rect 102874 0 102930 800
rect 103886 0 103942 800
rect 104898 0 104954 800
rect 105910 0 105966 800
rect 106922 0 106978 800
rect 107934 0 107990 800
rect 108946 0 109002 800
rect 109958 0 110014 800
rect 110970 0 111026 800
rect 111982 0 112038 800
rect 112994 0 113050 800
rect 114006 0 114062 800
rect 115018 0 115074 800
rect 116030 0 116086 800
rect 117042 0 117098 800
rect 118054 0 118110 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 121090 0 121146 800
rect 122102 0 122158 800
rect 123114 0 123170 800
rect 124126 0 124182 800
rect 125138 0 125194 800
rect 126150 0 126206 800
rect 127162 0 127218 800
rect 128174 0 128230 800
rect 129186 0 129242 800
rect 130198 0 130254 800
rect 131210 0 131266 800
rect 132222 0 132278 800
rect 133234 0 133290 800
rect 134246 0 134302 800
<< obsm2 >>
rect 1400 169144 13946 169200
rect 14114 169144 41914 169200
rect 42082 169144 69882 169200
rect 70050 169144 97850 169200
rect 98018 169144 125818 169200
rect 125986 169144 138624 169200
rect 1400 856 138624 169144
rect 1400 734 5666 856
rect 5834 734 6678 856
rect 6846 734 7690 856
rect 7858 734 8702 856
rect 8870 734 9714 856
rect 9882 734 10726 856
rect 10894 734 11738 856
rect 11906 734 12750 856
rect 12918 734 13762 856
rect 13930 734 14774 856
rect 14942 734 15786 856
rect 15954 734 16798 856
rect 16966 734 17810 856
rect 17978 734 18822 856
rect 18990 734 19834 856
rect 20002 734 20846 856
rect 21014 734 21858 856
rect 22026 734 22870 856
rect 23038 734 23882 856
rect 24050 734 24894 856
rect 25062 734 25906 856
rect 26074 734 26918 856
rect 27086 734 27930 856
rect 28098 734 28942 856
rect 29110 734 29954 856
rect 30122 734 30966 856
rect 31134 734 31978 856
rect 32146 734 32990 856
rect 33158 734 34002 856
rect 34170 734 35014 856
rect 35182 734 36026 856
rect 36194 734 37038 856
rect 37206 734 38050 856
rect 38218 734 39062 856
rect 39230 734 40074 856
rect 40242 734 41086 856
rect 41254 734 42098 856
rect 42266 734 43110 856
rect 43278 734 44122 856
rect 44290 734 45134 856
rect 45302 734 46146 856
rect 46314 734 47158 856
rect 47326 734 48170 856
rect 48338 734 49182 856
rect 49350 734 50194 856
rect 50362 734 51206 856
rect 51374 734 52218 856
rect 52386 734 53230 856
rect 53398 734 54242 856
rect 54410 734 55254 856
rect 55422 734 56266 856
rect 56434 734 57278 856
rect 57446 734 58290 856
rect 58458 734 59302 856
rect 59470 734 60314 856
rect 60482 734 61326 856
rect 61494 734 62338 856
rect 62506 734 63350 856
rect 63518 734 64362 856
rect 64530 734 65374 856
rect 65542 734 66386 856
rect 66554 734 67398 856
rect 67566 734 68410 856
rect 68578 734 69422 856
rect 69590 734 70434 856
rect 70602 734 71446 856
rect 71614 734 72458 856
rect 72626 734 73470 856
rect 73638 734 74482 856
rect 74650 734 75494 856
rect 75662 734 76506 856
rect 76674 734 77518 856
rect 77686 734 78530 856
rect 78698 734 79542 856
rect 79710 734 80554 856
rect 80722 734 81566 856
rect 81734 734 82578 856
rect 82746 734 83590 856
rect 83758 734 84602 856
rect 84770 734 85614 856
rect 85782 734 86626 856
rect 86794 734 87638 856
rect 87806 734 88650 856
rect 88818 734 89662 856
rect 89830 734 90674 856
rect 90842 734 91686 856
rect 91854 734 92698 856
rect 92866 734 93710 856
rect 93878 734 94722 856
rect 94890 734 95734 856
rect 95902 734 96746 856
rect 96914 734 97758 856
rect 97926 734 98770 856
rect 98938 734 99782 856
rect 99950 734 100794 856
rect 100962 734 101806 856
rect 101974 734 102818 856
rect 102986 734 103830 856
rect 103998 734 104842 856
rect 105010 734 105854 856
rect 106022 734 106866 856
rect 107034 734 107878 856
rect 108046 734 108890 856
rect 109058 734 109902 856
rect 110070 734 110914 856
rect 111082 734 111926 856
rect 112094 734 112938 856
rect 113106 734 113950 856
rect 114118 734 114962 856
rect 115130 734 115974 856
rect 116142 734 116986 856
rect 117154 734 117998 856
rect 118166 734 119010 856
rect 119178 734 120022 856
rect 120190 734 121034 856
rect 121202 734 122046 856
rect 122214 734 123058 856
rect 123226 734 124070 856
rect 124238 734 125082 856
rect 125250 734 126094 856
rect 126262 734 127106 856
rect 127274 734 128118 856
rect 128286 734 129130 856
rect 129298 734 130142 856
rect 130310 734 131154 856
rect 131322 734 132166 856
rect 132334 734 133178 856
rect 133346 734 134190 856
rect 134358 734 138624 856
<< metal3 >>
rect 139200 165656 140000 165776
rect 139200 159672 140000 159792
rect 0 153960 800 154080
rect 139200 153688 140000 153808
rect 0 152872 800 152992
rect 0 151784 800 151904
rect 0 150696 800 150816
rect 0 149608 800 149728
rect 0 148520 800 148640
rect 139200 147704 140000 147824
rect 0 147432 800 147552
rect 0 146344 800 146464
rect 0 145256 800 145376
rect 0 144168 800 144288
rect 0 143080 800 143200
rect 0 141992 800 142112
rect 139200 141720 140000 141840
rect 0 140904 800 141024
rect 0 139816 800 139936
rect 0 138728 800 138848
rect 0 137640 800 137760
rect 0 136552 800 136672
rect 139200 135736 140000 135856
rect 0 135464 800 135584
rect 0 134376 800 134496
rect 0 133288 800 133408
rect 0 132200 800 132320
rect 0 131112 800 131232
rect 0 130024 800 130144
rect 139200 129752 140000 129872
rect 0 128936 800 129056
rect 0 127848 800 127968
rect 0 126760 800 126880
rect 0 125672 800 125792
rect 0 124584 800 124704
rect 139200 123768 140000 123888
rect 0 123496 800 123616
rect 0 122408 800 122528
rect 0 121320 800 121440
rect 0 120232 800 120352
rect 0 119144 800 119264
rect 0 118056 800 118176
rect 139200 117784 140000 117904
rect 0 116968 800 117088
rect 0 115880 800 116000
rect 0 114792 800 114912
rect 0 113704 800 113824
rect 0 112616 800 112736
rect 139200 111800 140000 111920
rect 0 111528 800 111648
rect 0 110440 800 110560
rect 0 109352 800 109472
rect 0 108264 800 108384
rect 0 107176 800 107296
rect 0 106088 800 106208
rect 139200 105816 140000 105936
rect 0 105000 800 105120
rect 0 103912 800 104032
rect 0 102824 800 102944
rect 0 101736 800 101856
rect 0 100648 800 100768
rect 139200 99832 140000 99952
rect 0 99560 800 99680
rect 0 98472 800 98592
rect 0 97384 800 97504
rect 0 96296 800 96416
rect 0 95208 800 95328
rect 0 94120 800 94240
rect 139200 93848 140000 93968
rect 0 93032 800 93152
rect 0 91944 800 92064
rect 0 90856 800 90976
rect 0 89768 800 89888
rect 0 88680 800 88800
rect 139200 87864 140000 87984
rect 0 87592 800 87712
rect 0 86504 800 86624
rect 0 85416 800 85536
rect 0 84328 800 84448
rect 0 83240 800 83360
rect 0 82152 800 82272
rect 139200 81880 140000 82000
rect 0 81064 800 81184
rect 0 79976 800 80096
rect 0 78888 800 79008
rect 0 77800 800 77920
rect 0 76712 800 76832
rect 139200 75896 140000 76016
rect 0 75624 800 75744
rect 0 74536 800 74656
rect 0 73448 800 73568
rect 0 72360 800 72480
rect 0 71272 800 71392
rect 0 70184 800 70304
rect 139200 69912 140000 70032
rect 0 69096 800 69216
rect 0 68008 800 68128
rect 0 66920 800 67040
rect 0 65832 800 65952
rect 0 64744 800 64864
rect 139200 63928 140000 64048
rect 0 63656 800 63776
rect 0 62568 800 62688
rect 0 61480 800 61600
rect 0 60392 800 60512
rect 0 59304 800 59424
rect 0 58216 800 58336
rect 139200 57944 140000 58064
rect 0 57128 800 57248
rect 0 56040 800 56160
rect 0 54952 800 55072
rect 0 53864 800 53984
rect 0 52776 800 52896
rect 139200 51960 140000 52080
rect 0 51688 800 51808
rect 0 50600 800 50720
rect 0 49512 800 49632
rect 0 48424 800 48544
rect 0 47336 800 47456
rect 0 46248 800 46368
rect 139200 45976 140000 46096
rect 0 45160 800 45280
rect 0 44072 800 44192
rect 0 42984 800 43104
rect 0 41896 800 42016
rect 0 40808 800 40928
rect 139200 39992 140000 40112
rect 0 39720 800 39840
rect 0 38632 800 38752
rect 0 37544 800 37664
rect 0 36456 800 36576
rect 0 35368 800 35488
rect 0 34280 800 34400
rect 139200 34008 140000 34128
rect 0 33192 800 33312
rect 0 32104 800 32224
rect 0 31016 800 31136
rect 0 29928 800 30048
rect 0 28840 800 28960
rect 139200 28024 140000 28144
rect 0 27752 800 27872
rect 0 26664 800 26784
rect 0 25576 800 25696
rect 0 24488 800 24608
rect 0 23400 800 23520
rect 0 22312 800 22432
rect 139200 22040 140000 22160
rect 0 21224 800 21344
rect 0 20136 800 20256
rect 0 19048 800 19168
rect 0 17960 800 18080
rect 0 16872 800 16992
rect 139200 16056 140000 16176
rect 0 15784 800 15904
rect 139200 10072 140000 10192
rect 139200 4088 140000 4208
<< obsm3 >>
rect 614 165856 139200 167585
rect 614 165576 139120 165856
rect 614 159872 139200 165576
rect 614 159592 139120 159872
rect 614 154160 139200 159592
rect 880 153888 139200 154160
rect 880 153880 139120 153888
rect 614 153608 139120 153880
rect 614 153072 139200 153608
rect 880 152792 139200 153072
rect 614 151984 139200 152792
rect 880 151704 139200 151984
rect 614 150896 139200 151704
rect 880 150616 139200 150896
rect 614 149808 139200 150616
rect 880 149528 139200 149808
rect 614 148720 139200 149528
rect 880 148440 139200 148720
rect 614 147904 139200 148440
rect 614 147632 139120 147904
rect 880 147624 139120 147632
rect 880 147352 139200 147624
rect 614 146544 139200 147352
rect 880 146264 139200 146544
rect 614 145456 139200 146264
rect 880 145176 139200 145456
rect 614 144368 139200 145176
rect 880 144088 139200 144368
rect 614 143280 139200 144088
rect 880 143000 139200 143280
rect 614 142192 139200 143000
rect 880 141920 139200 142192
rect 880 141912 139120 141920
rect 614 141640 139120 141912
rect 614 141104 139200 141640
rect 880 140824 139200 141104
rect 614 140016 139200 140824
rect 880 139736 139200 140016
rect 614 138928 139200 139736
rect 880 138648 139200 138928
rect 614 137840 139200 138648
rect 880 137560 139200 137840
rect 614 136752 139200 137560
rect 880 136472 139200 136752
rect 614 135936 139200 136472
rect 614 135664 139120 135936
rect 880 135656 139120 135664
rect 880 135384 139200 135656
rect 614 134576 139200 135384
rect 880 134296 139200 134576
rect 614 133488 139200 134296
rect 880 133208 139200 133488
rect 614 132400 139200 133208
rect 880 132120 139200 132400
rect 614 131312 139200 132120
rect 880 131032 139200 131312
rect 614 130224 139200 131032
rect 880 129952 139200 130224
rect 880 129944 139120 129952
rect 614 129672 139120 129944
rect 614 129136 139200 129672
rect 880 128856 139200 129136
rect 614 128048 139200 128856
rect 880 127768 139200 128048
rect 614 126960 139200 127768
rect 880 126680 139200 126960
rect 614 125872 139200 126680
rect 880 125592 139200 125872
rect 614 124784 139200 125592
rect 880 124504 139200 124784
rect 614 123968 139200 124504
rect 614 123696 139120 123968
rect 880 123688 139120 123696
rect 880 123416 139200 123688
rect 614 122608 139200 123416
rect 880 122328 139200 122608
rect 614 121520 139200 122328
rect 880 121240 139200 121520
rect 614 120432 139200 121240
rect 880 120152 139200 120432
rect 614 119344 139200 120152
rect 880 119064 139200 119344
rect 614 118256 139200 119064
rect 880 117984 139200 118256
rect 880 117976 139120 117984
rect 614 117704 139120 117976
rect 614 117168 139200 117704
rect 880 116888 139200 117168
rect 614 116080 139200 116888
rect 880 115800 139200 116080
rect 614 114992 139200 115800
rect 880 114712 139200 114992
rect 614 113904 139200 114712
rect 880 113624 139200 113904
rect 614 112816 139200 113624
rect 880 112536 139200 112816
rect 614 112000 139200 112536
rect 614 111728 139120 112000
rect 880 111720 139120 111728
rect 880 111448 139200 111720
rect 614 110640 139200 111448
rect 880 110360 139200 110640
rect 614 109552 139200 110360
rect 880 109272 139200 109552
rect 614 108464 139200 109272
rect 880 108184 139200 108464
rect 614 107376 139200 108184
rect 880 107096 139200 107376
rect 614 106288 139200 107096
rect 880 106016 139200 106288
rect 880 106008 139120 106016
rect 614 105736 139120 106008
rect 614 105200 139200 105736
rect 880 104920 139200 105200
rect 614 104112 139200 104920
rect 880 103832 139200 104112
rect 614 103024 139200 103832
rect 880 102744 139200 103024
rect 614 101936 139200 102744
rect 880 101656 139200 101936
rect 614 100848 139200 101656
rect 880 100568 139200 100848
rect 614 100032 139200 100568
rect 614 99760 139120 100032
rect 880 99752 139120 99760
rect 880 99480 139200 99752
rect 614 98672 139200 99480
rect 880 98392 139200 98672
rect 614 97584 139200 98392
rect 880 97304 139200 97584
rect 614 96496 139200 97304
rect 880 96216 139200 96496
rect 614 95408 139200 96216
rect 880 95128 139200 95408
rect 614 94320 139200 95128
rect 880 94048 139200 94320
rect 880 94040 139120 94048
rect 614 93768 139120 94040
rect 614 93232 139200 93768
rect 880 92952 139200 93232
rect 614 92144 139200 92952
rect 880 91864 139200 92144
rect 614 91056 139200 91864
rect 880 90776 139200 91056
rect 614 89968 139200 90776
rect 880 89688 139200 89968
rect 614 88880 139200 89688
rect 880 88600 139200 88880
rect 614 88064 139200 88600
rect 614 87792 139120 88064
rect 880 87784 139120 87792
rect 880 87512 139200 87784
rect 614 86704 139200 87512
rect 880 86424 139200 86704
rect 614 85616 139200 86424
rect 880 85336 139200 85616
rect 614 84528 139200 85336
rect 880 84248 139200 84528
rect 614 83440 139200 84248
rect 880 83160 139200 83440
rect 614 82352 139200 83160
rect 880 82080 139200 82352
rect 880 82072 139120 82080
rect 614 81800 139120 82072
rect 614 81264 139200 81800
rect 880 80984 139200 81264
rect 614 80176 139200 80984
rect 880 79896 139200 80176
rect 614 79088 139200 79896
rect 880 78808 139200 79088
rect 614 78000 139200 78808
rect 880 77720 139200 78000
rect 614 76912 139200 77720
rect 880 76632 139200 76912
rect 614 76096 139200 76632
rect 614 75824 139120 76096
rect 880 75816 139120 75824
rect 880 75544 139200 75816
rect 614 74736 139200 75544
rect 880 74456 139200 74736
rect 614 73648 139200 74456
rect 880 73368 139200 73648
rect 614 72560 139200 73368
rect 880 72280 139200 72560
rect 614 71472 139200 72280
rect 880 71192 139200 71472
rect 614 70384 139200 71192
rect 880 70112 139200 70384
rect 880 70104 139120 70112
rect 614 69832 139120 70104
rect 614 69296 139200 69832
rect 880 69016 139200 69296
rect 614 68208 139200 69016
rect 880 67928 139200 68208
rect 614 67120 139200 67928
rect 880 66840 139200 67120
rect 614 66032 139200 66840
rect 880 65752 139200 66032
rect 614 64944 139200 65752
rect 880 64664 139200 64944
rect 614 64128 139200 64664
rect 614 63856 139120 64128
rect 880 63848 139120 63856
rect 880 63576 139200 63848
rect 614 62768 139200 63576
rect 880 62488 139200 62768
rect 614 61680 139200 62488
rect 880 61400 139200 61680
rect 614 60592 139200 61400
rect 880 60312 139200 60592
rect 614 59504 139200 60312
rect 880 59224 139200 59504
rect 614 58416 139200 59224
rect 880 58144 139200 58416
rect 880 58136 139120 58144
rect 614 57864 139120 58136
rect 614 57328 139200 57864
rect 880 57048 139200 57328
rect 614 56240 139200 57048
rect 880 55960 139200 56240
rect 614 55152 139200 55960
rect 880 54872 139200 55152
rect 614 54064 139200 54872
rect 880 53784 139200 54064
rect 614 52976 139200 53784
rect 880 52696 139200 52976
rect 614 52160 139200 52696
rect 614 51888 139120 52160
rect 880 51880 139120 51888
rect 880 51608 139200 51880
rect 614 50800 139200 51608
rect 880 50520 139200 50800
rect 614 49712 139200 50520
rect 880 49432 139200 49712
rect 614 48624 139200 49432
rect 880 48344 139200 48624
rect 614 47536 139200 48344
rect 880 47256 139200 47536
rect 614 46448 139200 47256
rect 880 46176 139200 46448
rect 880 46168 139120 46176
rect 614 45896 139120 46168
rect 614 45360 139200 45896
rect 880 45080 139200 45360
rect 614 44272 139200 45080
rect 880 43992 139200 44272
rect 614 43184 139200 43992
rect 880 42904 139200 43184
rect 614 42096 139200 42904
rect 880 41816 139200 42096
rect 614 41008 139200 41816
rect 880 40728 139200 41008
rect 614 40192 139200 40728
rect 614 39920 139120 40192
rect 880 39912 139120 39920
rect 880 39640 139200 39912
rect 614 38832 139200 39640
rect 880 38552 139200 38832
rect 614 37744 139200 38552
rect 880 37464 139200 37744
rect 614 36656 139200 37464
rect 880 36376 139200 36656
rect 614 35568 139200 36376
rect 880 35288 139200 35568
rect 614 34480 139200 35288
rect 880 34208 139200 34480
rect 880 34200 139120 34208
rect 614 33928 139120 34200
rect 614 33392 139200 33928
rect 880 33112 139200 33392
rect 614 32304 139200 33112
rect 880 32024 139200 32304
rect 614 31216 139200 32024
rect 880 30936 139200 31216
rect 614 30128 139200 30936
rect 880 29848 139200 30128
rect 614 29040 139200 29848
rect 880 28760 139200 29040
rect 614 28224 139200 28760
rect 614 27952 139120 28224
rect 880 27944 139120 27952
rect 880 27672 139200 27944
rect 614 26864 139200 27672
rect 880 26584 139200 26864
rect 614 25776 139200 26584
rect 880 25496 139200 25776
rect 614 24688 139200 25496
rect 880 24408 139200 24688
rect 614 23600 139200 24408
rect 880 23320 139200 23600
rect 614 22512 139200 23320
rect 880 22240 139200 22512
rect 880 22232 139120 22240
rect 614 21960 139120 22232
rect 614 21424 139200 21960
rect 880 21144 139200 21424
rect 614 20336 139200 21144
rect 880 20056 139200 20336
rect 614 19248 139200 20056
rect 880 18968 139200 19248
rect 614 18160 139200 18968
rect 880 17880 139200 18160
rect 614 17072 139200 17880
rect 880 16792 139200 17072
rect 614 16256 139200 16792
rect 614 15984 139120 16256
rect 880 15976 139120 15984
rect 880 15704 139200 15976
rect 614 10272 139200 15704
rect 614 9992 139120 10272
rect 614 4288 139200 9992
rect 614 4008 139120 4288
rect 614 1939 139200 4008
<< metal4 >>
rect 4208 2128 4528 167600
rect 19568 2128 19888 167600
rect 34928 2128 35248 167600
rect 50288 2128 50608 167600
rect 65648 2128 65968 167600
rect 81008 2128 81328 167600
rect 96368 2128 96688 167600
rect 111728 2128 112048 167600
rect 127088 2128 127408 167600
<< obsm4 >>
rect 2819 2048 4128 166293
rect 4608 2048 19488 166293
rect 19968 2048 34848 166293
rect 35328 2048 50208 166293
rect 50688 2048 65568 166293
rect 66048 2048 80928 166293
rect 81408 2048 96288 166293
rect 96768 2048 111648 166293
rect 112128 2048 127008 166293
rect 127488 2048 137941 166293
rect 2819 1939 137941 2048
<< labels >>
rlabel metal2 s 5722 0 5778 800 6 cache_entry[0]
port 1 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 cache_entry[100]
port 2 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 cache_entry[101]
port 3 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 cache_entry[102]
port 4 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 cache_entry[103]
port 5 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 cache_entry[104]
port 6 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 cache_entry[105]
port 7 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 cache_entry[106]
port 8 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 cache_entry[107]
port 9 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 cache_entry[108]
port 10 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 cache_entry[109]
port 11 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 cache_entry[10]
port 12 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 cache_entry[110]
port 13 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 cache_entry[111]
port 14 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 cache_entry[112]
port 15 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 cache_entry[113]
port 16 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 cache_entry[114]
port 17 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 cache_entry[115]
port 18 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 cache_entry[116]
port 19 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 cache_entry[117]
port 20 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 cache_entry[118]
port 21 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 cache_entry[119]
port 22 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 cache_entry[11]
port 23 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 cache_entry[120]
port 24 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 cache_entry[121]
port 25 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 cache_entry[122]
port 26 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 cache_entry[123]
port 27 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 cache_entry[124]
port 28 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 cache_entry[125]
port 29 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 cache_entry[126]
port 30 nsew signal output
rlabel metal2 s 134246 0 134302 800 6 cache_entry[127]
port 31 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 cache_entry[12]
port 32 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 cache_entry[13]
port 33 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 cache_entry[14]
port 34 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 cache_entry[15]
port 35 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 cache_entry[16]
port 36 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 cache_entry[17]
port 37 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 cache_entry[18]
port 38 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 cache_entry[19]
port 39 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 cache_entry[1]
port 40 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 cache_entry[20]
port 41 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 cache_entry[21]
port 42 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 cache_entry[22]
port 43 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 cache_entry[23]
port 44 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 cache_entry[24]
port 45 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 cache_entry[25]
port 46 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 cache_entry[26]
port 47 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 cache_entry[27]
port 48 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 cache_entry[28]
port 49 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 cache_entry[29]
port 50 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 cache_entry[2]
port 51 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 cache_entry[30]
port 52 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 cache_entry[31]
port 53 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 cache_entry[32]
port 54 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 cache_entry[33]
port 55 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 cache_entry[34]
port 56 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 cache_entry[35]
port 57 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 cache_entry[36]
port 58 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 cache_entry[37]
port 59 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 cache_entry[38]
port 60 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 cache_entry[39]
port 61 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 cache_entry[3]
port 62 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 cache_entry[40]
port 63 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 cache_entry[41]
port 64 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 cache_entry[42]
port 65 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 cache_entry[43]
port 66 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 cache_entry[44]
port 67 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 cache_entry[45]
port 68 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 cache_entry[46]
port 69 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 cache_entry[47]
port 70 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 cache_entry[48]
port 71 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 cache_entry[49]
port 72 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 cache_entry[4]
port 73 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 cache_entry[50]
port 74 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 cache_entry[51]
port 75 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 cache_entry[52]
port 76 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 cache_entry[53]
port 77 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 cache_entry[54]
port 78 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 cache_entry[55]
port 79 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 cache_entry[56]
port 80 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 cache_entry[57]
port 81 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 cache_entry[58]
port 82 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 cache_entry[59]
port 83 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 cache_entry[5]
port 84 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 cache_entry[60]
port 85 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 cache_entry[61]
port 86 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 cache_entry[62]
port 87 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 cache_entry[63]
port 88 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 cache_entry[64]
port 89 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 cache_entry[65]
port 90 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 cache_entry[66]
port 91 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 cache_entry[67]
port 92 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 cache_entry[68]
port 93 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 cache_entry[69]
port 94 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 cache_entry[6]
port 95 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 cache_entry[70]
port 96 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 cache_entry[71]
port 97 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 cache_entry[72]
port 98 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 cache_entry[73]
port 99 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 cache_entry[74]
port 100 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 cache_entry[75]
port 101 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 cache_entry[76]
port 102 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 cache_entry[77]
port 103 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 cache_entry[78]
port 104 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 cache_entry[79]
port 105 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 cache_entry[7]
port 106 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 cache_entry[80]
port 107 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 cache_entry[81]
port 108 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 cache_entry[82]
port 109 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 cache_entry[83]
port 110 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 cache_entry[84]
port 111 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 cache_entry[85]
port 112 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 cache_entry[86]
port 113 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 cache_entry[87]
port 114 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 cache_entry[88]
port 115 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 cache_entry[89]
port 116 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 cache_entry[8]
port 117 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 cache_entry[90]
port 118 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 cache_entry[91]
port 119 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 cache_entry[92]
port 120 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 cache_entry[93]
port 121 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 cache_entry[94]
port 122 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 cache_entry[95]
port 123 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 cache_entry[96]
port 124 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 cache_entry[97]
port 125 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 cache_entry[98]
port 126 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 cache_entry[99]
port 127 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 cache_entry[9]
port 128 nsew signal output
rlabel metal2 s 97906 169200 97962 170000 6 cache_hit
port 129 nsew signal output
rlabel metal3 s 139200 4088 140000 4208 6 curr_PC[0]
port 130 nsew signal input
rlabel metal3 s 139200 63928 140000 64048 6 curr_PC[10]
port 131 nsew signal input
rlabel metal3 s 139200 69912 140000 70032 6 curr_PC[11]
port 132 nsew signal input
rlabel metal3 s 139200 75896 140000 76016 6 curr_PC[12]
port 133 nsew signal input
rlabel metal3 s 139200 81880 140000 82000 6 curr_PC[13]
port 134 nsew signal input
rlabel metal3 s 139200 87864 140000 87984 6 curr_PC[14]
port 135 nsew signal input
rlabel metal3 s 139200 93848 140000 93968 6 curr_PC[15]
port 136 nsew signal input
rlabel metal3 s 139200 99832 140000 99952 6 curr_PC[16]
port 137 nsew signal input
rlabel metal3 s 139200 105816 140000 105936 6 curr_PC[17]
port 138 nsew signal input
rlabel metal3 s 139200 111800 140000 111920 6 curr_PC[18]
port 139 nsew signal input
rlabel metal3 s 139200 117784 140000 117904 6 curr_PC[19]
port 140 nsew signal input
rlabel metal3 s 139200 10072 140000 10192 6 curr_PC[1]
port 141 nsew signal input
rlabel metal3 s 139200 123768 140000 123888 6 curr_PC[20]
port 142 nsew signal input
rlabel metal3 s 139200 129752 140000 129872 6 curr_PC[21]
port 143 nsew signal input
rlabel metal3 s 139200 135736 140000 135856 6 curr_PC[22]
port 144 nsew signal input
rlabel metal3 s 139200 141720 140000 141840 6 curr_PC[23]
port 145 nsew signal input
rlabel metal3 s 139200 147704 140000 147824 6 curr_PC[24]
port 146 nsew signal input
rlabel metal3 s 139200 153688 140000 153808 6 curr_PC[25]
port 147 nsew signal input
rlabel metal3 s 139200 159672 140000 159792 6 curr_PC[26]
port 148 nsew signal input
rlabel metal3 s 139200 165656 140000 165776 6 curr_PC[27]
port 149 nsew signal input
rlabel metal3 s 139200 16056 140000 16176 6 curr_PC[2]
port 150 nsew signal input
rlabel metal3 s 139200 22040 140000 22160 6 curr_PC[3]
port 151 nsew signal input
rlabel metal3 s 139200 28024 140000 28144 6 curr_PC[4]
port 152 nsew signal input
rlabel metal3 s 139200 34008 140000 34128 6 curr_PC[5]
port 153 nsew signal input
rlabel metal3 s 139200 39992 140000 40112 6 curr_PC[6]
port 154 nsew signal input
rlabel metal3 s 139200 45976 140000 46096 6 curr_PC[7]
port 155 nsew signal input
rlabel metal3 s 139200 51960 140000 52080 6 curr_PC[8]
port 156 nsew signal input
rlabel metal3 s 139200 57944 140000 58064 6 curr_PC[9]
port 157 nsew signal input
rlabel metal2 s 125874 169200 125930 170000 6 entry_valid
port 158 nsew signal input
rlabel metal2 s 69938 169200 69994 170000 6 invalidate
port 159 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 new_entry[0]
port 160 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 new_entry[100]
port 161 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 new_entry[101]
port 162 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 new_entry[102]
port 163 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 new_entry[103]
port 164 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 new_entry[104]
port 165 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 new_entry[105]
port 166 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 new_entry[106]
port 167 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 new_entry[107]
port 168 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 new_entry[108]
port 169 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 new_entry[109]
port 170 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 new_entry[10]
port 171 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 new_entry[110]
port 172 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 new_entry[111]
port 173 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 new_entry[112]
port 174 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 new_entry[113]
port 175 nsew signal input
rlabel metal3 s 0 139816 800 139936 6 new_entry[114]
port 176 nsew signal input
rlabel metal3 s 0 140904 800 141024 6 new_entry[115]
port 177 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 new_entry[116]
port 178 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 new_entry[117]
port 179 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 new_entry[118]
port 180 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 new_entry[119]
port 181 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 new_entry[11]
port 182 nsew signal input
rlabel metal3 s 0 146344 800 146464 6 new_entry[120]
port 183 nsew signal input
rlabel metal3 s 0 147432 800 147552 6 new_entry[121]
port 184 nsew signal input
rlabel metal3 s 0 148520 800 148640 6 new_entry[122]
port 185 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 new_entry[123]
port 186 nsew signal input
rlabel metal3 s 0 150696 800 150816 6 new_entry[124]
port 187 nsew signal input
rlabel metal3 s 0 151784 800 151904 6 new_entry[125]
port 188 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 new_entry[126]
port 189 nsew signal input
rlabel metal3 s 0 153960 800 154080 6 new_entry[127]
port 190 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 new_entry[12]
port 191 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 new_entry[13]
port 192 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 new_entry[14]
port 193 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 new_entry[15]
port 194 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 new_entry[16]
port 195 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 new_entry[17]
port 196 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 new_entry[18]
port 197 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 new_entry[19]
port 198 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 new_entry[1]
port 199 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 new_entry[20]
port 200 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 new_entry[21]
port 201 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 new_entry[22]
port 202 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 new_entry[23]
port 203 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 new_entry[24]
port 204 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 new_entry[25]
port 205 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 new_entry[26]
port 206 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 new_entry[27]
port 207 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 new_entry[28]
port 208 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 new_entry[29]
port 209 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 new_entry[2]
port 210 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 new_entry[30]
port 211 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 new_entry[31]
port 212 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 new_entry[32]
port 213 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 new_entry[33]
port 214 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 new_entry[34]
port 215 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 new_entry[35]
port 216 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 new_entry[36]
port 217 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 new_entry[37]
port 218 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 new_entry[38]
port 219 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 new_entry[39]
port 220 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 new_entry[3]
port 221 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 new_entry[40]
port 222 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 new_entry[41]
port 223 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 new_entry[42]
port 224 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 new_entry[43]
port 225 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 new_entry[44]
port 226 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 new_entry[45]
port 227 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 new_entry[46]
port 228 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 new_entry[47]
port 229 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 new_entry[48]
port 230 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 new_entry[49]
port 231 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 new_entry[4]
port 232 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 new_entry[50]
port 233 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 new_entry[51]
port 234 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 new_entry[52]
port 235 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 new_entry[53]
port 236 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 new_entry[54]
port 237 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 new_entry[55]
port 238 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 new_entry[56]
port 239 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 new_entry[57]
port 240 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 new_entry[58]
port 241 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 new_entry[59]
port 242 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 new_entry[5]
port 243 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 new_entry[60]
port 244 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 new_entry[61]
port 245 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 new_entry[62]
port 246 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 new_entry[63]
port 247 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 new_entry[64]
port 248 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 new_entry[65]
port 249 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 new_entry[66]
port 250 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 new_entry[67]
port 251 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 new_entry[68]
port 252 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 new_entry[69]
port 253 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 new_entry[6]
port 254 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 new_entry[70]
port 255 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 new_entry[71]
port 256 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 new_entry[72]
port 257 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 new_entry[73]
port 258 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 new_entry[74]
port 259 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 new_entry[75]
port 260 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 new_entry[76]
port 261 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 new_entry[77]
port 262 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 new_entry[78]
port 263 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 new_entry[79]
port 264 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 new_entry[7]
port 265 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 new_entry[80]
port 266 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 new_entry[81]
port 267 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 new_entry[82]
port 268 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 new_entry[83]
port 269 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 new_entry[84]
port 270 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 new_entry[85]
port 271 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 new_entry[86]
port 272 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 new_entry[87]
port 273 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 new_entry[88]
port 274 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 new_entry[89]
port 275 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 new_entry[8]
port 276 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 new_entry[90]
port 277 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 new_entry[91]
port 278 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 new_entry[92]
port 279 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 new_entry[93]
port 280 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 new_entry[94]
port 281 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 new_entry[95]
port 282 nsew signal input
rlabel metal3 s 0 120232 800 120352 6 new_entry[96]
port 283 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 new_entry[97]
port 284 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 new_entry[98]
port 285 nsew signal input
rlabel metal3 s 0 123496 800 123616 6 new_entry[99]
port 286 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 new_entry[9]
port 287 nsew signal input
rlabel metal2 s 41970 169200 42026 170000 6 rst
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 167600 6 vccd1
port 289 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 167600 6 vccd1
port 289 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 167600 6 vccd1
port 289 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 167600 6 vccd1
port 289 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 167600 6 vccd1
port 289 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 167600 6 vssd1
port 290 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 167600 6 vssd1
port 290 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 167600 6 vssd1
port 290 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 167600 6 vssd1
port 290 nsew ground bidirectional
rlabel metal2 s 14002 169200 14058 170000 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 140000 170000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 73956902
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/icache/runs/24_06_01_22_42/results/signoff/icache.magic.gds
string GDS_START 588570
<< end >>

