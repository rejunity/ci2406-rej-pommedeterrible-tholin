// This is the unpowered netlist.
module execution_unit (busy,
    dest_pred_val,
    is_load,
    is_store,
    pred_val,
    rst,
    sign_extend,
    take_branch,
    wb_clk_i,
    curr_PC,
    dest_idx,
    dest_mask,
    dest_pred,
    dest_val,
    instruction,
    loadstore_address,
    loadstore_dest,
    loadstore_size,
    new_PC,
    pred_idx,
    reg1_idx,
    reg1_val,
    reg2_idx,
    reg2_val);
 output busy;
 output dest_pred_val;
 output is_load;
 output is_store;
 input pred_val;
 input rst;
 output sign_extend;
 output take_branch;
 input wb_clk_i;
 input [27:0] curr_PC;
 output [4:0] dest_idx;
 output [1:0] dest_mask;
 output [2:0] dest_pred;
 output [31:0] dest_val;
 input [41:0] instruction;
 output [31:0] loadstore_address;
 output [4:0] loadstore_dest;
 output [1:0] loadstore_size;
 output [27:0] new_PC;
 output [2:0] pred_idx;
 output [4:0] reg1_idx;
 input [31:0] reg1_val;
 output [4:0] reg2_idx;
 input [31:0] reg2_val;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire busy_l;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire div_complete;
 wire \div_counter[0] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_res[0] ;
 wire \div_res[10] ;
 wire \div_res[11] ;
 wire \div_res[12] ;
 wire \div_res[13] ;
 wire \div_res[14] ;
 wire \div_res[15] ;
 wire \div_res[16] ;
 wire \div_res[17] ;
 wire \div_res[18] ;
 wire \div_res[19] ;
 wire \div_res[1] ;
 wire \div_res[20] ;
 wire \div_res[21] ;
 wire \div_res[22] ;
 wire \div_res[23] ;
 wire \div_res[24] ;
 wire \div_res[25] ;
 wire \div_res[26] ;
 wire \div_res[27] ;
 wire \div_res[28] ;
 wire \div_res[29] ;
 wire \div_res[2] ;
 wire \div_res[30] ;
 wire \div_res[31] ;
 wire \div_res[3] ;
 wire \div_res[4] ;
 wire \div_res[5] ;
 wire \div_res[6] ;
 wire \div_res[7] ;
 wire \div_res[8] ;
 wire \div_res[9] ;
 wire \div_shifter[0] ;
 wire \div_shifter[10] ;
 wire \div_shifter[11] ;
 wire \div_shifter[12] ;
 wire \div_shifter[13] ;
 wire \div_shifter[14] ;
 wire \div_shifter[15] ;
 wire \div_shifter[16] ;
 wire \div_shifter[17] ;
 wire \div_shifter[18] ;
 wire \div_shifter[19] ;
 wire \div_shifter[1] ;
 wire \div_shifter[20] ;
 wire \div_shifter[21] ;
 wire \div_shifter[22] ;
 wire \div_shifter[23] ;
 wire \div_shifter[24] ;
 wire \div_shifter[25] ;
 wire \div_shifter[26] ;
 wire \div_shifter[27] ;
 wire \div_shifter[28] ;
 wire \div_shifter[29] ;
 wire \div_shifter[2] ;
 wire \div_shifter[30] ;
 wire \div_shifter[31] ;
 wire \div_shifter[32] ;
 wire \div_shifter[33] ;
 wire \div_shifter[34] ;
 wire \div_shifter[35] ;
 wire \div_shifter[36] ;
 wire \div_shifter[37] ;
 wire \div_shifter[38] ;
 wire \div_shifter[39] ;
 wire \div_shifter[3] ;
 wire \div_shifter[40] ;
 wire \div_shifter[41] ;
 wire \div_shifter[42] ;
 wire \div_shifter[43] ;
 wire \div_shifter[44] ;
 wire \div_shifter[45] ;
 wire \div_shifter[46] ;
 wire \div_shifter[47] ;
 wire \div_shifter[48] ;
 wire \div_shifter[49] ;
 wire \div_shifter[4] ;
 wire \div_shifter[50] ;
 wire \div_shifter[51] ;
 wire \div_shifter[52] ;
 wire \div_shifter[53] ;
 wire \div_shifter[54] ;
 wire \div_shifter[55] ;
 wire \div_shifter[56] ;
 wire \div_shifter[57] ;
 wire \div_shifter[58] ;
 wire \div_shifter[59] ;
 wire \div_shifter[5] ;
 wire \div_shifter[60] ;
 wire \div_shifter[61] ;
 wire \div_shifter[62] ;
 wire \div_shifter[63] ;
 wire \div_shifter[6] ;
 wire \div_shifter[7] ;
 wire \div_shifter[8] ;
 wire \div_shifter[9] ;
 wire divi1_sign;
 wire \divi2_l[0] ;
 wire \divi2_l[10] ;
 wire \divi2_l[11] ;
 wire \divi2_l[12] ;
 wire \divi2_l[13] ;
 wire \divi2_l[14] ;
 wire \divi2_l[15] ;
 wire \divi2_l[16] ;
 wire \divi2_l[17] ;
 wire \divi2_l[18] ;
 wire \divi2_l[19] ;
 wire \divi2_l[1] ;
 wire \divi2_l[20] ;
 wire \divi2_l[21] ;
 wire \divi2_l[22] ;
 wire \divi2_l[23] ;
 wire \divi2_l[24] ;
 wire \divi2_l[25] ;
 wire \divi2_l[26] ;
 wire \divi2_l[27] ;
 wire \divi2_l[28] ;
 wire \divi2_l[29] ;
 wire \divi2_l[2] ;
 wire \divi2_l[30] ;
 wire \divi2_l[31] ;
 wire \divi2_l[3] ;
 wire \divi2_l[4] ;
 wire \divi2_l[5] ;
 wire \divi2_l[6] ;
 wire \divi2_l[7] ;
 wire \divi2_l[8] ;
 wire \divi2_l[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(reg1_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(reg1_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(reg2_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(reg2_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(reg2_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(reg2_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(reg2_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(reg2_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(reg2_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(reg2_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(reg2_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(reg2_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(instruction[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(instruction[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(pred_val));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(pred_val));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(pred_val));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(reg1_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(reg1_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(reg1_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(reg1_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(reg1_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(reg1_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(reg1_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(reg1_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(reg2_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(reg1_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(reg1_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(reg1_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06572__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__B (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__B (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__A2 (.DIODE(_04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__B (.DIODE(_04709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A2_N (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__B (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__A_N (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__B (.DIODE(_04785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__B (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__B (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06615__B (.DIODE(_04861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__B1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__B (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__B (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__B (.DIODE(_04948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__A_N (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__B (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06629__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__A2_N (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__A_N (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06632__B (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__B (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__A2_N (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__A_N (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__B (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__B (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06644__B (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__B (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__B (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06653__A_N (.DIODE(_05275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06654__B (.DIODE(_05275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06657__B (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__A2_N (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__B1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__A2_N (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__B1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__B (.DIODE(_05426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__B (.DIODE(_05426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__B (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06673__A_N (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__B (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__B (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__B (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__A_N (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__B (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__B (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__B (.DIODE(_05658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__B (.DIODE(_05658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__B (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__B (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06698__A_N (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__B (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__B (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__B (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A_N (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__B (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__A2 (.DIODE(_04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__A_N (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06711__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__A3 (.DIODE(_04785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__B1 (.DIODE(_05898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__A_N (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__B (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__B (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A3 (.DIODE(_04861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A_N (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__B (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06724__B (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__A3 (.DIODE(_04948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__B1 (.DIODE(_05988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__A_N (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__B (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__B (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06733__A3 (.DIODE(_04709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06733__B1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06734__A_N (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__B (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__B (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__A3 (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A_N (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__B (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__B (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A3 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__B1 (.DIODE(_06144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__A_N (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__B (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__B (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__B (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__A3 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__B1 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__A_N (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06755__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__A3 (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__B1 (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A_N (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__B (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A3 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__B1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__A_N (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__B (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__B (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__B (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06770__C1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__C_N (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06773__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06773__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__B (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__B (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A3 (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__B1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__A3 (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__B1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A3 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__B1 (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__A3 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__B1 (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A3 (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__B1 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__A3 (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__B1 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A3 (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__B1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__A3 (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__B1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__B (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__B (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__B (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__A2 (.DIODE(_05275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__B (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__B (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06840__B (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__B (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__B (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__B1 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__B (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__B (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__B (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__A2 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__B1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__B (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__B (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__B (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__S (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__B (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__C (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__C (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__C (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__D (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__C (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__D (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__B (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__B (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__B1 (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A1 (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__A1 (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__A (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__A2 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__A2 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__A3 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A1 (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A2 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__C (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__C (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__B (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A1 (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A2 (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A3 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__B2 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__D (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__B (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__B (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__A_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__C (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__B (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__B1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__C1 (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__B (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__C (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__C1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__C (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__B (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__B (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__B (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__B1 (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__C1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A_N (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__C (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__B (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__C_N (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__A (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A4 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A1 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A2 (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__B (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__C (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__B1_N (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__C_N (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__B1 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__B (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A2 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A2 (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A2 (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__A (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__B (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__A1 (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__A (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__C_N (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__B (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__B (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__B (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__A (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__S (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__A (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__B (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__B (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__A (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__B (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A (.DIODE(_05275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__C (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__D (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__A1 (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__A (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A1 (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B2 (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__A (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A1 (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A2 (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__C1 (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__A1 (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__C1 (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__B (.DIODE(_00244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A1_N (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A2_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__B2 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A1 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A1 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A2 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(_05275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__S (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__B1 (.DIODE(_05658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A1 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B2 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A1 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A2 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__B1 (.DIODE(_05426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(_05426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__C (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__A1 (.DIODE(_05426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__A2 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__C1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A2 (.DIODE(_00224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__C1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A2 (.DIODE(_00350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__B1_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A2 (.DIODE(_00350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__B1_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B (.DIODE(_00350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A_N (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__B (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A2 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__B1 (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07354__A (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__B1 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__B (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B2 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B2 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A1 (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07436__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B1 (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A1 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B1 (.DIODE(_00167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B2 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A2 (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__B (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__C (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__C_N (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A2 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B2 (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__A0 (.DIODE(_00595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__A1 (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__B2 (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__A (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07734__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A1 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A2 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A2 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A3 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__B (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A1 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A2 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__B (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A1 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__B (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A2 (.DIODE(_01130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__C (.DIODE(_01130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08321__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A2 (.DIODE(_01482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__C (.DIODE(_01482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__B1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__A (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A_N (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__B1 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__A2 (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__B2 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A2 (.DIODE(_06526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__B2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08722__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A2 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A3 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__C1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__S (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__S (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__S (.DIODE(_02175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__S (.DIODE(_02175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__S (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__S (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A2 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A1 (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A2 (.DIODE(_02258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B1 (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09177__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A2 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A3 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__A0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__S (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__B1 (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09197__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__B2 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A2 (.DIODE(_00244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__B1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__B1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A (.DIODE(_06526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__A (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A1 (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__B1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__C_N (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__B (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A1 (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__B1 (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__B2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__A2 (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__B1 (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B1 (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A2 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A1 (.DIODE(_06526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__B1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A2 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__B2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__B (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B1 (.DIODE(_02627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__B1 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A2 (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__A (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__B (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__B (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__B (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__S (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A2 (.DIODE(_02760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A3 (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__B1 (.DIODE(_02258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__A2 (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A1 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A2 (.DIODE(_02760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__B2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__A2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__A2_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__B2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__B (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__B (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__B (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__B (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__B1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__B1 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09834__D (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__C1 (.DIODE(_02924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A2 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A3 (.DIODE(_02930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A2 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__B1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09852__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A2 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A3 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A1 (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B2 (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__B1 (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__B1 (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__B2 (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__B2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__B1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__C1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__A1 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10012__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__B (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__B (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__B1 (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A2 (.DIODE(_00178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A (.DIODE(_03086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B (.DIODE(_03178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A (.DIODE(_03086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__B (.DIODE(_03178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A (.DIODE(_03086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__B (.DIODE(_03178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__B1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B1 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__C1 (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A2 (.DIODE(_00244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__B2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A1 (.DIODE(_00178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__B (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__B (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__B (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A1_N (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A2_N (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__A1 (.DIODE(_00178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__A (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__B (.DIODE(_03405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__B (.DIODE(_03405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__B (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__B (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__B1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__S (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__A1_N (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__A2_N (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__C1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__B2 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A1 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A3 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B2 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A2 (.DIODE(_00244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A_N (.DIODE(_03572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__B (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A_N (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B (.DIODE(_03572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__B (.DIODE(_03572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__B1 (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A3 (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__C1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__S (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A1 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__B1 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__C1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__B1 (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__B2 (.DIODE(_03606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__B1 (.DIODE(_03612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A2 (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__B2 (.DIODE(_00178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__A (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__B (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__B (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__C1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A1 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__B1 (.DIODE(_03729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A1 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__S (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__C_N (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__D_N (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A1 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__A (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__C1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A1_N (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A2_N (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__C1 (.DIODE(_03852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__B (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A1 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B1 (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A1 (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B1_N (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__A3 (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__B1 (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__A2 (.DIODE(_03950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A2 (.DIODE(_03950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__B1 (.DIODE(_03975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__B2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__A1 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__B2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__B1 (.DIODE(_03983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A3 (.DIODE(_03950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A2 (.DIODE(_00244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B1_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__B1_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__B (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__A2 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__A2 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__B (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A (.DIODE(_05955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__B (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__C1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__C1 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A2 (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A2 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A3 (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__B2 (.DIODE(_00178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11065__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11065__B (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11105__A2 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11105__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A2 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__C1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__B (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A1 (.DIODE(_05907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__C1 (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A2 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__B1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__S (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A2 (.DIODE(_03950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A3 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A4 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A1 (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A2 (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__C1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__B (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A1 (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__C1 (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__B1 (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A1_N (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A2_N (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__B2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__C1 (.DIODE(_04326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__B (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__C (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A1 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__B1 (.DIODE(_04404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__C (.DIODE(_04404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11326__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11330__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__S (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A (.DIODE(_05799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A2 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A1 (.DIODE(_02258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B1 (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A1_N (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A2 (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B1 (.DIODE(_04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__B1 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__B (.DIODE(_04404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__A (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__A2 (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A1 (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A2 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A1 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__B1 (.DIODE(_02258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__B1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__A2 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A3 (.DIODE(_04549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A2 (.DIODE(_04404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A3 (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__B (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A1_N (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A2_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__A (.DIODE(_04614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__B (.DIODE(_04614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__A2 (.DIODE(_04614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__B (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__C1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A1 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A2 (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__B1 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__B2 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__C1 (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11574__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A3 (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__11624__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__B (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__C1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__C1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__A (.DIODE(_04404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__B (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__C (.DIODE(_04614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__B (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__C (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__B1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__S (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__B (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__C1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__A1 (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__B2 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11737__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11816__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__B2 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A2 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__B (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__B (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__C1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__A_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__B (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__C1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__C1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__S (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__B (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__C1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A1 (.DIODE(_05275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__B (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__A2_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12042__S (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A0 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A2 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__B1 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A1 (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__A (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__B (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A2 (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__S (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__B1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__S (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__B1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__A0 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__S (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A1 (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__C1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A2 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__B1 (.DIODE(_05417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A1 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__A1 (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__B1 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A3 (.DIODE(_00350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A4 (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__C1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__B1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__A2 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__C1 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A2 (.DIODE(_02760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B2 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__C1 (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A1 (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__C1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12350__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__D_N (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A1 (.DIODE(_04883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__C1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A2 (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__S (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__B1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A1 (.DIODE(_02175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__C1 (.DIODE(_05581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__A1 (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__A2 (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__C1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__A (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__B (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__B1 (.DIODE(_02258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__A2 (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A2 (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A3 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__C1 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__B2 (.DIODE(_02243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__A1 (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A1 (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A2 (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__C1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__A0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A (.DIODE(_04600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__A (.DIODE(_04600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__A (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__S (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__A (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__A (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__A (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__A (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__A (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__A (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__A (.DIODE(_04709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A (.DIODE(_04709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A (.DIODE(_04948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A (.DIODE(_04948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A (.DIODE(_04861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A (.DIODE(_04861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A (.DIODE(_04785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A (.DIODE(_04785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__B (.DIODE(_04600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__B (.DIODE(_04600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__B (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__B (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__B (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__B (.DIODE(_05716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__B (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__B (.DIODE(_05629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__B (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__B (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__B (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__B (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__B (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__B (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__B (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__B (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__B (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__B (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__B (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__B (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__B (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__B (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__B (.DIODE(_04709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__B (.DIODE(_04709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__B (.DIODE(_04948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__B (.DIODE(_04948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__B (.DIODE(_04861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__B (.DIODE(_04861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__B (.DIODE(_04785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A2 (.DIODE(_04785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A1 (.DIODE(_06526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A1 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A1 (.DIODE(_00510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12915__B (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__A (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__A1 (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A1 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A1 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A1 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__A1 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__C1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A1 (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A1 (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__A1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A1 (.DIODE(_00350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A1 (.DIODE(_00456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__B1 (.DIODE(_00595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__B2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A0 (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13242__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13247__C1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__13248__B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(_02175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(_02175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(_00178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(_04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(_04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(_04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(_04471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(_04471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(_04471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(_00595_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(_00167_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(_00166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold260_A (.DIODE(\div_shifter[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew214_A (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap151_A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap261_A (.DIODE(_00213_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_98 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06566_ (.A(net605),
    .Y(_04340_));
 sky130_fd_sc_hd__inv_2 _06567_ (.A(net392),
    .Y(_04351_));
 sky130_fd_sc_hd__inv_2 _06568_ (.A(net382),
    .Y(_04362_));
 sky130_fd_sc_hd__inv_2 _06569_ (.A(net389),
    .Y(_04373_));
 sky130_fd_sc_hd__inv_2 _06570_ (.A(net367),
    .Y(_04384_));
 sky130_fd_sc_hd__inv_2 _06571_ (.A(net606),
    .Y(_04395_));
 sky130_fd_sc_hd__inv_2 _06572_ (.A(net278),
    .Y(_04406_));
 sky130_fd_sc_hd__inv_2 _06573_ (.A(instruction[3]),
    .Y(_04417_));
 sky130_fd_sc_hd__inv_2 _06574_ (.A(net308),
    .Y(_04428_));
 sky130_fd_sc_hd__inv_2 _06575_ (.A(instruction[41]),
    .Y(_04439_));
 sky130_fd_sc_hd__inv_2 _06576_ (.A(reg1_val[29]),
    .Y(_04449_));
 sky130_fd_sc_hd__inv_2 _06577_ (.A(net310),
    .Y(_04460_));
 sky130_fd_sc_hd__inv_2 _06578_ (.A(rst),
    .Y(_04471_));
 sky130_fd_sc_hd__or4bb_4 _06579_ (.A(instruction[0]),
    .B(instruction[1]),
    .C_N(instruction[2]),
    .D_N(pred_val),
    .X(_04482_));
 sky130_fd_sc_hd__nor2_8 _06580_ (.A(instruction[3]),
    .B(_04482_),
    .Y(is_load));
 sky130_fd_sc_hd__nor2_8 _06581_ (.A(_04417_),
    .B(_04482_),
    .Y(is_store));
 sky130_fd_sc_hd__and3b_1 _06582_ (.A_N(instruction[0]),
    .B(pred_val),
    .C(instruction[1]),
    .X(_04513_));
 sky130_fd_sc_hd__and4bb_4 _06583_ (.A_N(instruction[0]),
    .B_N(instruction[2]),
    .C(instruction[1]),
    .D(pred_val),
    .X(_04524_));
 sky130_fd_sc_hd__or4bb_1 _06584_ (.A(instruction[0]),
    .B(instruction[2]),
    .C_N(instruction[1]),
    .D_N(pred_val),
    .X(_04535_));
 sky130_fd_sc_hd__and2_1 _06585_ (.A(reg2_val[31]),
    .B(net290),
    .X(_04546_));
 sky130_fd_sc_hd__o31a_1 _06586_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(pred_val),
    .X(_04556_));
 sky130_fd_sc_hd__o311a_4 _06587_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[41]),
    .C1(pred_val),
    .X(_04567_));
 sky130_fd_sc_hd__and4bb_2 _06588_ (.A_N(instruction[1]),
    .B_N(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04578_));
 sky130_fd_sc_hd__or4bb_4 _06589_ (.A(instruction[1]),
    .B(instruction[2]),
    .C_N(instruction[0]),
    .D_N(pred_val),
    .X(_04589_));
 sky130_fd_sc_hd__and2_4 _06590_ (.A(instruction[25]),
    .B(net287),
    .X(_04600_));
 sky130_fd_sc_hd__o211a_1 _06591_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .X(_04611_));
 sky130_fd_sc_hd__o211ai_1 _06592_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .Y(_04622_));
 sky130_fd_sc_hd__a21o_1 _06593_ (.A1(instruction[41]),
    .A2(_04578_),
    .B1(_04611_),
    .X(_04633_));
 sky130_fd_sc_hd__a21oi_4 _06594_ (.A1(instruction[41]),
    .A2(_04578_),
    .B1(_04611_),
    .Y(_04644_));
 sky130_fd_sc_hd__a221o_1 _06595_ (.A1(instruction[24]),
    .A2(_04567_),
    .B1(_04578_),
    .B2(instruction[41]),
    .C1(_04611_),
    .X(_04654_));
 sky130_fd_sc_hd__nand2_2 _06596_ (.A(_04524_),
    .B(_04654_),
    .Y(_04665_));
 sky130_fd_sc_hd__o21ba_2 _06597_ (.A1(_04439_),
    .A2(_04665_),
    .B1_N(_04546_),
    .X(_04676_));
 sky130_fd_sc_hd__a31o_4 _06598_ (.A1(instruction[41]),
    .A2(_04524_),
    .A3(_04654_),
    .B1(_04546_),
    .X(_04687_));
 sky130_fd_sc_hd__xor2_4 _06599_ (.A(reg1_val[31]),
    .B(_04687_),
    .X(_04698_));
 sky130_fd_sc_hd__and2_4 _06600_ (.A(instruction[37]),
    .B(net288),
    .X(_04709_));
 sky130_fd_sc_hd__nor2_1 _06601_ (.A(_04644_),
    .B(_04709_),
    .Y(_04720_));
 sky130_fd_sc_hd__o2bb2a_4 _06602_ (.A1_N(reg2_val[27]),
    .A2_N(net290),
    .B1(_04665_),
    .B2(_04720_),
    .X(_04731_));
 sky130_fd_sc_hd__nand2b_1 _06603_ (.A_N(reg1_val[27]),
    .B(_04731_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2b_2 _06604_ (.A_N(_04731_),
    .B(reg1_val[27]),
    .Y(_04753_));
 sky130_fd_sc_hd__inv_2 _06605_ (.A(_04753_),
    .Y(_04763_));
 sky130_fd_sc_hd__nand2_1 _06606_ (.A(_04742_),
    .B(_04753_),
    .Y(_04774_));
 sky130_fd_sc_hd__and2_4 _06607_ (.A(instruction[40]),
    .B(net288),
    .X(_04785_));
 sky130_fd_sc_hd__nor2_1 _06608_ (.A(net270),
    .B(_04785_),
    .Y(_04796_));
 sky130_fd_sc_hd__a2bb2o_2 _06609_ (.A1_N(_04796_),
    .A2_N(net245),
    .B1(net289),
    .B2(reg2_val[30]),
    .X(_04807_));
 sky130_fd_sc_hd__inv_2 _06610_ (.A(_04807_),
    .Y(_04818_));
 sky130_fd_sc_hd__and2_1 _06611_ (.A(reg1_val[30]),
    .B(_04807_),
    .X(_04829_));
 sky130_fd_sc_hd__nor2_1 _06612_ (.A(reg1_val[30]),
    .B(_04807_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_2 _06613_ (.A(_04829_),
    .B(_04840_),
    .Y(_04851_));
 sky130_fd_sc_hd__and2_4 _06614_ (.A(instruction[39]),
    .B(net288),
    .X(_04861_));
 sky130_fd_sc_hd__nor2_1 _06615_ (.A(_04644_),
    .B(_04861_),
    .Y(_04872_));
 sky130_fd_sc_hd__a2bb2o_4 _06616_ (.A1_N(_04872_),
    .A2_N(net245),
    .B1(net290),
    .B2(reg2_val[29]),
    .X(_04883_));
 sky130_fd_sc_hd__nand2_1 _06617_ (.A(reg1_val[29]),
    .B(_04883_),
    .Y(_04894_));
 sky130_fd_sc_hd__or2_1 _06618_ (.A(reg1_val[29]),
    .B(_04883_),
    .X(_04905_));
 sky130_fd_sc_hd__inv_2 _06619_ (.A(_04905_),
    .Y(_04916_));
 sky130_fd_sc_hd__and2_1 _06620_ (.A(_04894_),
    .B(_04905_),
    .X(_04927_));
 sky130_fd_sc_hd__nand2_1 _06621_ (.A(_04894_),
    .B(_04905_),
    .Y(_04938_));
 sky130_fd_sc_hd__and2_4 _06622_ (.A(instruction[38]),
    .B(net288),
    .X(_04948_));
 sky130_fd_sc_hd__nor2_1 _06623_ (.A(net270),
    .B(_04948_),
    .Y(_04959_));
 sky130_fd_sc_hd__o2bb2a_4 _06624_ (.A1_N(reg2_val[28]),
    .A2_N(net289),
    .B1(net245),
    .B2(_04959_),
    .X(_04970_));
 sky130_fd_sc_hd__and2b_1 _06625_ (.A_N(_04970_),
    .B(reg1_val[28]),
    .X(_04981_));
 sky130_fd_sc_hd__nand2b_1 _06626_ (.A_N(reg1_val[28]),
    .B(_04970_),
    .Y(_04992_));
 sky130_fd_sc_hd__and2b_1 _06627_ (.A_N(_04981_),
    .B(_04992_),
    .X(_05003_));
 sky130_fd_sc_hd__and2_4 _06628_ (.A(instruction[35]),
    .B(net288),
    .X(_05014_));
 sky130_fd_sc_hd__nor2_1 _06629_ (.A(_04644_),
    .B(_05014_),
    .Y(_05025_));
 sky130_fd_sc_hd__o2bb2a_2 _06630_ (.A1_N(reg2_val[25]),
    .A2_N(net290),
    .B1(net245),
    .B2(_05025_),
    .X(_05035_));
 sky130_fd_sc_hd__and2b_1 _06631_ (.A_N(_05035_),
    .B(reg1_val[25]),
    .X(_05046_));
 sky130_fd_sc_hd__and2b_1 _06632_ (.A_N(reg1_val[25]),
    .B(_05035_),
    .X(_05057_));
 sky130_fd_sc_hd__or2_2 _06633_ (.A(_05046_),
    .B(_05057_),
    .X(_05068_));
 sky130_fd_sc_hd__and2_4 _06634_ (.A(instruction[36]),
    .B(net288),
    .X(_05079_));
 sky130_fd_sc_hd__nor2_1 _06635_ (.A(_04644_),
    .B(_05079_),
    .Y(_05090_));
 sky130_fd_sc_hd__o2bb2a_2 _06636_ (.A1_N(reg2_val[26]),
    .A2_N(net290),
    .B1(_04665_),
    .B2(_05090_),
    .X(_05101_));
 sky130_fd_sc_hd__and2b_1 _06637_ (.A_N(_05101_),
    .B(reg1_val[26]),
    .X(_05112_));
 sky130_fd_sc_hd__and2b_1 _06638_ (.A_N(reg1_val[26]),
    .B(_05101_),
    .X(_05122_));
 sky130_fd_sc_hd__or2_2 _06639_ (.A(_05112_),
    .B(_05122_),
    .X(_05133_));
 sky130_fd_sc_hd__and2_4 _06640_ (.A(instruction[34]),
    .B(net287),
    .X(_05144_));
 sky130_fd_sc_hd__nor2_1 _06641_ (.A(net271),
    .B(_05144_),
    .Y(_05155_));
 sky130_fd_sc_hd__o2bb2a_1 _06642_ (.A1_N(reg2_val[24]),
    .A2_N(net289),
    .B1(net245),
    .B2(_05155_),
    .X(_05166_));
 sky130_fd_sc_hd__a2bb2o_2 _06643_ (.A1_N(_05155_),
    .A2_N(net245),
    .B1(net289),
    .B2(reg2_val[24]),
    .X(_05177_));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(reg1_val[24]),
    .B(_05177_),
    .Y(_05188_));
 sky130_fd_sc_hd__or2_1 _06645_ (.A(reg1_val[24]),
    .B(_05177_),
    .X(_05199_));
 sky130_fd_sc_hd__nand2_2 _06646_ (.A(_05188_),
    .B(_05199_),
    .Y(_05209_));
 sky130_fd_sc_hd__or3_1 _06647_ (.A(_04851_),
    .B(_04927_),
    .C(_05003_),
    .X(_05220_));
 sky130_fd_sc_hd__and4b_1 _06648_ (.A_N(_04698_),
    .B(_05068_),
    .C(_05133_),
    .D(_05209_),
    .X(_05231_));
 sky130_fd_sc_hd__nand3b_1 _06649_ (.A_N(_05220_),
    .B(_05231_),
    .C(_04774_),
    .Y(_05242_));
 sky130_fd_sc_hd__and2_4 _06650_ (.A(instruction[33]),
    .B(net287),
    .X(_05253_));
 sky130_fd_sc_hd__nor2_1 _06651_ (.A(net271),
    .B(_05253_),
    .Y(_05264_));
 sky130_fd_sc_hd__o2bb2a_2 _06652_ (.A1_N(reg2_val[23]),
    .A2_N(net289),
    .B1(net245),
    .B2(_05264_),
    .X(_05275_));
 sky130_fd_sc_hd__and2b_1 _06653_ (.A_N(_05275_),
    .B(reg1_val[23]),
    .X(_05286_));
 sky130_fd_sc_hd__and2b_1 _06654_ (.A_N(reg1_val[23]),
    .B(_05275_),
    .X(_05296_));
 sky130_fd_sc_hd__nor2_1 _06655_ (.A(_05286_),
    .B(_05296_),
    .Y(_05307_));
 sky130_fd_sc_hd__and2_4 _06656_ (.A(instruction[32]),
    .B(net287),
    .X(_05318_));
 sky130_fd_sc_hd__nor2_1 _06657_ (.A(net272),
    .B(_05318_),
    .Y(_05329_));
 sky130_fd_sc_hd__o2bb2a_1 _06658_ (.A1_N(reg2_val[22]),
    .A2_N(net290),
    .B1(net245),
    .B2(_05329_),
    .X(_05340_));
 sky130_fd_sc_hd__a2bb2o_2 _06659_ (.A1_N(_05329_),
    .A2_N(net245),
    .B1(net290),
    .B2(reg2_val[22]),
    .X(_05351_));
 sky130_fd_sc_hd__and2_1 _06660_ (.A(reg1_val[22]),
    .B(_05351_),
    .X(_05361_));
 sky130_fd_sc_hd__nor2_1 _06661_ (.A(reg1_val[22]),
    .B(_05351_),
    .Y(_05372_));
 sky130_fd_sc_hd__nor2_2 _06662_ (.A(_05361_),
    .B(_05372_),
    .Y(_05383_));
 sky130_fd_sc_hd__and2_4 _06663_ (.A(instruction[30]),
    .B(net287),
    .X(_05394_));
 sky130_fd_sc_hd__nor2_1 _06664_ (.A(net272),
    .B(_05394_),
    .Y(_05405_));
 sky130_fd_sc_hd__o2bb2a_2 _06665_ (.A1_N(reg2_val[20]),
    .A2_N(net290),
    .B1(net245),
    .B2(_05405_),
    .X(_05416_));
 sky130_fd_sc_hd__a2bb2o_2 _06666_ (.A1_N(_05405_),
    .A2_N(net245),
    .B1(net290),
    .B2(reg2_val[20]),
    .X(_05426_));
 sky130_fd_sc_hd__and2_1 _06667_ (.A(reg1_val[20]),
    .B(_05426_),
    .X(_05437_));
 sky130_fd_sc_hd__nor2_1 _06668_ (.A(reg1_val[20]),
    .B(_05426_),
    .Y(_05448_));
 sky130_fd_sc_hd__nor2_2 _06669_ (.A(_05437_),
    .B(_05448_),
    .Y(_05459_));
 sky130_fd_sc_hd__o311a_4 _06670_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[31]),
    .C1(pred_val),
    .X(_05470_));
 sky130_fd_sc_hd__nor2_1 _06671_ (.A(net270),
    .B(_05470_),
    .Y(_05480_));
 sky130_fd_sc_hd__o2bb2a_4 _06672_ (.A1_N(reg2_val[21]),
    .A2_N(net289),
    .B1(net245),
    .B2(_05480_),
    .X(_05491_));
 sky130_fd_sc_hd__and2b_1 _06673_ (.A_N(_05491_),
    .B(reg1_val[21]),
    .X(_05502_));
 sky130_fd_sc_hd__and2b_1 _06674_ (.A_N(reg1_val[21]),
    .B(_05491_),
    .X(_05513_));
 sky130_fd_sc_hd__nor2_2 _06675_ (.A(_05502_),
    .B(_05513_),
    .Y(_05524_));
 sky130_fd_sc_hd__or4_1 _06676_ (.A(_05307_),
    .B(_05383_),
    .C(_05459_),
    .D(_05524_),
    .X(_05534_));
 sky130_fd_sc_hd__and2_4 _06677_ (.A(instruction[29]),
    .B(net287),
    .X(_05545_));
 sky130_fd_sc_hd__nor2_1 _06678_ (.A(net271),
    .B(_05545_),
    .Y(_05556_));
 sky130_fd_sc_hd__o2bb2a_2 _06679_ (.A1_N(reg2_val[19]),
    .A2_N(net289),
    .B1(_04665_),
    .B2(_05556_),
    .X(_05567_));
 sky130_fd_sc_hd__and2_1 _06680_ (.A(reg1_val[19]),
    .B(_05567_),
    .X(_05578_));
 sky130_fd_sc_hd__and2b_1 _06681_ (.A_N(_05567_),
    .B(reg1_val[19]),
    .X(_05588_));
 sky130_fd_sc_hd__and2b_1 _06682_ (.A_N(reg1_val[19]),
    .B(_05567_),
    .X(_05599_));
 sky130_fd_sc_hd__nor2_1 _06683_ (.A(_05588_),
    .B(_05599_),
    .Y(_05610_));
 sky130_fd_sc_hd__inv_2 _06684_ (.A(_05610_),
    .Y(_05620_));
 sky130_fd_sc_hd__and2_4 _06685_ (.A(instruction[28]),
    .B(net287),
    .X(_05629_));
 sky130_fd_sc_hd__nor2_1 _06686_ (.A(net272),
    .B(_05629_),
    .Y(_05639_));
 sky130_fd_sc_hd__o2bb2a_2 _06687_ (.A1_N(reg2_val[18]),
    .A2_N(net289),
    .B1(net245),
    .B2(_05639_),
    .X(_05649_));
 sky130_fd_sc_hd__a2bb2o_2 _06688_ (.A1_N(_05639_),
    .A2_N(net245),
    .B1(net289),
    .B2(reg2_val[18]),
    .X(_05658_));
 sky130_fd_sc_hd__and2_1 _06689_ (.A(reg1_val[18]),
    .B(_05649_),
    .X(_05668_));
 sky130_fd_sc_hd__and2_1 _06690_ (.A(reg1_val[18]),
    .B(_05658_),
    .X(_05677_));
 sky130_fd_sc_hd__nor2_1 _06691_ (.A(reg1_val[18]),
    .B(_05658_),
    .Y(_05687_));
 sky130_fd_sc_hd__nor2_1 _06692_ (.A(_05677_),
    .B(_05687_),
    .Y(_05696_));
 sky130_fd_sc_hd__or2_1 _06693_ (.A(_05677_),
    .B(_05687_),
    .X(_05706_));
 sky130_fd_sc_hd__and2_4 _06694_ (.A(instruction[27]),
    .B(net287),
    .X(_05716_));
 sky130_fd_sc_hd__nor2_1 _06695_ (.A(net271),
    .B(_05716_),
    .Y(_05725_));
 sky130_fd_sc_hd__o2bb2a_4 _06696_ (.A1_N(reg2_val[17]),
    .A2_N(net289),
    .B1(net245),
    .B2(_05725_),
    .X(_05734_));
 sky130_fd_sc_hd__and2_1 _06697_ (.A(reg1_val[17]),
    .B(_05734_),
    .X(_05744_));
 sky130_fd_sc_hd__and2b_1 _06698_ (.A_N(_05734_),
    .B(reg1_val[17]),
    .X(_05754_));
 sky130_fd_sc_hd__nand2b_1 _06699_ (.A_N(reg1_val[17]),
    .B(_05734_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2b_1 _06700_ (.A_N(_05754_),
    .B(_05763_),
    .Y(_05772_));
 sky130_fd_sc_hd__o311a_4 _06701_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[26]),
    .C1(pred_val),
    .X(_05781_));
 sky130_fd_sc_hd__nor2_1 _06702_ (.A(net270),
    .B(_05781_),
    .Y(_05790_));
 sky130_fd_sc_hd__o2bb2a_4 _06703_ (.A1_N(reg2_val[16]),
    .A2_N(net289),
    .B1(net245),
    .B2(_05790_),
    .X(_05799_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(reg1_val[16]),
    .B(_05799_),
    .Y(_05808_));
 sky130_fd_sc_hd__and2b_1 _06705_ (.A_N(_05799_),
    .B(reg1_val[16]),
    .X(_05817_));
 sky130_fd_sc_hd__nand2b_1 _06706_ (.A_N(reg1_val[16]),
    .B(_05799_),
    .Y(_05826_));
 sky130_fd_sc_hd__and2b_1 _06707_ (.A_N(_05817_),
    .B(_05826_),
    .X(_05835_));
 sky130_fd_sc_hd__and2_1 _06708_ (.A(reg2_val[15]),
    .B(net289),
    .X(_05844_));
 sky130_fd_sc_hd__a31o_4 _06709_ (.A1(net292),
    .A2(_04567_),
    .A3(net272),
    .B1(_05844_),
    .X(_05854_));
 sky130_fd_sc_hd__and2b_1 _06710_ (.A_N(_05854_),
    .B(reg1_val[15]),
    .X(_05863_));
 sky130_fd_sc_hd__and2_1 _06711_ (.A(reg1_val[15]),
    .B(_05854_),
    .X(_05872_));
 sky130_fd_sc_hd__nor2_1 _06712_ (.A(reg1_val[15]),
    .B(_05854_),
    .Y(_05880_));
 sky130_fd_sc_hd__nor2_1 _06713_ (.A(_05872_),
    .B(_05880_),
    .Y(_05889_));
 sky130_fd_sc_hd__and2_1 _06714_ (.A(reg2_val[14]),
    .B(net291),
    .X(_05898_));
 sky130_fd_sc_hd__a31o_4 _06715_ (.A1(net292),
    .A2(net272),
    .A3(_04785_),
    .B1(_05898_),
    .X(_05907_));
 sky130_fd_sc_hd__nand2b_1 _06716_ (.A_N(_05907_),
    .B(reg1_val[14]),
    .Y(_05916_));
 sky130_fd_sc_hd__and2_1 _06717_ (.A(reg1_val[14]),
    .B(_05907_),
    .X(_05925_));
 sky130_fd_sc_hd__nor2_1 _06718_ (.A(reg1_val[14]),
    .B(_05907_),
    .Y(_05934_));
 sky130_fd_sc_hd__nor2_1 _06719_ (.A(_05925_),
    .B(_05934_),
    .Y(_05943_));
 sky130_fd_sc_hd__and2_1 _06720_ (.A(reg2_val[13]),
    .B(net289),
    .X(_05949_));
 sky130_fd_sc_hd__a31o_4 _06721_ (.A1(net292),
    .A2(net270),
    .A3(_04861_),
    .B1(_05949_),
    .X(_05955_));
 sky130_fd_sc_hd__nand2b_1 _06722_ (.A_N(_05955_),
    .B(reg1_val[13]),
    .Y(_05961_));
 sky130_fd_sc_hd__and2_1 _06723_ (.A(reg1_val[13]),
    .B(_05955_),
    .X(_05967_));
 sky130_fd_sc_hd__nor2_1 _06724_ (.A(reg1_val[13]),
    .B(_05955_),
    .Y(_05973_));
 sky130_fd_sc_hd__nor2_1 _06725_ (.A(_05967_),
    .B(_05973_),
    .Y(_05979_));
 sky130_fd_sc_hd__and2_1 _06726_ (.A(reg2_val[12]),
    .B(net291),
    .X(_05988_));
 sky130_fd_sc_hd__a31o_4 _06727_ (.A1(net292),
    .A2(net270),
    .A3(_04948_),
    .B1(_05988_),
    .X(_05999_));
 sky130_fd_sc_hd__nand2b_1 _06728_ (.A_N(_05999_),
    .B(reg1_val[12]),
    .Y(_06010_));
 sky130_fd_sc_hd__and2_1 _06729_ (.A(reg1_val[12]),
    .B(_05999_),
    .X(_06021_));
 sky130_fd_sc_hd__nor2_1 _06730_ (.A(reg1_val[12]),
    .B(_05999_),
    .Y(_06032_));
 sky130_fd_sc_hd__nor2_1 _06731_ (.A(_06021_),
    .B(_06032_),
    .Y(_06043_));
 sky130_fd_sc_hd__and2_1 _06732_ (.A(reg2_val[11]),
    .B(net291),
    .X(_06054_));
 sky130_fd_sc_hd__a31o_4 _06733_ (.A1(net292),
    .A2(net270),
    .A3(_04709_),
    .B1(_06054_),
    .X(_06065_));
 sky130_fd_sc_hd__and2b_1 _06734_ (.A_N(_06065_),
    .B(reg1_val[11]),
    .X(_06076_));
 sky130_fd_sc_hd__and2_1 _06735_ (.A(reg1_val[11]),
    .B(_06065_),
    .X(_06087_));
 sky130_fd_sc_hd__nor2_1 _06736_ (.A(reg1_val[11]),
    .B(_06065_),
    .Y(_06096_));
 sky130_fd_sc_hd__nor2_1 _06737_ (.A(_06087_),
    .B(_06096_),
    .Y(_06102_));
 sky130_fd_sc_hd__and2_1 _06738_ (.A(reg2_val[10]),
    .B(net291),
    .X(_06108_));
 sky130_fd_sc_hd__a31o_4 _06739_ (.A1(net292),
    .A2(net270),
    .A3(_05079_),
    .B1(_06108_),
    .X(_06114_));
 sky130_fd_sc_hd__nand2b_1 _06740_ (.A_N(_06114_),
    .B(reg1_val[10]),
    .Y(_06120_));
 sky130_fd_sc_hd__and2_1 _06741_ (.A(reg1_val[10]),
    .B(_06114_),
    .X(_06126_));
 sky130_fd_sc_hd__nor2_1 _06742_ (.A(reg1_val[10]),
    .B(_06114_),
    .Y(_06132_));
 sky130_fd_sc_hd__nor2_1 _06743_ (.A(_06126_),
    .B(_06132_),
    .Y(_06138_));
 sky130_fd_sc_hd__and2_1 _06744_ (.A(reg2_val[9]),
    .B(net291),
    .X(_06144_));
 sky130_fd_sc_hd__a31o_4 _06745_ (.A1(net292),
    .A2(net270),
    .A3(_05014_),
    .B1(_06144_),
    .X(_06150_));
 sky130_fd_sc_hd__and2b_1 _06746_ (.A_N(_06150_),
    .B(reg1_val[9]),
    .X(_06156_));
 sky130_fd_sc_hd__nor2_1 _06747_ (.A(reg1_val[9]),
    .B(_06150_),
    .Y(_06162_));
 sky130_fd_sc_hd__and2_1 _06748_ (.A(reg1_val[9]),
    .B(_06150_),
    .X(_06168_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(reg1_val[9]),
    .B(_06150_),
    .Y(_06176_));
 sky130_fd_sc_hd__or2_1 _06750_ (.A(_06162_),
    .B(_06168_),
    .X(_06185_));
 sky130_fd_sc_hd__and2_1 _06751_ (.A(reg2_val[8]),
    .B(net291),
    .X(_06193_));
 sky130_fd_sc_hd__a31o_4 _06752_ (.A1(net292),
    .A2(net270),
    .A3(_05144_),
    .B1(_06193_),
    .X(_06202_));
 sky130_fd_sc_hd__and2b_1 _06753_ (.A_N(_06202_),
    .B(reg1_val[8]),
    .X(_06211_));
 sky130_fd_sc_hd__nor2_1 _06754_ (.A(reg1_val[8]),
    .B(_06202_),
    .Y(_06220_));
 sky130_fd_sc_hd__nand2_1 _06755_ (.A(reg1_val[8]),
    .B(_06202_),
    .Y(_06229_));
 sky130_fd_sc_hd__nand2b_2 _06756_ (.A_N(_06220_),
    .B(_06229_),
    .Y(_06238_));
 sky130_fd_sc_hd__and2_1 _06757_ (.A(reg2_val[7]),
    .B(net291),
    .X(_06247_));
 sky130_fd_sc_hd__a31o_4 _06758_ (.A1(net292),
    .A2(net270),
    .A3(_05253_),
    .B1(_06247_),
    .X(_06256_));
 sky130_fd_sc_hd__and2b_1 _06759_ (.A_N(_06256_),
    .B(reg1_val[7]),
    .X(_06265_));
 sky130_fd_sc_hd__nor2_1 _06760_ (.A(reg1_val[7]),
    .B(_06256_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand2_1 _06761_ (.A(reg1_val[7]),
    .B(_06256_),
    .Y(_06282_));
 sky130_fd_sc_hd__nand2b_2 _06762_ (.A_N(_06274_),
    .B(_06282_),
    .Y(_06291_));
 sky130_fd_sc_hd__and2_1 _06763_ (.A(reg2_val[6]),
    .B(net291),
    .X(_06300_));
 sky130_fd_sc_hd__a31o_4 _06764_ (.A1(net292),
    .A2(net270),
    .A3(_05318_),
    .B1(_06300_),
    .X(_06307_));
 sky130_fd_sc_hd__nand2b_1 _06765_ (.A_N(_06307_),
    .B(reg1_val[6]),
    .Y(_06309_));
 sky130_fd_sc_hd__nor2_1 _06766_ (.A(reg1_val[6]),
    .B(_06307_),
    .Y(_06310_));
 sky130_fd_sc_hd__or2_1 _06767_ (.A(reg1_val[6]),
    .B(_06307_),
    .X(_06311_));
 sky130_fd_sc_hd__and2_1 _06768_ (.A(reg1_val[6]),
    .B(_06307_),
    .X(_06312_));
 sky130_fd_sc_hd__nor2_1 _06769_ (.A(_06310_),
    .B(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__o2111a_2 _06770_ (.A1(_04439_),
    .A2(_04589_),
    .B1(_04622_),
    .C1(_05470_),
    .D1(_04524_),
    .X(_06314_));
 sky130_fd_sc_hd__or3b_1 _06771_ (.A(net290),
    .B(_04633_),
    .C_N(_05470_),
    .X(_06315_));
 sky130_fd_sc_hd__a21oi_4 _06772_ (.A1(reg2_val[5]),
    .A2(net289),
    .B1(net269),
    .Y(_06316_));
 sky130_fd_sc_hd__a21o_2 _06773_ (.A1(reg2_val[5]),
    .A2(net290),
    .B1(net269),
    .X(_06317_));
 sky130_fd_sc_hd__and2_1 _06774_ (.A(reg1_val[5]),
    .B(_06316_),
    .X(_06318_));
 sky130_fd_sc_hd__nor2_1 _06775_ (.A(reg1_val[5]),
    .B(_06317_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand2_1 _06776_ (.A(reg1_val[5]),
    .B(_06317_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2b_1 _06777_ (.A_N(_06319_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__and2_2 _06778_ (.A(reg2_val[4]),
    .B(net291),
    .X(_06322_));
 sky130_fd_sc_hd__a31o_1 _06779_ (.A1(net292),
    .A2(net272),
    .A3(_05394_),
    .B1(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__a31oi_4 _06780_ (.A1(net292),
    .A2(net272),
    .A3(_05394_),
    .B1(_06322_),
    .Y(_06324_));
 sky130_fd_sc_hd__and2_1 _06781_ (.A(reg1_val[4]),
    .B(net239),
    .X(_06325_));
 sky130_fd_sc_hd__nor2_1 _06782_ (.A(reg1_val[4]),
    .B(net241),
    .Y(_06326_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(reg1_val[4]),
    .B(net241),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2b_2 _06784_ (.A_N(_06326_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__and2_2 _06785_ (.A(reg2_val[3]),
    .B(net291),
    .X(_06329_));
 sky130_fd_sc_hd__a31oi_4 _06786_ (.A1(_04524_),
    .A2(net271),
    .A3(_05545_),
    .B1(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__a31o_1 _06787_ (.A1(_04524_),
    .A2(net271),
    .A3(_05545_),
    .B1(_06329_),
    .X(_06331_));
 sky130_fd_sc_hd__and2_1 _06788_ (.A(reg1_val[3]),
    .B(net238),
    .X(_06332_));
 sky130_fd_sc_hd__nor2_1 _06789_ (.A(reg1_val[3]),
    .B(net236),
    .Y(_06333_));
 sky130_fd_sc_hd__nand2_1 _06790_ (.A(reg1_val[3]),
    .B(net236),
    .Y(_06334_));
 sky130_fd_sc_hd__nand2b_2 _06791_ (.A_N(_06333_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__and2_2 _06792_ (.A(reg2_val[2]),
    .B(net291),
    .X(_06336_));
 sky130_fd_sc_hd__a31oi_4 _06793_ (.A1(net292),
    .A2(net271),
    .A3(_05629_),
    .B1(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__a31o_1 _06794_ (.A1(_04524_),
    .A2(net271),
    .A3(_05629_),
    .B1(_06336_),
    .X(_06338_));
 sky130_fd_sc_hd__and2_1 _06795_ (.A(reg1_val[2]),
    .B(net235),
    .X(_06339_));
 sky130_fd_sc_hd__nor2_1 _06796_ (.A(reg1_val[2]),
    .B(net233),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_1 _06797_ (.A(reg1_val[2]),
    .B(net233),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2b_2 _06798_ (.A_N(_06340_),
    .B(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__and2_2 _06799_ (.A(reg2_val[1]),
    .B(net291),
    .X(_06343_));
 sky130_fd_sc_hd__a31oi_2 _06800_ (.A1(net292),
    .A2(net270),
    .A3(_05716_),
    .B1(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__a31o_2 _06801_ (.A1(net292),
    .A2(net270),
    .A3(_05716_),
    .B1(_06343_),
    .X(_06345_));
 sky130_fd_sc_hd__and2_1 _06802_ (.A(net307),
    .B(net231),
    .X(_06346_));
 sky130_fd_sc_hd__or2_1 _06803_ (.A(net307),
    .B(net230),
    .X(_06347_));
 sky130_fd_sc_hd__xnor2_2 _06804_ (.A(net307),
    .B(net230),
    .Y(_06348_));
 sky130_fd_sc_hd__and2_1 _06805_ (.A(net292),
    .B(_05781_),
    .X(_06349_));
 sky130_fd_sc_hd__a22oi_1 _06806_ (.A1(reg2_val[0]),
    .A2(net289),
    .B1(net270),
    .B2(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__a22o_1 _06807_ (.A1(reg2_val[0]),
    .A2(net289),
    .B1(net270),
    .B2(_06349_),
    .X(_06351_));
 sky130_fd_sc_hd__nand2_1 _06808_ (.A(net306),
    .B(net224),
    .Y(_06352_));
 sky130_fd_sc_hd__a21o_1 _06809_ (.A1(_06348_),
    .A2(_06352_),
    .B1(_06346_),
    .X(_06353_));
 sky130_fd_sc_hd__a21o_1 _06810_ (.A1(_06342_),
    .A2(_06353_),
    .B1(_06339_),
    .X(_06354_));
 sky130_fd_sc_hd__a21o_1 _06811_ (.A1(_06335_),
    .A2(_06354_),
    .B1(_06332_),
    .X(_06355_));
 sky130_fd_sc_hd__a21o_1 _06812_ (.A1(_06328_),
    .A2(_06355_),
    .B1(_06325_),
    .X(_06356_));
 sky130_fd_sc_hd__a21oi_1 _06813_ (.A1(_06321_),
    .A2(_06356_),
    .B1(_06318_),
    .Y(_06357_));
 sky130_fd_sc_hd__o21ai_1 _06814_ (.A1(_06313_),
    .A2(_06357_),
    .B1(_06309_),
    .Y(_06358_));
 sky130_fd_sc_hd__a21o_1 _06815_ (.A1(_06291_),
    .A2(_06358_),
    .B1(_06265_),
    .X(_06359_));
 sky130_fd_sc_hd__a21o_1 _06816_ (.A1(_06238_),
    .A2(_06359_),
    .B1(_06211_),
    .X(_06360_));
 sky130_fd_sc_hd__a21oi_1 _06817_ (.A1(_06185_),
    .A2(_06360_),
    .B1(_06156_),
    .Y(_06361_));
 sky130_fd_sc_hd__o21a_1 _06818_ (.A1(_06138_),
    .A2(_06361_),
    .B1(_06120_),
    .X(_06362_));
 sky130_fd_sc_hd__o21ba_1 _06819_ (.A1(_06102_),
    .A2(_06362_),
    .B1_N(_06076_),
    .X(_06363_));
 sky130_fd_sc_hd__o21a_1 _06820_ (.A1(_06043_),
    .A2(_06363_),
    .B1(_06010_),
    .X(_06364_));
 sky130_fd_sc_hd__o21a_1 _06821_ (.A1(_05979_),
    .A2(_06364_),
    .B1(_05961_),
    .X(_06365_));
 sky130_fd_sc_hd__o21a_1 _06822_ (.A1(_05943_),
    .A2(_06365_),
    .B1(_05916_),
    .X(_06366_));
 sky130_fd_sc_hd__o21ba_1 _06823_ (.A1(_05889_),
    .A2(_06366_),
    .B1_N(_05863_),
    .X(_06367_));
 sky130_fd_sc_hd__o21ai_1 _06824_ (.A1(_05835_),
    .A2(_06367_),
    .B1(_05808_),
    .Y(_06368_));
 sky130_fd_sc_hd__a21o_1 _06825_ (.A1(_05772_),
    .A2(_06368_),
    .B1(_05744_),
    .X(_06369_));
 sky130_fd_sc_hd__a21o_1 _06826_ (.A1(_05706_),
    .A2(_06369_),
    .B1(_05668_),
    .X(_06370_));
 sky130_fd_sc_hd__a21oi_1 _06827_ (.A1(_05620_),
    .A2(_06370_),
    .B1(_05578_),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2_1 _06828_ (.A(reg1_val[22]),
    .B(_05340_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2_1 _06829_ (.A(reg1_val[21]),
    .B(_05491_),
    .Y(_06373_));
 sky130_fd_sc_hd__nand2_1 _06830_ (.A(reg1_val[20]),
    .B(_05416_),
    .Y(_06374_));
 sky130_fd_sc_hd__or2_1 _06831_ (.A(_05524_),
    .B(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__a21o_1 _06832_ (.A1(_06373_),
    .A2(_06375_),
    .B1(_05383_),
    .X(_06376_));
 sky130_fd_sc_hd__a21oi_1 _06833_ (.A1(_06372_),
    .A2(_06376_),
    .B1(_05307_),
    .Y(_06377_));
 sky130_fd_sc_hd__a21oi_1 _06834_ (.A1(reg1_val[23]),
    .A2(_05275_),
    .B1(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__o21ai_1 _06835_ (.A1(_05534_),
    .A2(_06371_),
    .B1(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__and2b_1 _06836_ (.A_N(_05242_),
    .B(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__nand2_1 _06837_ (.A(reg1_val[30]),
    .B(_04818_),
    .Y(_06381_));
 sky130_fd_sc_hd__nor2_1 _06838_ (.A(_04449_),
    .B(_04883_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _06839_ (.A(reg1_val[28]),
    .B(_04970_),
    .Y(_06383_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(reg1_val[27]),
    .B(_04731_),
    .Y(_06384_));
 sky130_fd_sc_hd__and2_1 _06841_ (.A(reg1_val[26]),
    .B(_05101_),
    .X(_06385_));
 sky130_fd_sc_hd__and2_1 _06842_ (.A(reg1_val[25]),
    .B(_05035_),
    .X(_06386_));
 sky130_fd_sc_hd__and2_1 _06843_ (.A(reg1_val[24]),
    .B(_05166_),
    .X(_06387_));
 sky130_fd_sc_hd__a21o_1 _06844_ (.A1(_05068_),
    .A2(_06387_),
    .B1(_06386_),
    .X(_06388_));
 sky130_fd_sc_hd__a21o_1 _06845_ (.A1(_05133_),
    .A2(_06388_),
    .B1(_06385_),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _06846_ (.A(_04774_),
    .B(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__a21o_1 _06847_ (.A1(_06384_),
    .A2(_06390_),
    .B1(_05003_),
    .X(_06391_));
 sky130_fd_sc_hd__a21oi_1 _06848_ (.A1(_06383_),
    .A2(_06391_),
    .B1(_04927_),
    .Y(_06392_));
 sky130_fd_sc_hd__o21ba_1 _06849_ (.A1(_06382_),
    .A2(_06392_),
    .B1_N(_04851_),
    .X(_06393_));
 sky130_fd_sc_hd__a21oi_1 _06850_ (.A1(reg1_val[30]),
    .A2(_04818_),
    .B1(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__nor2_1 _06851_ (.A(_04698_),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand2_1 _06852_ (.A(reg1_val[31]),
    .B(_04676_),
    .Y(_06396_));
 sky130_fd_sc_hd__or4b_1 _06853_ (.A(instruction[6]),
    .B(_06380_),
    .C(_06395_),
    .D_N(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__a21o_1 _06854_ (.A1(_05209_),
    .A2(_06379_),
    .B1(_06387_),
    .X(_06398_));
 sky130_fd_sc_hd__a21o_1 _06855_ (.A1(_05068_),
    .A2(_06398_),
    .B1(_06386_),
    .X(_06399_));
 sky130_fd_sc_hd__a21o_1 _06856_ (.A1(_05133_),
    .A2(_06399_),
    .B1(_06385_),
    .X(_06400_));
 sky130_fd_sc_hd__a21boi_1 _06857_ (.A1(_04774_),
    .A2(_06400_),
    .B1_N(_06384_),
    .Y(_06401_));
 sky130_fd_sc_hd__o21ai_1 _06858_ (.A1(_05003_),
    .A2(_06401_),
    .B1(_06383_),
    .Y(_06402_));
 sky130_fd_sc_hd__a21oi_1 _06859_ (.A1(_04938_),
    .A2(_06402_),
    .B1(_06382_),
    .Y(_06403_));
 sky130_fd_sc_hd__o21ai_1 _06860_ (.A1(_04851_),
    .A2(_06403_),
    .B1(_06381_),
    .Y(_06404_));
 sky130_fd_sc_hd__o21ai_1 _06861_ (.A1(_04698_),
    .A2(_06404_),
    .B1(_06396_),
    .Y(_06405_));
 sky130_fd_sc_hd__a21boi_1 _06862_ (.A1(instruction[6]),
    .A2(_06405_),
    .B1_N(_06397_),
    .Y(_06406_));
 sky130_fd_sc_hd__or2_4 _06863_ (.A(instruction[3]),
    .B(instruction[4]),
    .X(_06407_));
 sky130_fd_sc_hd__nor2_2 _06864_ (.A(net306),
    .B(net228),
    .Y(_06408_));
 sky130_fd_sc_hd__nor2_1 _06865_ (.A(net308),
    .B(net224),
    .Y(_06409_));
 sky130_fd_sc_hd__or3b_1 _06866_ (.A(_05610_),
    .B(_05696_),
    .C_N(_05772_),
    .X(_06410_));
 sky130_fd_sc_hd__nand2_1 _06867_ (.A(_06185_),
    .B(_06291_),
    .Y(_06411_));
 sky130_fd_sc_hd__or4_1 _06868_ (.A(_05889_),
    .B(_05943_),
    .C(_05979_),
    .D(_06043_),
    .X(_06412_));
 sky130_fd_sc_hd__or4_1 _06869_ (.A(_06102_),
    .B(_06138_),
    .C(_06411_),
    .D(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__and4b_1 _06870_ (.A_N(_06313_),
    .B(_06321_),
    .C(_06328_),
    .D(_06335_),
    .X(_06414_));
 sky130_fd_sc_hd__o2111a_1 _06871_ (.A1(_06408_),
    .A2(_06409_),
    .B1(_06238_),
    .C1(_06342_),
    .D1(_06348_),
    .X(_06415_));
 sky130_fd_sc_hd__nand2_1 _06872_ (.A(_06414_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__or4_1 _06873_ (.A(_05835_),
    .B(_06410_),
    .C(_06413_),
    .D(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__or3_1 _06874_ (.A(_05242_),
    .B(_05534_),
    .C(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__mux2_1 _06875_ (.A0(_06418_),
    .A1(_04698_),
    .S(instruction[6]),
    .X(_06419_));
 sky130_fd_sc_hd__nand2_2 _06876_ (.A(instruction[3]),
    .B(instruction[4]),
    .Y(_06420_));
 sky130_fd_sc_hd__o22a_1 _06877_ (.A1(_06407_),
    .A2(_06419_),
    .B1(_06420_),
    .B2(_06418_),
    .X(_06421_));
 sky130_fd_sc_hd__or2_2 _06878_ (.A(_04417_),
    .B(instruction[4]),
    .X(_06422_));
 sky130_fd_sc_hd__o21a_1 _06879_ (.A1(_04417_),
    .A2(_06406_),
    .B1(_06421_),
    .X(_06423_));
 sky130_fd_sc_hd__xnor2_4 _06880_ (.A(instruction[5]),
    .B(_06423_),
    .Y(dest_pred_val));
 sky130_fd_sc_hd__and2_4 _06881_ (.A(instruction[2]),
    .B(_04513_),
    .X(_06424_));
 sky130_fd_sc_hd__nand2_2 _06882_ (.A(instruction[2]),
    .B(_04513_),
    .Y(_06425_));
 sky130_fd_sc_hd__and4b_4 _06883_ (.A_N(instruction[1]),
    .B(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_06426_));
 sky130_fd_sc_hd__nand4b_4 _06884_ (.A_N(instruction[1]),
    .B(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .Y(_06427_));
 sky130_fd_sc_hd__a21o_4 _06885_ (.A1(dest_pred_val),
    .A2(_06426_),
    .B1(_06424_),
    .X(take_branch));
 sky130_fd_sc_hd__nand2b_4 _06886_ (.A_N(instruction[5]),
    .B(instruction[6]),
    .Y(_06428_));
 sky130_fd_sc_hd__a21oi_2 _06887_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(instruction[4]),
    .Y(_06429_));
 sky130_fd_sc_hd__a221oi_4 _06888_ (.A1(net290),
    .A2(_04589_),
    .B1(_06428_),
    .B2(instruction[4]),
    .C1(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__a221o_1 _06889_ (.A1(net290),
    .A2(_04589_),
    .B1(_06428_),
    .B2(instruction[4]),
    .C1(_06429_),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_4 _06890_ (.A(net280),
    .B(_06430_),
    .Y(_06432_));
 sky130_fd_sc_hd__nand2_1 _06891_ (.A(net274),
    .B(_06431_),
    .Y(_06433_));
 sky130_fd_sc_hd__nor2_8 _06892_ (.A(div_complete),
    .B(net222),
    .Y(busy));
 sky130_fd_sc_hd__and4b_4 _06893_ (.A_N(instruction[2]),
    .B(instruction[1]),
    .C(pred_val),
    .D(instruction[0]),
    .X(_06434_));
 sky130_fd_sc_hd__and2_4 _06894_ (.A(instruction[11]),
    .B(_06434_),
    .X(dest_pred[0]));
 sky130_fd_sc_hd__and2_4 _06895_ (.A(instruction[12]),
    .B(_06434_),
    .X(dest_pred[1]));
 sky130_fd_sc_hd__and2_4 _06896_ (.A(instruction[13]),
    .B(_06434_),
    .X(dest_pred[2]));
 sky130_fd_sc_hd__or2_2 _06897_ (.A(_04513_),
    .B(_04578_),
    .X(_06435_));
 sky130_fd_sc_hd__and2_4 _06898_ (.A(instruction[11]),
    .B(_06435_),
    .X(dest_idx[0]));
 sky130_fd_sc_hd__and2_4 _06899_ (.A(instruction[12]),
    .B(_06435_),
    .X(dest_idx[1]));
 sky130_fd_sc_hd__and2_4 _06900_ (.A(instruction[13]),
    .B(_06435_),
    .X(dest_idx[2]));
 sky130_fd_sc_hd__and2_4 _06901_ (.A(instruction[14]),
    .B(_06435_),
    .X(dest_idx[3]));
 sky130_fd_sc_hd__and2_4 _06902_ (.A(instruction[15]),
    .B(_06435_),
    .X(dest_idx[4]));
 sky130_fd_sc_hd__or2_1 _06903_ (.A(instruction[18]),
    .B(_06426_),
    .X(_06436_));
 sky130_fd_sc_hd__o211a_4 _06904_ (.A1(instruction[11]),
    .A2(_06427_),
    .B1(_06436_),
    .C1(net287),
    .X(reg1_idx[0]));
 sky130_fd_sc_hd__or2_1 _06905_ (.A(instruction[19]),
    .B(_06426_),
    .X(_06437_));
 sky130_fd_sc_hd__o211a_4 _06906_ (.A1(instruction[12]),
    .A2(_06427_),
    .B1(_06437_),
    .C1(net287),
    .X(reg1_idx[1]));
 sky130_fd_sc_hd__or2_1 _06907_ (.A(instruction[20]),
    .B(_06426_),
    .X(_06438_));
 sky130_fd_sc_hd__o211a_4 _06908_ (.A1(instruction[13]),
    .A2(_06427_),
    .B1(_06438_),
    .C1(net287),
    .X(reg1_idx[2]));
 sky130_fd_sc_hd__or2_1 _06909_ (.A(instruction[21]),
    .B(_06426_),
    .X(_06439_));
 sky130_fd_sc_hd__o211a_4 _06910_ (.A1(instruction[14]),
    .A2(_06427_),
    .B1(_06439_),
    .C1(net288),
    .X(reg1_idx[3]));
 sky130_fd_sc_hd__or2_1 _06911_ (.A(instruction[22]),
    .B(_06426_),
    .X(_06440_));
 sky130_fd_sc_hd__o211a_4 _06912_ (.A1(instruction[15]),
    .A2(_06427_),
    .B1(_06440_),
    .C1(net288),
    .X(reg1_idx[4]));
 sky130_fd_sc_hd__or2_1 _06913_ (.A(instruction[25]),
    .B(_06426_),
    .X(_06441_));
 sky130_fd_sc_hd__o211a_4 _06914_ (.A1(instruction[18]),
    .A2(_06427_),
    .B1(_06441_),
    .C1(net287),
    .X(reg2_idx[0]));
 sky130_fd_sc_hd__or2_1 _06915_ (.A(instruction[26]),
    .B(_06426_),
    .X(_06442_));
 sky130_fd_sc_hd__o211a_4 _06916_ (.A1(instruction[19]),
    .A2(_06427_),
    .B1(_06442_),
    .C1(net287),
    .X(reg2_idx[1]));
 sky130_fd_sc_hd__or2_1 _06917_ (.A(instruction[27]),
    .B(_06426_),
    .X(_06443_));
 sky130_fd_sc_hd__o211a_4 _06918_ (.A1(instruction[20]),
    .A2(_06427_),
    .B1(_06443_),
    .C1(net287),
    .X(reg2_idx[2]));
 sky130_fd_sc_hd__or2_1 _06919_ (.A(instruction[28]),
    .B(_06426_),
    .X(_06444_));
 sky130_fd_sc_hd__o211a_4 _06920_ (.A1(instruction[21]),
    .A2(_06427_),
    .B1(_06444_),
    .C1(net287),
    .X(reg2_idx[3]));
 sky130_fd_sc_hd__or2_1 _06921_ (.A(instruction[29]),
    .B(_06426_),
    .X(_06445_));
 sky130_fd_sc_hd__o211a_4 _06922_ (.A1(instruction[22]),
    .A2(_06427_),
    .B1(_06445_),
    .C1(net287),
    .X(reg2_idx[4]));
 sky130_fd_sc_hd__nor3_2 _06923_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06422_),
    .Y(_06446_));
 sky130_fd_sc_hd__or3_4 _06924_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06422_),
    .X(_06447_));
 sky130_fd_sc_hd__or2_2 _06925_ (.A(instruction[6]),
    .B(instruction[5]),
    .X(_06448_));
 sky130_fd_sc_hd__nand2_4 _06926_ (.A(_04417_),
    .B(instruction[4]),
    .Y(_06449_));
 sky130_fd_sc_hd__nor2_1 _06927_ (.A(_06448_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__or2_2 _06928_ (.A(_06448_),
    .B(_06449_),
    .X(_06451_));
 sky130_fd_sc_hd__a31o_1 _06929_ (.A1(instruction[17]),
    .A2(_06447_),
    .A3(_06451_),
    .B1(net290),
    .X(_06452_));
 sky130_fd_sc_hd__nor2_1 _06930_ (.A(instruction[6]),
    .B(is_load),
    .Y(_06453_));
 sky130_fd_sc_hd__o211a_1 _06931_ (.A1(instruction[40]),
    .A2(_04589_),
    .B1(_06452_),
    .C1(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__a32o_2 _06932_ (.A1(instruction[24]),
    .A2(net310),
    .A3(is_load),
    .B1(_04633_),
    .B2(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__nand2_8 _06933_ (.A(net266),
    .B(_06455_),
    .Y(dest_mask[0]));
 sky130_fd_sc_hd__a22o_2 _06934_ (.A1(net310),
    .A2(is_load),
    .B1(_04644_),
    .B2(_06454_),
    .X(_06456_));
 sky130_fd_sc_hd__nand2_8 _06935_ (.A(net266),
    .B(_06456_),
    .Y(dest_mask[1]));
 sky130_fd_sc_hd__nand2b_2 _06936_ (.A_N(instruction[6]),
    .B(instruction[5]),
    .Y(_06457_));
 sky130_fd_sc_hd__nor2_2 _06937_ (.A(_06407_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__and2_4 _06938_ (.A(net309),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__nand2_4 _06939_ (.A(net309),
    .B(_06458_),
    .Y(_06460_));
 sky130_fd_sc_hd__and2_1 _06940_ (.A(reg1_val[31]),
    .B(net310),
    .X(_06461_));
 sky130_fd_sc_hd__or4_2 _06941_ (.A(net308),
    .B(net307),
    .C(reg1_val[2]),
    .D(reg1_val[3]),
    .X(_06462_));
 sky130_fd_sc_hd__or4_1 _06942_ (.A(reg1_val[4]),
    .B(reg1_val[5]),
    .C(reg1_val[6]),
    .D(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__or4_2 _06943_ (.A(reg1_val[7]),
    .B(reg1_val[8]),
    .C(reg1_val[9]),
    .D(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__or4_4 _06944_ (.A(reg1_val[10]),
    .B(reg1_val[11]),
    .C(reg1_val[12]),
    .D(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__nand2_1 _06945_ (.A(net282),
    .B(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__xor2_2 _06946_ (.A(reg1_val[13]),
    .B(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__o21a_1 _06947_ (.A1(reg1_val[10]),
    .A2(_06464_),
    .B1(net282),
    .X(_06468_));
 sky130_fd_sc_hd__xnor2_4 _06948_ (.A(reg1_val[11]),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__inv_6 _06949_ (.A(net186),
    .Y(_06470_));
 sky130_fd_sc_hd__o31a_2 _06950_ (.A1(reg1_val[10]),
    .A2(reg1_val[11]),
    .A3(_06464_),
    .B1(net282),
    .X(_06471_));
 sky130_fd_sc_hd__xnor2_4 _06951_ (.A(reg1_val[12]),
    .B(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__nor2_1 _06952_ (.A(net186),
    .B(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__or2_1 _06953_ (.A(net186),
    .B(_06472_),
    .X(_06474_));
 sky130_fd_sc_hd__nand2_1 _06954_ (.A(net186),
    .B(_06472_),
    .Y(_06475_));
 sky130_fd_sc_hd__mux2_1 _06955_ (.A0(_06475_),
    .A1(_06474_),
    .S(net153),
    .X(_06476_));
 sky130_fd_sc_hd__and2_2 _06956_ (.A(net310),
    .B(_04687_),
    .X(_06477_));
 sky130_fd_sc_hd__nand2_8 _06957_ (.A(net310),
    .B(_04687_),
    .Y(_06478_));
 sky130_fd_sc_hd__and4_1 _06958_ (.A(net238),
    .B(net235),
    .C(net232),
    .D(net228),
    .X(_06479_));
 sky130_fd_sc_hd__or4_4 _06959_ (.A(net237),
    .B(net234),
    .C(net230),
    .D(net224),
    .X(_06480_));
 sky130_fd_sc_hd__or4_4 _06960_ (.A(_06256_),
    .B(_06307_),
    .C(_06317_),
    .D(net242),
    .X(_06481_));
 sky130_fd_sc_hd__nor2_1 _06961_ (.A(_06480_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__or2_1 _06962_ (.A(_06480_),
    .B(_06481_),
    .X(_06483_));
 sky130_fd_sc_hd__or4_1 _06963_ (.A(_06065_),
    .B(_06114_),
    .C(_06150_),
    .D(_06202_),
    .X(_06484_));
 sky130_fd_sc_hd__or3_2 _06964_ (.A(_06480_),
    .B(_06481_),
    .C(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__or2_1 _06965_ (.A(_05854_),
    .B(_05907_),
    .X(_06486_));
 sky130_fd_sc_hd__nor4_2 _06966_ (.A(_05955_),
    .B(_05999_),
    .C(_06484_),
    .D(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__or4_2 _06967_ (.A(_05955_),
    .B(_05999_),
    .C(_06484_),
    .D(_06486_),
    .X(_06488_));
 sky130_fd_sc_hd__a21o_1 _06968_ (.A1(_06482_),
    .A2(_06487_),
    .B1(_06478_),
    .X(_06489_));
 sky130_fd_sc_hd__a21oi_1 _06969_ (.A1(_06482_),
    .A2(_06487_),
    .B1(_05799_),
    .Y(_06490_));
 sky130_fd_sc_hd__a22o_4 _06970_ (.A1(_05799_),
    .A2(_06489_),
    .B1(_06490_),
    .B2(net196),
    .X(_06491_));
 sky130_fd_sc_hd__nand2_2 _06971_ (.A(_06474_),
    .B(_06475_),
    .Y(_06492_));
 sky130_fd_sc_hd__a31o_1 _06972_ (.A1(_05799_),
    .A2(_06482_),
    .A3(_06487_),
    .B1(_06478_),
    .X(_06493_));
 sky130_fd_sc_hd__xnor2_4 _06973_ (.A(_05734_),
    .B(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__o22a_1 _06974_ (.A1(net125),
    .A2(_06491_),
    .B1(net121),
    .B2(net119),
    .X(_06495_));
 sky130_fd_sc_hd__xnor2_1 _06975_ (.A(net153),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__o21a_1 _06976_ (.A1(reg1_val[13]),
    .A2(_06465_),
    .B1(net282),
    .X(_06497_));
 sky130_fd_sc_hd__o31a_4 _06977_ (.A1(reg1_val[13]),
    .A2(reg1_val[14]),
    .A3(_06465_),
    .B1(net281),
    .X(_06498_));
 sky130_fd_sc_hd__xor2_4 _06978_ (.A(reg1_val[15]),
    .B(_06498_),
    .X(_06499_));
 sky130_fd_sc_hd__xnor2_4 _06979_ (.A(reg1_val[15]),
    .B(_06498_),
    .Y(_06500_));
 sky130_fd_sc_hd__o31a_2 _06980_ (.A1(_05955_),
    .A2(_05999_),
    .A3(_06485_),
    .B1(net196),
    .X(_06501_));
 sky130_fd_sc_hd__xnor2_4 _06981_ (.A(_05907_),
    .B(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__xnor2_4 _06982_ (.A(reg1_val[14]),
    .B(_06497_),
    .Y(_06503_));
 sky130_fd_sc_hd__or3_1 _06983_ (.A(net152),
    .B(net151),
    .C(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__nand3_1 _06984_ (.A(net152),
    .B(net151),
    .C(_06503_),
    .Y(_06505_));
 sky130_fd_sc_hd__and2_1 _06985_ (.A(_06504_),
    .B(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__xnor2_2 _06986_ (.A(net153),
    .B(_06503_),
    .Y(_06507_));
 sky130_fd_sc_hd__o41a_2 _06987_ (.A1(_05907_),
    .A2(_05955_),
    .A3(_05999_),
    .A4(_06485_),
    .B1(net196),
    .X(_06508_));
 sky130_fd_sc_hd__xnor2_4 _06988_ (.A(_05854_),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__o22a_1 _06989_ (.A1(_06502_),
    .A2(net74),
    .B1(net115),
    .B2(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__xnor2_1 _06990_ (.A(net149),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__or2_1 _06991_ (.A(_06496_),
    .B(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__nand2_1 _06992_ (.A(_06496_),
    .B(_06511_),
    .Y(_06513_));
 sky130_fd_sc_hd__and2_1 _06993_ (.A(_06512_),
    .B(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__or4_4 _06994_ (.A(reg1_val[13]),
    .B(reg1_val[14]),
    .C(reg1_val[15]),
    .D(_06465_),
    .X(_06515_));
 sky130_fd_sc_hd__or3_1 _06995_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .C(reg1_val[22]),
    .X(_06516_));
 sky130_fd_sc_hd__or2_1 _06996_ (.A(reg1_val[16]),
    .B(reg1_val[17]),
    .X(_06517_));
 sky130_fd_sc_hd__or3_4 _06997_ (.A(reg1_val[18]),
    .B(reg1_val[19]),
    .C(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__or3_4 _06998_ (.A(reg1_val[23]),
    .B(_06516_),
    .C(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__or3_1 _06999_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .C(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__o21a_1 _07000_ (.A1(_06515_),
    .A2(_06520_),
    .B1(net281),
    .X(_06521_));
 sky130_fd_sc_hd__o31a_2 _07001_ (.A1(reg1_val[26]),
    .A2(_06515_),
    .A3(_06520_),
    .B1(net281),
    .X(_06522_));
 sky130_fd_sc_hd__xor2_4 _07002_ (.A(reg1_val[27]),
    .B(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__inv_8 _07003_ (.A(net111),
    .Y(_06524_));
 sky130_fd_sc_hd__and3_2 _07004_ (.A(net310),
    .B(_04687_),
    .C(net224),
    .X(_06525_));
 sky130_fd_sc_hd__xnor2_4 _07005_ (.A(net232),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__xnor2_1 _07006_ (.A(net230),
    .B(_06525_),
    .Y(_06527_));
 sky130_fd_sc_hd__o21ai_2 _07007_ (.A1(_06515_),
    .A2(_06519_),
    .B1(net281),
    .Y(_06528_));
 sky130_fd_sc_hd__o31a_1 _07008_ (.A1(reg1_val[24]),
    .A2(_06515_),
    .A3(_06519_),
    .B1(net281),
    .X(_06529_));
 sky130_fd_sc_hd__xor2_1 _07009_ (.A(reg1_val[25]),
    .B(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__xor2_4 _07010_ (.A(reg1_val[26]),
    .B(_06521_),
    .X(_06531_));
 sky130_fd_sc_hd__and2_1 _07011_ (.A(net110),
    .B(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__and3b_1 _07012_ (.A_N(net112),
    .B(net108),
    .C(_06531_),
    .X(_06533_));
 sky130_fd_sc_hd__nor2_1 _07013_ (.A(net108),
    .B(_06531_),
    .Y(_06534_));
 sky130_fd_sc_hd__a21oi_1 _07014_ (.A1(net112),
    .A2(_06534_),
    .B1(_06533_),
    .Y(_06535_));
 sky130_fd_sc_hd__o211a_1 _07015_ (.A1(net230),
    .A2(net224),
    .B1(net310),
    .C1(_04687_),
    .X(_06536_));
 sky130_fd_sc_hd__xnor2_1 _07016_ (.A(net234),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__or2_2 _07017_ (.A(_06532_),
    .B(_06534_),
    .X(_06538_));
 sky130_fd_sc_hd__o22a_1 _07018_ (.A1(net185),
    .A2(net30),
    .B1(net183),
    .B2(net28),
    .X(_06539_));
 sky130_fd_sc_hd__xnor2_2 _07019_ (.A(_06524_),
    .B(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__o21ai_2 _07020_ (.A1(_06515_),
    .A2(_06518_),
    .B1(net281),
    .Y(_06541_));
 sky130_fd_sc_hd__o31a_2 _07021_ (.A1(_06515_),
    .A2(_06516_),
    .A3(_06518_),
    .B1(net281),
    .X(_06542_));
 sky130_fd_sc_hd__xor2_4 _07022_ (.A(reg1_val[23]),
    .B(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__and3_1 _07023_ (.A(net310),
    .B(_04687_),
    .C(net242),
    .X(_06544_));
 sky130_fd_sc_hd__a211o_1 _07024_ (.A1(_06324_),
    .A2(_06479_),
    .B1(_06478_),
    .C1(_06317_),
    .X(_06545_));
 sky130_fd_sc_hd__a211o_1 _07025_ (.A1(net196),
    .A2(_06480_),
    .B1(_06544_),
    .C1(_06316_),
    .X(_06546_));
 sky130_fd_sc_hd__and2_2 _07026_ (.A(_06545_),
    .B(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__o31a_1 _07027_ (.A1(reg1_val[20]),
    .A2(_06515_),
    .A3(_06518_),
    .B1(net281),
    .X(_06548_));
 sky130_fd_sc_hd__xor2_1 _07028_ (.A(reg1_val[21]),
    .B(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__o41a_2 _07029_ (.A1(reg1_val[20]),
    .A2(reg1_val[21]),
    .A3(_06515_),
    .A4(_06518_),
    .B1(net281),
    .X(_06550_));
 sky130_fd_sc_hd__xor2_4 _07030_ (.A(reg1_val[22]),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__nand3b_4 _07031_ (.A_N(_06543_),
    .B(net103),
    .C(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__or3b_4 _07032_ (.A(net103),
    .B(_06551_),
    .C_N(_06543_),
    .X(_06553_));
 sky130_fd_sc_hd__and2_1 _07033_ (.A(_06552_),
    .B(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__a31o_4 _07034_ (.A1(_06316_),
    .A2(_06324_),
    .A3(_06479_),
    .B1(_06478_),
    .X(_06555_));
 sky130_fd_sc_hd__xnor2_4 _07035_ (.A(_06307_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__xor2_4 _07036_ (.A(_06307_),
    .B(_06555_),
    .X(_06557_));
 sky130_fd_sc_hd__xnor2_2 _07037_ (.A(net103),
    .B(_06551_),
    .Y(_06558_));
 sky130_fd_sc_hd__o22a_1 _07038_ (.A1(net148),
    .A2(net25),
    .B1(net146),
    .B2(net72),
    .X(_06559_));
 sky130_fd_sc_hd__xor2_2 _07039_ (.A(net107),
    .B(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__nor2_1 _07040_ (.A(_06540_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__xor2_2 _07041_ (.A(_06540_),
    .B(_06560_),
    .X(_06562_));
 sky130_fd_sc_hd__o311a_2 _07042_ (.A1(net234),
    .A2(net230),
    .A3(net224),
    .B1(_04687_),
    .C1(net310),
    .X(_06563_));
 sky130_fd_sc_hd__xnor2_2 _07043_ (.A(net237),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_4 _07044_ (.A(_06330_),
    .B(_06563_),
    .Y(_06565_));
 sky130_fd_sc_hd__xnor2_4 _07045_ (.A(reg1_val[24]),
    .B(_06528_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand3b_2 _07046_ (.A_N(net108),
    .B(net105),
    .C(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__or3b_2 _07047_ (.A(net105),
    .B(_00136_),
    .C_N(net108),
    .X(_00138_));
 sky130_fd_sc_hd__and2_1 _07048_ (.A(_00137_),
    .B(_00138_),
    .X(_00139_));
 sky130_fd_sc_hd__a21o_2 _07049_ (.A1(net196),
    .A2(_06480_),
    .B1(net242),
    .X(_00140_));
 sky130_fd_sc_hd__or3_2 _07050_ (.A(_06324_),
    .B(_06478_),
    .C(_06479_),
    .X(_00141_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(_00140_),
    .B(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__xnor2_4 _07052_ (.A(net107),
    .B(_00136_),
    .Y(_00143_));
 sky130_fd_sc_hd__o22a_1 _07053_ (.A1(net180),
    .A2(net23),
    .B1(net144),
    .B2(net70),
    .X(_00144_));
 sky130_fd_sc_hd__xnor2_2 _07054_ (.A(net110),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__a21o_1 _07055_ (.A1(_06562_),
    .A2(_00145_),
    .B1(_06561_),
    .X(_00146_));
 sky130_fd_sc_hd__and2_1 _07056_ (.A(_06514_),
    .B(_00146_),
    .X(_00147_));
 sky130_fd_sc_hd__xnor2_1 _07057_ (.A(_06514_),
    .B(_00146_),
    .Y(_00148_));
 sky130_fd_sc_hd__o41a_4 _07058_ (.A1(reg1_val[13]),
    .A2(reg1_val[14]),
    .A3(reg1_val[15]),
    .A4(_06465_),
    .B1(net282),
    .X(_00149_));
 sky130_fd_sc_hd__o211ai_4 _07059_ (.A1(reg1_val[16]),
    .A2(_06515_),
    .B1(net281),
    .C1(reg1_val[17]),
    .Y(_00150_));
 sky130_fd_sc_hd__a211o_2 _07060_ (.A1(reg1_val[16]),
    .A2(net281),
    .B1(_00149_),
    .C1(reg1_val[17]),
    .X(_00151_));
 sky130_fd_sc_hd__and2_4 _07061_ (.A(_00150_),
    .B(_00151_),
    .X(_00152_));
 sky130_fd_sc_hd__nand2_8 _07062_ (.A(_00150_),
    .B(_00151_),
    .Y(_00153_));
 sky130_fd_sc_hd__o41a_4 _07063_ (.A1(_06150_),
    .A2(_06202_),
    .A3(_06480_),
    .A4(_06481_),
    .B1(net196),
    .X(_00154_));
 sky130_fd_sc_hd__and3_1 _07064_ (.A(net309),
    .B(_04687_),
    .C(_06114_),
    .X(_00155_));
 sky130_fd_sc_hd__o21bai_2 _07065_ (.A1(_00154_),
    .A2(_00155_),
    .B1_N(_06065_),
    .Y(_00156_));
 sky130_fd_sc_hd__or3b_2 _07066_ (.A(_00154_),
    .B(_00155_),
    .C_N(_06065_),
    .X(_00157_));
 sky130_fd_sc_hd__and2_4 _07067_ (.A(_00156_),
    .B(_00157_),
    .X(_00158_));
 sky130_fd_sc_hd__xor2_4 _07068_ (.A(reg1_val[16]),
    .B(_00149_),
    .X(_00159_));
 sky130_fd_sc_hd__xnor2_1 _07069_ (.A(reg1_val[16]),
    .B(_00149_),
    .Y(_00160_));
 sky130_fd_sc_hd__a211o_1 _07070_ (.A1(_00150_),
    .A2(_00151_),
    .B1(_00160_),
    .C1(net149),
    .X(_00161_));
 sky130_fd_sc_hd__nand4_1 _07071_ (.A(net149),
    .B(_00150_),
    .C(_00151_),
    .D(_00160_),
    .Y(_00162_));
 sky130_fd_sc_hd__and2_1 _07072_ (.A(_00161_),
    .B(_00162_),
    .X(_00163_));
 sky130_fd_sc_hd__a21o_1 _07073_ (.A1(net196),
    .A2(_06485_),
    .B1(_05999_),
    .X(_00164_));
 sky130_fd_sc_hd__nand3_2 _07074_ (.A(_05999_),
    .B(net196),
    .C(_06485_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_4 _07075_ (.A(_00164_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__xnor2_4 _07076_ (.A(_06499_),
    .B(_00159_),
    .Y(_00167_));
 sky130_fd_sc_hd__o22a_1 _07077_ (.A1(net98),
    .A2(net68),
    .B1(net96),
    .B2(net94),
    .X(_00168_));
 sky130_fd_sc_hd__xnor2_1 _07078_ (.A(net100),
    .B(_00168_),
    .Y(_00169_));
 sky130_fd_sc_hd__o41a_2 _07079_ (.A1(_06307_),
    .A2(_06317_),
    .A3(net242),
    .A4(_06480_),
    .B1(net196),
    .X(_00170_));
 sky130_fd_sc_hd__xnor2_4 _07080_ (.A(_06256_),
    .B(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__o21ai_2 _07081_ (.A1(_06515_),
    .A2(_06517_),
    .B1(net281),
    .Y(_00172_));
 sky130_fd_sc_hd__o31a_1 _07082_ (.A1(reg1_val[18]),
    .A2(_06515_),
    .A3(_06517_),
    .B1(net281),
    .X(_00173_));
 sky130_fd_sc_hd__xor2_4 _07083_ (.A(reg1_val[19]),
    .B(_00173_),
    .X(_00174_));
 sky130_fd_sc_hd__xnor2_4 _07084_ (.A(reg1_val[20]),
    .B(_06541_),
    .Y(_00175_));
 sky130_fd_sc_hd__o21a_4 _07085_ (.A1(net91),
    .A2(_00175_),
    .B1(net102),
    .X(_00176_));
 sky130_fd_sc_hd__a21oi_4 _07086_ (.A1(net91),
    .A2(_00175_),
    .B1(net102),
    .Y(_00177_));
 sky130_fd_sc_hd__or2_4 _07087_ (.A(_00176_),
    .B(_00177_),
    .X(_00178_));
 sky130_fd_sc_hd__o21a_1 _07088_ (.A1(_06480_),
    .A2(_06481_),
    .B1(net196),
    .X(_00179_));
 sky130_fd_sc_hd__xnor2_4 _07089_ (.A(_06202_),
    .B(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__xnor2_1 _07090_ (.A(net93),
    .B(_00175_),
    .Y(_00181_));
 sky130_fd_sc_hd__o22a_1 _07091_ (.A1(net142),
    .A2(net22),
    .B1(net140),
    .B2(net67),
    .X(_00182_));
 sky130_fd_sc_hd__xnor2_1 _07092_ (.A(net102),
    .B(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__xor2_1 _07093_ (.A(_00169_),
    .B(_00183_),
    .X(_00184_));
 sky130_fd_sc_hd__o31a_2 _07094_ (.A1(_06202_),
    .A2(_06480_),
    .A3(_06481_),
    .B1(net196),
    .X(_00185_));
 sky130_fd_sc_hd__xnor2_4 _07095_ (.A(_06150_),
    .B(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__xnor2_4 _07096_ (.A(reg1_val[18]),
    .B(_00172_),
    .Y(_00187_));
 sky130_fd_sc_hd__or3b_4 _07097_ (.A(_00153_),
    .B(net93),
    .C_N(_00187_),
    .X(_00188_));
 sky130_fd_sc_hd__or3b_4 _07098_ (.A(net100),
    .B(_00187_),
    .C_N(net93),
    .X(_00189_));
 sky130_fd_sc_hd__and2_1 _07099_ (.A(_00188_),
    .B(_00189_),
    .X(_00190_));
 sky130_fd_sc_hd__xnor2_4 _07100_ (.A(_06114_),
    .B(_00154_),
    .Y(_00191_));
 sky130_fd_sc_hd__xnor2_2 _07101_ (.A(net101),
    .B(_00187_),
    .Y(_00192_));
 sky130_fd_sc_hd__o22a_1 _07102_ (.A1(net137),
    .A2(net20),
    .B1(net135),
    .B2(net64),
    .X(_00193_));
 sky130_fd_sc_hd__xnor2_1 _07103_ (.A(net91),
    .B(_00193_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _07104_ (.A(_00184_),
    .B(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__a21bo_1 _07105_ (.A1(_00169_),
    .A2(_00183_),
    .B1_N(_00195_),
    .X(_00196_));
 sky130_fd_sc_hd__and2b_1 _07106_ (.A_N(_00148_),
    .B(_00196_),
    .X(_00197_));
 sky130_fd_sc_hd__or2_2 _07107_ (.A(_00147_),
    .B(_00197_),
    .X(_00198_));
 sky130_fd_sc_hd__o22a_1 _07108_ (.A1(net30),
    .A2(net183),
    .B1(net28),
    .B2(net180),
    .X(_00199_));
 sky130_fd_sc_hd__xnor2_1 _07109_ (.A(_06523_),
    .B(_00199_),
    .Y(_00200_));
 sky130_fd_sc_hd__o22a_1 _07110_ (.A1(net25),
    .A2(net146),
    .B1(net72),
    .B2(net142),
    .X(_00201_));
 sky130_fd_sc_hd__xnor2_1 _07111_ (.A(net107),
    .B(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__and2_1 _07112_ (.A(_00200_),
    .B(_00202_),
    .X(_00203_));
 sky130_fd_sc_hd__xor2_1 _07113_ (.A(_00200_),
    .B(_00202_),
    .X(_00204_));
 sky130_fd_sc_hd__o22a_1 _07114_ (.A1(net23),
    .A2(net144),
    .B1(net70),
    .B2(net148),
    .X(_00205_));
 sky130_fd_sc_hd__xnor2_1 _07115_ (.A(net110),
    .B(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__xor2_1 _07116_ (.A(_00204_),
    .B(_00206_),
    .X(_00207_));
 sky130_fd_sc_hd__inv_2 _07117_ (.A(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__o31a_2 _07118_ (.A1(net308),
    .A2(net307),
    .A3(reg1_val[2]),
    .B1(net282),
    .X(_00209_));
 sky130_fd_sc_hd__xor2_4 _07119_ (.A(reg1_val[3]),
    .B(_00209_),
    .X(_00210_));
 sky130_fd_sc_hd__xnor2_1 _07120_ (.A(reg1_val[3]),
    .B(_00209_),
    .Y(_00211_));
 sky130_fd_sc_hd__and3_2 _07121_ (.A(net308),
    .B(reg1_val[31]),
    .C(instruction[7]),
    .X(_00212_));
 sky130_fd_sc_hd__xor2_4 _07122_ (.A(net307),
    .B(_00212_),
    .X(_00213_));
 sky130_fd_sc_hd__xnor2_1 _07123_ (.A(net307),
    .B(_00212_),
    .Y(_00214_));
 sky130_fd_sc_hd__o21a_1 _07124_ (.A1(net308),
    .A2(net307),
    .B1(net282),
    .X(_00215_));
 sky130_fd_sc_hd__xnor2_2 _07125_ (.A(reg1_val[2]),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__or2_1 _07126_ (.A(net260),
    .B(_00216_),
    .X(_00217_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(net260),
    .B(_00216_),
    .Y(_00218_));
 sky130_fd_sc_hd__mux2_1 _07128_ (.A0(_00217_),
    .A1(_00218_),
    .S(_00210_),
    .X(_00219_));
 sky130_fd_sc_hd__and2_1 _07129_ (.A(_05734_),
    .B(_05799_),
    .X(_00220_));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(_05734_),
    .B(_05799_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _07131_ (.A(_05567_),
    .B(_05649_),
    .Y(_00222_));
 sky130_fd_sc_hd__nor4_2 _07132_ (.A(_06483_),
    .B(_06488_),
    .C(_00221_),
    .D(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__or4_4 _07133_ (.A(_06483_),
    .B(_06488_),
    .C(_00221_),
    .D(_00222_),
    .X(_00224_));
 sky130_fd_sc_hd__nand2_1 _07134_ (.A(_05416_),
    .B(_05491_),
    .Y(_00225_));
 sky130_fd_sc_hd__and4_2 _07135_ (.A(_05275_),
    .B(_05340_),
    .C(_05416_),
    .D(_05491_),
    .X(_00226_));
 sky130_fd_sc_hd__a21oi_1 _07136_ (.A1(_00223_),
    .A2(_00226_),
    .B1(_06478_),
    .Y(_00227_));
 sky130_fd_sc_hd__a41o_1 _07137_ (.A1(_05035_),
    .A2(_05166_),
    .A3(_00223_),
    .A4(_00226_),
    .B1(_06478_),
    .X(_00228_));
 sky130_fd_sc_hd__xnor2_1 _07138_ (.A(_05101_),
    .B(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(_00217_),
    .B(_00218_),
    .Y(_00230_));
 sky130_fd_sc_hd__and3_1 _07140_ (.A(_05035_),
    .B(_05101_),
    .C(_05166_),
    .X(_00231_));
 sky130_fd_sc_hd__and3_1 _07141_ (.A(_00223_),
    .B(_00226_),
    .C(_00231_),
    .X(_00232_));
 sky130_fd_sc_hd__nand4_2 _07142_ (.A(_04731_),
    .B(_00223_),
    .C(_00226_),
    .D(_00231_),
    .Y(_00233_));
 sky130_fd_sc_hd__a41o_2 _07143_ (.A1(_04731_),
    .A2(_00223_),
    .A3(_00226_),
    .A4(_00231_),
    .B1(_06478_),
    .X(_00234_));
 sky130_fd_sc_hd__or2_1 _07144_ (.A(_04731_),
    .B(_06478_),
    .X(_00235_));
 sky130_fd_sc_hd__a2bb2o_1 _07145_ (.A1_N(_00232_),
    .A2_N(_00235_),
    .B1(_00234_),
    .B2(_04731_),
    .X(_00236_));
 sky130_fd_sc_hd__o22a_1 _07146_ (.A1(net178),
    .A2(net63),
    .B1(net175),
    .B2(net60),
    .X(_00237_));
 sky130_fd_sc_hd__xnor2_1 _07147_ (.A(_00210_),
    .B(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__and2_1 _07148_ (.A(net306),
    .B(net307),
    .X(_00239_));
 sky130_fd_sc_hd__nand2_1 _07149_ (.A(net306),
    .B(net307),
    .Y(_00240_));
 sky130_fd_sc_hd__xnor2_1 _07150_ (.A(_04970_),
    .B(_00234_),
    .Y(_00241_));
 sky130_fd_sc_hd__xor2_2 _07151_ (.A(_04970_),
    .B(_00234_),
    .X(_00242_));
 sky130_fd_sc_hd__a311o_4 _07152_ (.A1(_04731_),
    .A2(_04970_),
    .A3(_00232_),
    .B1(_06478_),
    .C1(_04883_),
    .X(_00243_));
 sky130_fd_sc_hd__o211ai_4 _07153_ (.A1(_04970_),
    .A2(_06478_),
    .B1(_00234_),
    .C1(_04883_),
    .Y(_00244_));
 sky130_fd_sc_hd__and2_1 _07154_ (.A(_00243_),
    .B(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__a2bb2o_1 _07155_ (.A1_N(net306),
    .A2_N(net19),
    .B1(_00239_),
    .B2(_00242_),
    .X(_00246_));
 sky130_fd_sc_hd__xnor2_1 _07156_ (.A(net261),
    .B(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__o21a_2 _07157_ (.A1(reg1_val[4]),
    .A2(_06462_),
    .B1(net282),
    .X(_00248_));
 sky130_fd_sc_hd__xor2_4 _07158_ (.A(reg1_val[5]),
    .B(_00248_),
    .X(_00249_));
 sky130_fd_sc_hd__xnor2_4 _07159_ (.A(reg1_val[5]),
    .B(_00248_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _07160_ (.A(net282),
    .B(_06462_),
    .Y(_00251_));
 sky130_fd_sc_hd__xor2_1 _07161_ (.A(reg1_val[4]),
    .B(_00251_),
    .X(_00252_));
 sky130_fd_sc_hd__or2_1 _07162_ (.A(net213),
    .B(_00252_),
    .X(_00253_));
 sky130_fd_sc_hd__or2_1 _07163_ (.A(_00249_),
    .B(_00253_),
    .X(_00254_));
 sky130_fd_sc_hd__nand2_1 _07164_ (.A(net213),
    .B(_00252_),
    .Y(_00255_));
 sky130_fd_sc_hd__o21a_1 _07165_ (.A1(net211),
    .A2(_00255_),
    .B1(_00254_),
    .X(_00256_));
 sky130_fd_sc_hd__xnor2_1 _07166_ (.A(_05177_),
    .B(_00227_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _07167_ (.A(_00253_),
    .B(_00255_),
    .Y(_00258_));
 sky130_fd_sc_hd__a31o_1 _07168_ (.A1(_05166_),
    .A2(_00223_),
    .A3(_00226_),
    .B1(_06478_),
    .X(_00259_));
 sky130_fd_sc_hd__xnor2_1 _07169_ (.A(_05035_),
    .B(_00259_),
    .Y(_00260_));
 sky130_fd_sc_hd__o22a_1 _07170_ (.A1(net134),
    .A2(net55),
    .B1(net172),
    .B2(net52),
    .X(_00261_));
 sky130_fd_sc_hd__xnor2_1 _07171_ (.A(net211),
    .B(_00261_),
    .Y(_00262_));
 sky130_fd_sc_hd__nor2_1 _07172_ (.A(_00247_),
    .B(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__xor2_1 _07173_ (.A(_00247_),
    .B(_00262_),
    .X(_00264_));
 sky130_fd_sc_hd__xor2_1 _07174_ (.A(_00238_),
    .B(_00264_),
    .X(_00265_));
 sky130_fd_sc_hd__o22a_1 _07175_ (.A1(net123),
    .A2(net121),
    .B1(net114),
    .B2(net125),
    .X(_00266_));
 sky130_fd_sc_hd__xnor2_1 _07176_ (.A(net152),
    .B(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__o21a_1 _07177_ (.A1(_05999_),
    .A2(_06485_),
    .B1(net196),
    .X(_00268_));
 sky130_fd_sc_hd__xnor2_4 _07178_ (.A(_05955_),
    .B(_00268_),
    .Y(_00269_));
 sky130_fd_sc_hd__o22a_1 _07179_ (.A1(net118),
    .A2(net115),
    .B1(net89),
    .B2(net74),
    .X(_00270_));
 sky130_fd_sc_hd__xnor2_1 _07180_ (.A(net149),
    .B(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__or2_1 _07181_ (.A(_00267_),
    .B(_00271_),
    .X(_00272_));
 sky130_fd_sc_hd__nand2_1 _07182_ (.A(net282),
    .B(_06463_),
    .Y(_00273_));
 sky130_fd_sc_hd__xor2_1 _07183_ (.A(reg1_val[7]),
    .B(_00273_),
    .X(_00274_));
 sky130_fd_sc_hd__o31a_1 _07184_ (.A1(reg1_val[4]),
    .A2(reg1_val[5]),
    .A3(_06462_),
    .B1(net282),
    .X(_00275_));
 sky130_fd_sc_hd__xnor2_1 _07185_ (.A(reg1_val[6]),
    .B(_00275_),
    .Y(_00276_));
 sky130_fd_sc_hd__nor2_1 _07186_ (.A(net211),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _07187_ (.A(net195),
    .B(_00277_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _07188_ (.A(net211),
    .B(_00276_),
    .Y(_00279_));
 sky130_fd_sc_hd__o21a_1 _07189_ (.A1(net195),
    .A2(_00279_),
    .B1(_00278_),
    .X(_00280_));
 sky130_fd_sc_hd__o21a_1 _07190_ (.A1(_00224_),
    .A2(_00225_),
    .B1(net196),
    .X(_00281_));
 sky130_fd_sc_hd__xnor2_1 _07191_ (.A(_05351_),
    .B(_00281_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2b_2 _07192_ (.A_N(_00277_),
    .B(_00279_),
    .Y(_00283_));
 sky130_fd_sc_hd__o31a_1 _07193_ (.A1(_05351_),
    .A2(_00224_),
    .A3(_00225_),
    .B1(net196),
    .X(_00284_));
 sky130_fd_sc_hd__xor2_1 _07194_ (.A(_05275_),
    .B(_00284_),
    .X(_00285_));
 sky130_fd_sc_hd__o22a_1 _07195_ (.A1(net132),
    .A2(net49),
    .B1(net170),
    .B2(net46),
    .X(_00286_));
 sky130_fd_sc_hd__xnor2_1 _07196_ (.A(net194),
    .B(_00286_),
    .Y(_00287_));
 sky130_fd_sc_hd__o21a_1 _07197_ (.A1(reg1_val[7]),
    .A2(_06463_),
    .B1(net282),
    .X(_00288_));
 sky130_fd_sc_hd__a21o_1 _07198_ (.A1(reg1_val[8]),
    .A2(net282),
    .B1(_00288_),
    .X(_00289_));
 sky130_fd_sc_hd__xnor2_1 _07199_ (.A(reg1_val[9]),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _07200_ (.A(net282),
    .B(_06464_),
    .Y(_00291_));
 sky130_fd_sc_hd__xor2_1 _07201_ (.A(reg1_val[10]),
    .B(_00291_),
    .X(_00292_));
 sky130_fd_sc_hd__or2_1 _07202_ (.A(net167),
    .B(_00292_),
    .X(_00293_));
 sky130_fd_sc_hd__nand2_1 _07203_ (.A(net167),
    .B(_00292_),
    .Y(_00294_));
 sky130_fd_sc_hd__mux2_4 _07204_ (.A0(_00293_),
    .A1(_00294_),
    .S(_06470_),
    .X(_00295_));
 sky130_fd_sc_hd__a31o_1 _07205_ (.A1(_06482_),
    .A2(_06487_),
    .A3(_00220_),
    .B1(_06478_),
    .X(_00296_));
 sky130_fd_sc_hd__o31a_1 _07206_ (.A1(_06483_),
    .A2(_06488_),
    .A3(_00221_),
    .B1(_05658_),
    .X(_00297_));
 sky130_fd_sc_hd__a22o_1 _07207_ (.A1(_05649_),
    .A2(_00296_),
    .B1(_00297_),
    .B2(_06477_),
    .X(_00298_));
 sky130_fd_sc_hd__nand2_4 _07208_ (.A(_00293_),
    .B(_00294_),
    .Y(_00299_));
 sky130_fd_sc_hd__a41o_1 _07209_ (.A1(_05649_),
    .A2(_06482_),
    .A3(_06487_),
    .A4(_00220_),
    .B1(_06478_),
    .X(_00300_));
 sky130_fd_sc_hd__xnor2_1 _07210_ (.A(_05567_),
    .B(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__o22a_1 _07211_ (.A1(net88),
    .A2(net86),
    .B1(net83),
    .B2(net81),
    .X(_00302_));
 sky130_fd_sc_hd__xnor2_1 _07212_ (.A(net186),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__nor2_1 _07213_ (.A(_00287_),
    .B(_00303_),
    .Y(_00304_));
 sky130_fd_sc_hd__xor2_1 _07214_ (.A(_00287_),
    .B(_00303_),
    .X(_00305_));
 sky130_fd_sc_hd__xnor2_1 _07215_ (.A(reg1_val[8]),
    .B(_00288_),
    .Y(_00306_));
 sky130_fd_sc_hd__or2_1 _07216_ (.A(net194),
    .B(_00306_),
    .X(_00307_));
 sky130_fd_sc_hd__nand2_1 _07217_ (.A(net194),
    .B(_00306_),
    .Y(_00308_));
 sky130_fd_sc_hd__mux2_1 _07218_ (.A0(_00308_),
    .A1(_00307_),
    .S(net168),
    .X(_00309_));
 sky130_fd_sc_hd__a21oi_4 _07219_ (.A1(_06477_),
    .A2(_00224_),
    .B1(_05426_),
    .Y(_00310_));
 sky130_fd_sc_hd__and3_2 _07220_ (.A(_05426_),
    .B(_06477_),
    .C(_00224_),
    .X(_00311_));
 sky130_fd_sc_hd__or2_1 _07221_ (.A(_00310_),
    .B(_00311_),
    .X(_00312_));
 sky130_fd_sc_hd__nand2_2 _07222_ (.A(_00307_),
    .B(_00308_),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2_1 _07223_ (.A(_05416_),
    .B(_06478_),
    .Y(_00314_));
 sky130_fd_sc_hd__o211ai_1 _07224_ (.A1(_05426_),
    .A2(_00224_),
    .B1(net196),
    .C1(_05491_),
    .Y(_00315_));
 sky130_fd_sc_hd__a211o_1 _07225_ (.A1(net196),
    .A2(_00224_),
    .B1(_00314_),
    .C1(_05491_),
    .X(_00316_));
 sky130_fd_sc_hd__and2_1 _07226_ (.A(_00315_),
    .B(_00316_),
    .X(_00317_));
 sky130_fd_sc_hd__o22a_1 _07227_ (.A1(net130),
    .A2(net43),
    .B1(net128),
    .B2(net40),
    .X(_00318_));
 sky130_fd_sc_hd__xnor2_1 _07228_ (.A(net168),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__and2b_1 _07229_ (.A_N(_00319_),
    .B(_00305_),
    .X(_00320_));
 sky130_fd_sc_hd__xnor2_1 _07230_ (.A(_00305_),
    .B(_00319_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2b_1 _07231_ (.A_N(_00272_),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__xnor2_1 _07232_ (.A(_00272_),
    .B(_00321_),
    .Y(_00323_));
 sky130_fd_sc_hd__xnor2_1 _07233_ (.A(_00265_),
    .B(_00323_),
    .Y(_00324_));
 sky130_fd_sc_hd__or2_1 _07234_ (.A(_00208_),
    .B(_00324_),
    .X(_00325_));
 sky130_fd_sc_hd__o22a_2 _07235_ (.A1(net55),
    .A2(net172),
    .B1(net46),
    .B2(net134),
    .X(_00326_));
 sky130_fd_sc_hd__xnor2_4 _07236_ (.A(net211),
    .B(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__o22a_2 _07237_ (.A1(net60),
    .A2(net257),
    .B1(net57),
    .B2(net306),
    .X(_00328_));
 sky130_fd_sc_hd__xnor2_4 _07238_ (.A(net260),
    .B(_00328_),
    .Y(_00329_));
 sky130_fd_sc_hd__o22a_2 _07239_ (.A1(net63),
    .A2(net175),
    .B1(net52),
    .B2(net178),
    .X(_00330_));
 sky130_fd_sc_hd__xnor2_4 _07240_ (.A(net213),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__xor2_4 _07241_ (.A(_00327_),
    .B(_00329_),
    .X(_00332_));
 sky130_fd_sc_hd__and2b_1 _07242_ (.A_N(_00331_),
    .B(_00332_),
    .X(_00333_));
 sky130_fd_sc_hd__o21bai_2 _07243_ (.A1(_00327_),
    .A2(_00329_),
    .B1_N(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__o22a_2 _07244_ (.A1(net49),
    .A2(net170),
    .B1(net40),
    .B2(net132),
    .X(_00335_));
 sky130_fd_sc_hd__xnor2_4 _07245_ (.A(net194),
    .B(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__o22a_2 _07246_ (.A1(_06494_),
    .A2(net88),
    .B1(net86),
    .B2(net83),
    .X(_00337_));
 sky130_fd_sc_hd__xnor2_4 _07247_ (.A(_06469_),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__nor2_1 _07248_ (.A(_00336_),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__xor2_4 _07249_ (.A(_00336_),
    .B(_00338_),
    .X(_00340_));
 sky130_fd_sc_hd__o22a_1 _07250_ (.A1(net81),
    .A2(net130),
    .B1(net43),
    .B2(net128),
    .X(_00341_));
 sky130_fd_sc_hd__xnor2_2 _07251_ (.A(net168),
    .B(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__and2b_1 _07252_ (.A_N(_00342_),
    .B(_00340_),
    .X(_00343_));
 sky130_fd_sc_hd__or4_2 _07253_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .C(reg1_val[26]),
    .D(reg1_val[27]),
    .X(_00344_));
 sky130_fd_sc_hd__or4_1 _07254_ (.A(reg1_val[28]),
    .B(_06515_),
    .C(_06519_),
    .D(_00344_),
    .X(_00345_));
 sky130_fd_sc_hd__o41a_1 _07255_ (.A1(reg1_val[28]),
    .A2(_06515_),
    .A3(_06519_),
    .A4(_00344_),
    .B1(net281),
    .X(_00346_));
 sky130_fd_sc_hd__xnor2_1 _07256_ (.A(reg1_val[29]),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_4 _07257_ (.A(net76),
    .Y(_00348_));
 sky130_fd_sc_hd__o31a_2 _07258_ (.A1(_06515_),
    .A2(_06519_),
    .A3(_00344_),
    .B1(net281),
    .X(_00349_));
 sky130_fd_sc_hd__xor2_4 _07259_ (.A(reg1_val[28]),
    .B(_00349_),
    .X(_00350_));
 sky130_fd_sc_hd__o21ba_1 _07260_ (.A1(net112),
    .A2(_00350_),
    .B1_N(net77),
    .X(_00351_));
 sky130_fd_sc_hd__a21boi_1 _07261_ (.A1(net112),
    .A2(_00350_),
    .B1_N(net77),
    .Y(_00352_));
 sky130_fd_sc_hd__or2_1 _07262_ (.A(_00351_),
    .B(_00352_),
    .X(_00353_));
 sky130_fd_sc_hd__xnor2_4 _07263_ (.A(net112),
    .B(_00350_),
    .Y(_00354_));
 sky130_fd_sc_hd__o22a_1 _07264_ (.A1(net229),
    .A2(net16),
    .B1(net37),
    .B2(net185),
    .X(_00355_));
 sky130_fd_sc_hd__xnor2_1 _07265_ (.A(_00348_),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__o21a_1 _07266_ (.A1(_00339_),
    .A2(_00343_),
    .B1(_00356_),
    .X(_00357_));
 sky130_fd_sc_hd__nor3_1 _07267_ (.A(_00339_),
    .B(_00343_),
    .C(_00356_),
    .Y(_00358_));
 sky130_fd_sc_hd__nor2_1 _07268_ (.A(_00357_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__xnor2_2 _07269_ (.A(_00334_),
    .B(_00359_),
    .Y(_00360_));
 sky130_fd_sc_hd__xnor2_1 _07270_ (.A(_00208_),
    .B(_00324_),
    .Y(_00361_));
 sky130_fd_sc_hd__o21a_2 _07271_ (.A1(_00360_),
    .A2(_00361_),
    .B1(_00325_),
    .X(_00362_));
 sky130_fd_sc_hd__o21bai_1 _07272_ (.A1(_00147_),
    .A2(_00197_),
    .B1_N(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__o22a_1 _07273_ (.A1(net69),
    .A2(net96),
    .B1(net95),
    .B2(net89),
    .X(_00364_));
 sky130_fd_sc_hd__xnor2_1 _07274_ (.A(_00152_),
    .B(_00364_),
    .Y(_00365_));
 sky130_fd_sc_hd__o22a_1 _07275_ (.A1(net22),
    .A2(net140),
    .B1(net66),
    .B2(net137),
    .X(_00366_));
 sky130_fd_sc_hd__xnor2_1 _07276_ (.A(net103),
    .B(_00366_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(_00365_),
    .B(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__xor2_1 _07278_ (.A(_00365_),
    .B(_00367_),
    .X(_00369_));
 sky130_fd_sc_hd__o22a_1 _07279_ (.A1(net20),
    .A2(net135),
    .B1(net64),
    .B2(net98),
    .X(_00370_));
 sky130_fd_sc_hd__xnor2_1 _07280_ (.A(net93),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__xor2_1 _07281_ (.A(_00369_),
    .B(_00371_),
    .X(_00372_));
 sky130_fd_sc_hd__nor2_1 _07282_ (.A(net229),
    .B(net37),
    .Y(_00373_));
 sky130_fd_sc_hd__o22a_1 _07283_ (.A1(net134),
    .A2(net48),
    .B1(net45),
    .B2(net172),
    .X(_00374_));
 sky130_fd_sc_hd__xnor2_1 _07284_ (.A(net211),
    .B(_00374_),
    .Y(_00375_));
 sky130_fd_sc_hd__o22a_1 _07285_ (.A1(net306),
    .A2(net59),
    .B1(net257),
    .B2(net62),
    .X(_00376_));
 sky130_fd_sc_hd__xnor2_1 _07286_ (.A(net260),
    .B(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__nor2_1 _07287_ (.A(_00375_),
    .B(_00377_),
    .Y(_00378_));
 sky130_fd_sc_hd__o22a_1 _07288_ (.A1(net178),
    .A2(net53),
    .B1(net50),
    .B2(net175),
    .X(_00379_));
 sky130_fd_sc_hd__xnor2_1 _07289_ (.A(net213),
    .B(_00379_),
    .Y(_00380_));
 sky130_fd_sc_hd__xor2_1 _07290_ (.A(_00375_),
    .B(_00377_),
    .X(_00381_));
 sky130_fd_sc_hd__and2b_1 _07291_ (.A_N(_00380_),
    .B(_00381_),
    .X(_00382_));
 sky130_fd_sc_hd__or3b_1 _07292_ (.A(_00378_),
    .B(_00382_),
    .C_N(_00373_),
    .X(_00383_));
 sky130_fd_sc_hd__or2_1 _07293_ (.A(_00348_),
    .B(_00373_),
    .X(_00384_));
 sky130_fd_sc_hd__and3_1 _07294_ (.A(_00372_),
    .B(_00383_),
    .C(_00384_),
    .X(_00385_));
 sky130_fd_sc_hd__o22a_1 _07295_ (.A1(net132),
    .A2(net41),
    .B1(net38),
    .B2(net170),
    .X(_00386_));
 sky130_fd_sc_hd__xnor2_1 _07296_ (.A(net194),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__o22a_1 _07297_ (.A1(net84),
    .A2(net130),
    .B1(net128),
    .B2(net79),
    .X(_00388_));
 sky130_fd_sc_hd__xnor2_1 _07298_ (.A(net167),
    .B(_00388_),
    .Y(_00389_));
 sky130_fd_sc_hd__or2_4 _07299_ (.A(_00387_),
    .B(_00389_),
    .X(_00390_));
 sky130_fd_sc_hd__xnor2_4 _07300_ (.A(_00340_),
    .B(_00342_),
    .Y(_00391_));
 sky130_fd_sc_hd__and2b_1 _07301_ (.A_N(_00390_),
    .B(_00391_),
    .X(_00392_));
 sky130_fd_sc_hd__xnor2_4 _07302_ (.A(_00331_),
    .B(_00332_),
    .Y(_00393_));
 sky130_fd_sc_hd__xnor2_4 _07303_ (.A(_00390_),
    .B(_00391_),
    .Y(_00394_));
 sky130_fd_sc_hd__a21oi_4 _07304_ (.A1(_00393_),
    .A2(_00394_),
    .B1(_00392_),
    .Y(_00395_));
 sky130_fd_sc_hd__a21oi_1 _07305_ (.A1(_00383_),
    .A2(_00384_),
    .B1(_00372_),
    .Y(_00396_));
 sky130_fd_sc_hd__nor2_2 _07306_ (.A(_00385_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__and2b_1 _07307_ (.A_N(_00395_),
    .B(_00397_),
    .X(_00398_));
 sky130_fd_sc_hd__or2_2 _07308_ (.A(_00385_),
    .B(_00398_),
    .X(_00399_));
 sky130_fd_sc_hd__xnor2_4 _07309_ (.A(_00198_),
    .B(_00362_),
    .Y(_00400_));
 sky130_fd_sc_hd__a21bo_1 _07310_ (.A1(_00399_),
    .A2(_00400_),
    .B1_N(_00363_),
    .X(_00401_));
 sky130_fd_sc_hd__a21o_1 _07311_ (.A1(_00334_),
    .A2(_00359_),
    .B1(_00357_),
    .X(_00402_));
 sky130_fd_sc_hd__o22a_1 _07312_ (.A1(net30),
    .A2(net180),
    .B1(net144),
    .B2(net28),
    .X(_00403_));
 sky130_fd_sc_hd__xnor2_1 _07313_ (.A(_06523_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__o22a_1 _07314_ (.A1(net25),
    .A2(net142),
    .B1(net140),
    .B2(net72),
    .X(_00405_));
 sky130_fd_sc_hd__xnor2_1 _07315_ (.A(net107),
    .B(_00405_),
    .Y(_00406_));
 sky130_fd_sc_hd__and2_1 _07316_ (.A(_00404_),
    .B(_00406_),
    .X(_00407_));
 sky130_fd_sc_hd__nor2_1 _07317_ (.A(_00404_),
    .B(_00406_),
    .Y(_00408_));
 sky130_fd_sc_hd__or2_1 _07318_ (.A(_00407_),
    .B(_00408_),
    .X(_00409_));
 sky130_fd_sc_hd__o22a_1 _07319_ (.A1(net148),
    .A2(net23),
    .B1(net70),
    .B2(net146),
    .X(_00410_));
 sky130_fd_sc_hd__xor2_1 _07320_ (.A(net110),
    .B(_00410_),
    .X(_00411_));
 sky130_fd_sc_hd__nor2_1 _07321_ (.A(_00409_),
    .B(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__and2_1 _07322_ (.A(_00409_),
    .B(_00411_),
    .X(_00413_));
 sky130_fd_sc_hd__nor2_1 _07323_ (.A(_00412_),
    .B(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__a21bo_1 _07324_ (.A1(_00265_),
    .A2(_00323_),
    .B1_N(_00322_),
    .X(_00415_));
 sky130_fd_sc_hd__xnor2_2 _07325_ (.A(_00402_),
    .B(_00414_),
    .Y(_00416_));
 sky130_fd_sc_hd__and2b_1 _07326_ (.A_N(_00416_),
    .B(_00415_),
    .X(_00417_));
 sky130_fd_sc_hd__a21o_1 _07327_ (.A1(_00402_),
    .A2(_00414_),
    .B1(_00417_),
    .X(_00418_));
 sky130_fd_sc_hd__o22a_1 _07328_ (.A1(net88),
    .A2(net81),
    .B1(net43),
    .B2(net83),
    .X(_00419_));
 sky130_fd_sc_hd__xnor2_1 _07329_ (.A(net186),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__o22a_1 _07330_ (.A1(net55),
    .A2(net170),
    .B1(net46),
    .B2(net132),
    .X(_00421_));
 sky130_fd_sc_hd__xnor2_1 _07331_ (.A(net195),
    .B(_00421_),
    .Y(_00422_));
 sky130_fd_sc_hd__nor2_1 _07332_ (.A(_00420_),
    .B(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__and2_1 _07333_ (.A(_00420_),
    .B(_00422_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_1 _07334_ (.A(_00423_),
    .B(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__o22a_1 _07335_ (.A1(net49),
    .A2(net128),
    .B1(net40),
    .B2(net130),
    .X(_00426_));
 sky130_fd_sc_hd__xnor2_1 _07336_ (.A(net168),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__xnor2_1 _07337_ (.A(_00425_),
    .B(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__inv_2 _07338_ (.A(_00428_),
    .Y(_00429_));
 sky130_fd_sc_hd__o22a_1 _07339_ (.A1(net178),
    .A2(net60),
    .B1(net57),
    .B2(net175),
    .X(_00430_));
 sky130_fd_sc_hd__xnor2_2 _07340_ (.A(_00210_),
    .B(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__o22a_1 _07341_ (.A1(net63),
    .A2(net172),
    .B1(net52),
    .B2(net134),
    .X(_00432_));
 sky130_fd_sc_hd__xnor2_2 _07342_ (.A(net211),
    .B(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2b_1 _07343_ (.A_N(_04883_),
    .B(_04970_),
    .Y(_00434_));
 sky130_fd_sc_hd__o21ai_1 _07344_ (.A1(_00233_),
    .A2(_00434_),
    .B1(_06477_),
    .Y(_00435_));
 sky130_fd_sc_hd__xnor2_2 _07345_ (.A(_04818_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__o22a_1 _07346_ (.A1(net257),
    .A2(net19),
    .B1(net14),
    .B2(net306),
    .X(_00437_));
 sky130_fd_sc_hd__xnor2_2 _07347_ (.A(net260),
    .B(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__nor2_1 _07348_ (.A(_00433_),
    .B(_00438_),
    .Y(_00439_));
 sky130_fd_sc_hd__xor2_2 _07349_ (.A(_00433_),
    .B(_00438_),
    .X(_00440_));
 sky130_fd_sc_hd__xnor2_2 _07350_ (.A(_00431_),
    .B(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__o22a_1 _07351_ (.A1(net125),
    .A2(_06494_),
    .B1(net86),
    .B2(net121),
    .X(_00442_));
 sky130_fd_sc_hd__xnor2_1 _07352_ (.A(net153),
    .B(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__o22a_1 _07353_ (.A1(_06502_),
    .A2(net94),
    .B1(_00269_),
    .B2(net69),
    .X(_00444_));
 sky130_fd_sc_hd__xnor2_1 _07354_ (.A(_00152_),
    .B(_00444_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2b_1 _07355_ (.A_N(_00443_),
    .B(_00445_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2b_1 _07356_ (.A_N(_00445_),
    .B(_00443_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_00446_),
    .B(_00447_),
    .Y(_00448_));
 sky130_fd_sc_hd__o22a_1 _07358_ (.A1(_06491_),
    .A2(net115),
    .B1(_06509_),
    .B2(net74),
    .X(_00449_));
 sky130_fd_sc_hd__xnor2_2 _07359_ (.A(net149),
    .B(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__xnor2_2 _07360_ (.A(_00448_),
    .B(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__or2_1 _07361_ (.A(_00441_),
    .B(_00451_),
    .X(_00452_));
 sky130_fd_sc_hd__xnor2_2 _07362_ (.A(_00441_),
    .B(_00451_),
    .Y(_00453_));
 sky130_fd_sc_hd__xnor2_2 _07363_ (.A(_00429_),
    .B(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__o21a_1 _07364_ (.A1(reg1_val[29]),
    .A2(_00345_),
    .B1(net281),
    .X(_00455_));
 sky130_fd_sc_hd__xnor2_4 _07365_ (.A(reg1_val[30]),
    .B(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__xnor2_1 _07366_ (.A(net78),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__nor2_1 _07367_ (.A(net229),
    .B(net11),
    .Y(_00458_));
 sky130_fd_sc_hd__o22a_1 _07368_ (.A1(net185),
    .A2(net16),
    .B1(net37),
    .B2(net183),
    .X(_00459_));
 sky130_fd_sc_hd__xnor2_2 _07369_ (.A(net78),
    .B(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__inv_2 _07370_ (.A(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__xor2_2 _07371_ (.A(_00458_),
    .B(_00460_),
    .X(_00462_));
 sky130_fd_sc_hd__a21o_1 _07372_ (.A1(_00238_),
    .A2(_00264_),
    .B1(_00263_),
    .X(_00463_));
 sky130_fd_sc_hd__and2b_1 _07373_ (.A_N(_06512_),
    .B(_00463_),
    .X(_00464_));
 sky130_fd_sc_hd__xnor2_1 _07374_ (.A(_06512_),
    .B(_00463_),
    .Y(_00465_));
 sky130_fd_sc_hd__o21a_1 _07375_ (.A1(_00304_),
    .A2(_00320_),
    .B1(_00465_),
    .X(_00466_));
 sky130_fd_sc_hd__nor3_1 _07376_ (.A(_00304_),
    .B(_00320_),
    .C(_00465_),
    .Y(_00467_));
 sky130_fd_sc_hd__or2_1 _07377_ (.A(_00466_),
    .B(_00467_),
    .X(_00468_));
 sky130_fd_sc_hd__xnor2_2 _07378_ (.A(_00454_),
    .B(_00462_),
    .Y(_00469_));
 sky130_fd_sc_hd__o32a_1 _07379_ (.A1(_00466_),
    .A2(_00467_),
    .A3(_00469_),
    .B1(_00462_),
    .B2(_00454_),
    .X(_00470_));
 sky130_fd_sc_hd__o22a_1 _07380_ (.A1(net98),
    .A2(net20),
    .B1(net64),
    .B2(net96),
    .X(_00471_));
 sky130_fd_sc_hd__xnor2_1 _07381_ (.A(net93),
    .B(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__o22a_1 _07382_ (.A1(net22),
    .A2(net137),
    .B1(net135),
    .B2(net66),
    .X(_00473_));
 sky130_fd_sc_hd__xnor2_1 _07383_ (.A(net103),
    .B(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__and2_1 _07384_ (.A(_00472_),
    .B(_00474_),
    .X(_00475_));
 sky130_fd_sc_hd__nor2_1 _07385_ (.A(_00472_),
    .B(_00474_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_00475_),
    .B(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__a21o_1 _07387_ (.A1(_00204_),
    .A2(_00206_),
    .B1(_00203_),
    .X(_00478_));
 sky130_fd_sc_hd__a21bo_1 _07388_ (.A1(_00369_),
    .A2(_00371_),
    .B1_N(_00368_),
    .X(_00479_));
 sky130_fd_sc_hd__xnor2_1 _07389_ (.A(_00477_),
    .B(_00478_),
    .Y(_00480_));
 sky130_fd_sc_hd__and2b_1 _07390_ (.A_N(_00480_),
    .B(_00479_),
    .X(_00481_));
 sky130_fd_sc_hd__a21oi_2 _07391_ (.A1(_00477_),
    .A2(_00478_),
    .B1(_00481_),
    .Y(_00482_));
 sky130_fd_sc_hd__or2_1 _07392_ (.A(_00470_),
    .B(_00482_),
    .X(_00483_));
 sky130_fd_sc_hd__xor2_2 _07393_ (.A(_00470_),
    .B(_00482_),
    .X(_00484_));
 sky130_fd_sc_hd__xor2_2 _07394_ (.A(_00418_),
    .B(_00484_),
    .X(_00485_));
 sky130_fd_sc_hd__xor2_2 _07395_ (.A(_00468_),
    .B(_00469_),
    .X(_00486_));
 sky130_fd_sc_hd__xnor2_2 _07396_ (.A(_00479_),
    .B(_00480_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(_00486_),
    .B(_00487_),
    .Y(_00488_));
 sky130_fd_sc_hd__xnor2_2 _07398_ (.A(_00415_),
    .B(_00416_),
    .Y(_00489_));
 sky130_fd_sc_hd__xor2_2 _07399_ (.A(_00486_),
    .B(_00487_),
    .X(_00490_));
 sky130_fd_sc_hd__a21bo_1 _07400_ (.A1(_00489_),
    .A2(_00490_),
    .B1_N(_00488_),
    .X(_00491_));
 sky130_fd_sc_hd__xnor2_2 _07401_ (.A(_00401_),
    .B(_00485_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2b_1 _07402_ (.A_N(_00492_),
    .B(_00491_),
    .Y(_00493_));
 sky130_fd_sc_hd__a21bo_2 _07403_ (.A1(_00401_),
    .A2(_00485_),
    .B1_N(_00493_),
    .X(_00494_));
 sky130_fd_sc_hd__o22a_1 _07404_ (.A1(net125),
    .A2(net86),
    .B1(net81),
    .B2(net121),
    .X(_00495_));
 sky130_fd_sc_hd__xnor2_1 _07405_ (.A(net153),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__o22a_1 _07406_ (.A1(_06502_),
    .A2(net68),
    .B1(net95),
    .B2(_06509_),
    .X(_00497_));
 sky130_fd_sc_hd__xnor2_1 _07407_ (.A(_00152_),
    .B(_00497_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2b_1 _07408_ (.A_N(_00496_),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__xor2_1 _07409_ (.A(_00496_),
    .B(_00498_),
    .X(_00500_));
 sky130_fd_sc_hd__o22a_1 _07410_ (.A1(_06491_),
    .A2(net74),
    .B1(net115),
    .B2(_06494_),
    .X(_00501_));
 sky130_fd_sc_hd__xnor2_1 _07411_ (.A(net149),
    .B(_00501_),
    .Y(_00502_));
 sky130_fd_sc_hd__or2_1 _07412_ (.A(_00500_),
    .B(_00502_),
    .X(_00503_));
 sky130_fd_sc_hd__nand2_1 _07413_ (.A(_00500_),
    .B(_00502_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_2 _07414_ (.A(_00503_),
    .B(_00504_),
    .Y(_00505_));
 sky130_fd_sc_hd__o22a_2 _07415_ (.A1(net178),
    .A2(net57),
    .B1(net19),
    .B2(net175),
    .X(_00506_));
 sky130_fd_sc_hd__xnor2_4 _07416_ (.A(net213),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__inv_2 _07417_ (.A(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__o31a_1 _07418_ (.A1(_04807_),
    .A2(_00233_),
    .A3(_00434_),
    .B1(instruction[7]),
    .X(_00509_));
 sky130_fd_sc_hd__nor2_4 _07419_ (.A(_04676_),
    .B(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__or2_1 _07420_ (.A(_04676_),
    .B(_00509_),
    .X(_00511_));
 sky130_fd_sc_hd__o22a_2 _07421_ (.A1(net257),
    .A2(net14),
    .B1(net7),
    .B2(net306),
    .X(_00512_));
 sky130_fd_sc_hd__xnor2_4 _07422_ (.A(net260),
    .B(_00512_),
    .Y(_00513_));
 sky130_fd_sc_hd__o22a_2 _07423_ (.A1(net63),
    .A2(net134),
    .B1(net172),
    .B2(net60),
    .X(_00514_));
 sky130_fd_sc_hd__xnor2_4 _07424_ (.A(net211),
    .B(_00514_),
    .Y(_00515_));
 sky130_fd_sc_hd__nor2_1 _07425_ (.A(_00513_),
    .B(_00515_),
    .Y(_00516_));
 sky130_fd_sc_hd__xor2_4 _07426_ (.A(_00513_),
    .B(_00515_),
    .X(_00517_));
 sky130_fd_sc_hd__xnor2_4 _07427_ (.A(_00507_),
    .B(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__o22a_1 _07428_ (.A1(net88),
    .A2(net43),
    .B1(net40),
    .B2(net83),
    .X(_00519_));
 sky130_fd_sc_hd__xnor2_1 _07429_ (.A(net186),
    .B(_00519_),
    .Y(_00520_));
 sky130_fd_sc_hd__o22a_1 _07430_ (.A1(net55),
    .A2(net132),
    .B1(net170),
    .B2(net52),
    .X(_00521_));
 sky130_fd_sc_hd__xnor2_1 _07431_ (.A(net194),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__nor2_1 _07432_ (.A(_00520_),
    .B(_00522_),
    .Y(_00523_));
 sky130_fd_sc_hd__and2_1 _07433_ (.A(_00520_),
    .B(_00522_),
    .X(_00524_));
 sky130_fd_sc_hd__nor2_2 _07434_ (.A(_00523_),
    .B(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__o22a_2 _07435_ (.A1(net49),
    .A2(net130),
    .B1(net128),
    .B2(net46),
    .X(_00526_));
 sky130_fd_sc_hd__xnor2_4 _07436_ (.A(net167),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__xnor2_4 _07437_ (.A(_00525_),
    .B(_00527_),
    .Y(_00528_));
 sky130_fd_sc_hd__xnor2_4 _07438_ (.A(_00505_),
    .B(_00518_),
    .Y(_00529_));
 sky130_fd_sc_hd__a32o_2 _07439_ (.A1(_00503_),
    .A2(_00504_),
    .A3(_00518_),
    .B1(_00528_),
    .B2(_00529_),
    .X(_00530_));
 sky130_fd_sc_hd__o22a_1 _07440_ (.A1(net180),
    .A2(net16),
    .B1(net37),
    .B2(net144),
    .X(_00531_));
 sky130_fd_sc_hd__xnor2_1 _07441_ (.A(net78),
    .B(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__o22a_1 _07442_ (.A1(net23),
    .A2(net142),
    .B1(net140),
    .B2(net70),
    .X(_00533_));
 sky130_fd_sc_hd__xor2_1 _07443_ (.A(net110),
    .B(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__or2_1 _07444_ (.A(_00532_),
    .B(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__nand2_1 _07445_ (.A(_00532_),
    .B(_00534_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(_00535_),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__o22a_1 _07447_ (.A1(net30),
    .A2(net148),
    .B1(net146),
    .B2(net28),
    .X(_00538_));
 sky130_fd_sc_hd__xnor2_1 _07448_ (.A(_06524_),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__xnor2_1 _07449_ (.A(_00537_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__o21ba_1 _07450_ (.A1(_00424_),
    .A2(_00427_),
    .B1_N(_00423_),
    .X(_00541_));
 sky130_fd_sc_hd__nand2b_1 _07451_ (.A_N(_00541_),
    .B(_00475_),
    .Y(_00542_));
 sky130_fd_sc_hd__o21ai_1 _07452_ (.A1(_00448_),
    .A2(_00450_),
    .B1(_00446_),
    .Y(_00543_));
 sky130_fd_sc_hd__xnor2_1 _07453_ (.A(_00475_),
    .B(_00541_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand2_1 _07454_ (.A(_00543_),
    .B(_00544_),
    .Y(_00545_));
 sky130_fd_sc_hd__a21o_1 _07455_ (.A1(_00542_),
    .A2(_00545_),
    .B1(_00540_),
    .X(_00546_));
 sky130_fd_sc_hd__nand3_1 _07456_ (.A(_00540_),
    .B(_00542_),
    .C(_00545_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_2 _07457_ (.A(_00546_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2b_1 _07458_ (.A_N(_00548_),
    .B(_00530_),
    .Y(_00549_));
 sky130_fd_sc_hd__xnor2_4 _07459_ (.A(_00530_),
    .B(_00548_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _07460_ (.A(_00499_),
    .B(_00503_),
    .Y(_00551_));
 sky130_fd_sc_hd__o22a_1 _07461_ (.A1(net96),
    .A2(net20),
    .B1(net64),
    .B2(net89),
    .X(_00552_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(net93),
    .B(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__o22a_1 _07463_ (.A1(net98),
    .A2(net66),
    .B1(_00191_),
    .B2(net22),
    .X(_00554_));
 sky130_fd_sc_hd__xnor2_1 _07464_ (.A(net103),
    .B(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__and2_1 _07465_ (.A(_00553_),
    .B(_00555_),
    .X(_00556_));
 sky130_fd_sc_hd__o21ba_1 _07466_ (.A1(_00524_),
    .A2(_00527_),
    .B1_N(_00523_),
    .X(_00557_));
 sky130_fd_sc_hd__nand2b_1 _07467_ (.A_N(_00557_),
    .B(_00556_),
    .Y(_00558_));
 sky130_fd_sc_hd__xnor2_1 _07468_ (.A(_00556_),
    .B(_00557_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _07469_ (.A(_00551_),
    .B(_00559_),
    .Y(_00560_));
 sky130_fd_sc_hd__or2_1 _07470_ (.A(_00551_),
    .B(_00559_),
    .X(_00561_));
 sky130_fd_sc_hd__and2_1 _07471_ (.A(_00560_),
    .B(_00561_),
    .X(_00562_));
 sky130_fd_sc_hd__o22a_1 _07472_ (.A1(net49),
    .A2(net83),
    .B1(net40),
    .B2(net88),
    .X(_00563_));
 sky130_fd_sc_hd__xnor2_1 _07473_ (.A(net186),
    .B(_00563_),
    .Y(_00564_));
 sky130_fd_sc_hd__o22a_1 _07474_ (.A1(net52),
    .A2(net132),
    .B1(net170),
    .B2(net63),
    .X(_00565_));
 sky130_fd_sc_hd__xnor2_1 _07475_ (.A(net194),
    .B(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__nor2_1 _07476_ (.A(_00564_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__and2_1 _07477_ (.A(_00564_),
    .B(_00566_),
    .X(_00568_));
 sky130_fd_sc_hd__nor2_1 _07478_ (.A(_00567_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__o22a_1 _07479_ (.A1(net46),
    .A2(net130),
    .B1(net128),
    .B2(net55),
    .X(_00570_));
 sky130_fd_sc_hd__xnor2_2 _07480_ (.A(net167),
    .B(_00570_),
    .Y(_00571_));
 sky130_fd_sc_hd__xnor2_2 _07481_ (.A(_00569_),
    .B(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__o22a_1 _07482_ (.A1(net125),
    .A2(net81),
    .B1(net43),
    .B2(net121),
    .X(_00573_));
 sky130_fd_sc_hd__xnor2_1 _07483_ (.A(net153),
    .B(_00573_),
    .Y(_00574_));
 sky130_fd_sc_hd__o22a_1 _07484_ (.A1(_06509_),
    .A2(net68),
    .B1(_00167_),
    .B2(_06491_),
    .X(_00575_));
 sky130_fd_sc_hd__xnor2_1 _07485_ (.A(_00152_),
    .B(_00575_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2b_1 _07486_ (.A_N(_00574_),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__xor2_1 _07487_ (.A(_00574_),
    .B(_00576_),
    .X(_00578_));
 sky130_fd_sc_hd__o22a_1 _07488_ (.A1(_06494_),
    .A2(net74),
    .B1(net115),
    .B2(net86),
    .X(_00579_));
 sky130_fd_sc_hd__xnor2_1 _07489_ (.A(net150),
    .B(_00579_),
    .Y(_00580_));
 sky130_fd_sc_hd__or2_1 _07490_ (.A(_00578_),
    .B(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__nand2_1 _07491_ (.A(_00578_),
    .B(_00580_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(_00581_),
    .B(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__o22a_1 _07493_ (.A1(net178),
    .A2(net19),
    .B1(net14),
    .B2(net175),
    .X(_00584_));
 sky130_fd_sc_hd__xnor2_2 _07494_ (.A(_00210_),
    .B(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__o22a_1 _07495_ (.A1(net60),
    .A2(net134),
    .B1(net172),
    .B2(net57),
    .X(_00586_));
 sky130_fd_sc_hd__xnor2_2 _07496_ (.A(_00249_),
    .B(_00586_),
    .Y(_00587_));
 sky130_fd_sc_hd__a21oi_2 _07497_ (.A1(net306),
    .A2(_00510_),
    .B1(net260),
    .Y(_00588_));
 sky130_fd_sc_hd__and2_1 _07498_ (.A(_00587_),
    .B(_00588_),
    .X(_00589_));
 sky130_fd_sc_hd__xor2_2 _07499_ (.A(_00587_),
    .B(_00588_),
    .X(_00590_));
 sky130_fd_sc_hd__xor2_2 _07500_ (.A(_00585_),
    .B(_00590_),
    .X(_00591_));
 sky130_fd_sc_hd__xnor2_2 _07501_ (.A(_00583_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__xor2_2 _07502_ (.A(_00572_),
    .B(_00592_),
    .X(_00593_));
 sky130_fd_sc_hd__or3_2 _07503_ (.A(reg1_val[29]),
    .B(reg1_val[30]),
    .C(_00345_),
    .X(_00594_));
 sky130_fd_sc_hd__a21boi_4 _07504_ (.A1(instruction[7]),
    .A2(_00594_),
    .B1_N(reg1_val[31]),
    .Y(_00595_));
 sky130_fd_sc_hd__a21bo_4 _07505_ (.A1(instruction[7]),
    .A2(_00594_),
    .B1_N(reg1_val[31]),
    .X(_00596_));
 sky130_fd_sc_hd__nand2_1 _07506_ (.A(net224),
    .B(net35),
    .Y(_00597_));
 sky130_fd_sc_hd__a21oi_1 _07507_ (.A1(_00508_),
    .A2(_00517_),
    .B1(_00516_),
    .Y(_00598_));
 sky130_fd_sc_hd__or3_2 _07508_ (.A(net77),
    .B(_00456_),
    .C(net33),
    .X(_00599_));
 sky130_fd_sc_hd__or3b_2 _07509_ (.A(_00348_),
    .B(net32),
    .C_N(_00456_),
    .X(_00600_));
 sky130_fd_sc_hd__and2_1 _07510_ (.A(_00599_),
    .B(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__o22a_1 _07511_ (.A1(net183),
    .A2(net11),
    .B1(net5),
    .B2(net185),
    .X(_00602_));
 sky130_fd_sc_hd__xnor2_1 _07512_ (.A(net35),
    .B(_00602_),
    .Y(_00603_));
 sky130_fd_sc_hd__and2b_1 _07513_ (.A_N(_00598_),
    .B(_00603_),
    .X(_00604_));
 sky130_fd_sc_hd__xnor2_1 _07514_ (.A(_00598_),
    .B(_00603_),
    .Y(_00605_));
 sky130_fd_sc_hd__xnor2_1 _07515_ (.A(_00597_),
    .B(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _07516_ (.A(_00593_),
    .B(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__xor2_1 _07517_ (.A(_00593_),
    .B(_00606_),
    .X(_00608_));
 sky130_fd_sc_hd__nand2_1 _07518_ (.A(_00562_),
    .B(_00608_),
    .Y(_00609_));
 sky130_fd_sc_hd__or2_1 _07519_ (.A(_00562_),
    .B(_00608_),
    .X(_00610_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(_00609_),
    .B(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hd__o22a_1 _07521_ (.A1(net28),
    .A2(net148),
    .B1(net144),
    .B2(net30),
    .X(_00612_));
 sky130_fd_sc_hd__xnor2_1 _07522_ (.A(_06523_),
    .B(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__o22a_1 _07523_ (.A1(net25),
    .A2(net140),
    .B1(net137),
    .B2(net72),
    .X(_00614_));
 sky130_fd_sc_hd__xnor2_1 _07524_ (.A(_06543_),
    .B(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hd__and2_1 _07525_ (.A(_00613_),
    .B(_00615_),
    .X(_00616_));
 sky130_fd_sc_hd__nor2_1 _07526_ (.A(_00613_),
    .B(_00615_),
    .Y(_00617_));
 sky130_fd_sc_hd__nor2_1 _07527_ (.A(_00616_),
    .B(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__o22a_1 _07528_ (.A1(net146),
    .A2(net23),
    .B1(net70),
    .B2(net142),
    .X(_00619_));
 sky130_fd_sc_hd__xor2_1 _07529_ (.A(net110),
    .B(_00619_),
    .X(_00620_));
 sky130_fd_sc_hd__o21bai_2 _07530_ (.A1(_00617_),
    .A2(_00620_),
    .B1_N(_00616_),
    .Y(_00621_));
 sky130_fd_sc_hd__a21o_1 _07531_ (.A1(_00188_),
    .A2(_00189_),
    .B1(net89),
    .X(_00622_));
 sky130_fd_sc_hd__or2_1 _07532_ (.A(net117),
    .B(net64),
    .X(_00623_));
 sky130_fd_sc_hd__and3_1 _07533_ (.A(net93),
    .B(_00622_),
    .C(_00623_),
    .X(_00624_));
 sky130_fd_sc_hd__a21oi_1 _07534_ (.A1(_00622_),
    .A2(_00623_),
    .B1(net93),
    .Y(_00625_));
 sky130_fd_sc_hd__a21o_1 _07535_ (.A1(_06552_),
    .A2(_06553_),
    .B1(net137),
    .X(_00626_));
 sky130_fd_sc_hd__or2_1 _07536_ (.A(_06558_),
    .B(net135),
    .X(_00627_));
 sky130_fd_sc_hd__and3_1 _07537_ (.A(net107),
    .B(_00626_),
    .C(_00627_),
    .X(_00628_));
 sky130_fd_sc_hd__a21oi_1 _07538_ (.A1(_00626_),
    .A2(_00627_),
    .B1(net107),
    .Y(_00629_));
 sky130_fd_sc_hd__o22a_1 _07539_ (.A1(_00624_),
    .A2(_00625_),
    .B1(_00628_),
    .B2(_00629_),
    .X(_00630_));
 sky130_fd_sc_hd__or4_1 _07540_ (.A(_00624_),
    .B(_00625_),
    .C(_00628_),
    .D(_00629_),
    .X(_00631_));
 sky130_fd_sc_hd__nand2b_2 _07541_ (.A_N(_00630_),
    .B(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__o22a_1 _07542_ (.A1(net98),
    .A2(net22),
    .B1(net66),
    .B2(_00166_),
    .X(_00633_));
 sky130_fd_sc_hd__xnor2_2 _07543_ (.A(net103),
    .B(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hd__and2b_1 _07544_ (.A_N(_00632_),
    .B(_00634_),
    .X(_00635_));
 sky130_fd_sc_hd__xnor2_2 _07545_ (.A(_00632_),
    .B(_00634_),
    .Y(_00636_));
 sky130_fd_sc_hd__a21o_2 _07546_ (.A1(_00431_),
    .A2(_00440_),
    .B1(_00439_),
    .X(_00637_));
 sky130_fd_sc_hd__o22a_2 _07547_ (.A1(net183),
    .A2(net16),
    .B1(net37),
    .B2(net180),
    .X(_00638_));
 sky130_fd_sc_hd__xnor2_4 _07548_ (.A(net78),
    .B(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__and2b_1 _07549_ (.A_N(_00639_),
    .B(_00637_),
    .X(_00640_));
 sky130_fd_sc_hd__o22a_2 _07550_ (.A1(net185),
    .A2(net11),
    .B1(net5),
    .B2(net229),
    .X(_00641_));
 sky130_fd_sc_hd__xnor2_4 _07551_ (.A(net35),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__xnor2_4 _07552_ (.A(_00637_),
    .B(_00639_),
    .Y(_00643_));
 sky130_fd_sc_hd__a21oi_2 _07553_ (.A1(_00642_),
    .A2(_00643_),
    .B1(_00640_),
    .Y(_00644_));
 sky130_fd_sc_hd__and2b_1 _07554_ (.A_N(_00644_),
    .B(_00636_),
    .X(_00645_));
 sky130_fd_sc_hd__xnor2_2 _07555_ (.A(_00636_),
    .B(_00644_),
    .Y(_00646_));
 sky130_fd_sc_hd__xnor2_1 _07556_ (.A(_00621_),
    .B(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hd__nor2_1 _07557_ (.A(_00611_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _07558_ (.A(_00611_),
    .B(_00647_),
    .Y(_00649_));
 sky130_fd_sc_hd__and2b_1 _07559_ (.A_N(_00648_),
    .B(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__xor2_4 _07560_ (.A(_00550_),
    .B(_00650_),
    .X(_00651_));
 sky130_fd_sc_hd__or2_1 _07561_ (.A(_00543_),
    .B(_00544_),
    .X(_00652_));
 sky130_fd_sc_hd__and2_2 _07562_ (.A(_00545_),
    .B(_00652_),
    .X(_00653_));
 sky130_fd_sc_hd__xnor2_4 _07563_ (.A(_00528_),
    .B(_00529_),
    .Y(_00654_));
 sky130_fd_sc_hd__xnor2_4 _07564_ (.A(_00642_),
    .B(_00643_),
    .Y(_00655_));
 sky130_fd_sc_hd__nor2_1 _07565_ (.A(_00654_),
    .B(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hd__xor2_4 _07566_ (.A(_00654_),
    .B(_00655_),
    .X(_00657_));
 sky130_fd_sc_hd__xor2_2 _07567_ (.A(_00653_),
    .B(_00657_),
    .X(_00658_));
 sky130_fd_sc_hd__nor2_1 _07568_ (.A(_00553_),
    .B(_00555_),
    .Y(_00659_));
 sky130_fd_sc_hd__nor2_2 _07569_ (.A(_00556_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__mux2_2 _07570_ (.A0(_00595_),
    .A1(_00461_),
    .S(_00458_),
    .X(_00661_));
 sky130_fd_sc_hd__xor2_1 _07571_ (.A(_00660_),
    .B(_00661_),
    .X(_00662_));
 sky130_fd_sc_hd__o21a_1 _07572_ (.A1(_00407_),
    .A2(_00412_),
    .B1(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__nor3_1 _07573_ (.A(_00407_),
    .B(_00412_),
    .C(_00662_),
    .Y(_00664_));
 sky130_fd_sc_hd__or2_2 _07574_ (.A(_00663_),
    .B(_00664_),
    .X(_00665_));
 sky130_fd_sc_hd__inv_2 _07575_ (.A(_00665_),
    .Y(_00666_));
 sky130_fd_sc_hd__o21ai_4 _07576_ (.A1(_00429_),
    .A2(_00453_),
    .B1(_00452_),
    .Y(_00667_));
 sky130_fd_sc_hd__xnor2_1 _07577_ (.A(_00618_),
    .B(_00620_),
    .Y(_00668_));
 sky130_fd_sc_hd__o21a_1 _07578_ (.A1(_00464_),
    .A2(_00466_),
    .B1(_00668_),
    .X(_00669_));
 sky130_fd_sc_hd__nor3_1 _07579_ (.A(_00464_),
    .B(_00466_),
    .C(_00668_),
    .Y(_00670_));
 sky130_fd_sc_hd__nor2_2 _07580_ (.A(_00669_),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__xnor2_4 _07581_ (.A(_00667_),
    .B(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__xnor2_2 _07582_ (.A(_00658_),
    .B(_00665_),
    .Y(_00673_));
 sky130_fd_sc_hd__and2b_1 _07583_ (.A_N(_00672_),
    .B(_00673_),
    .X(_00674_));
 sky130_fd_sc_hd__a21oi_2 _07584_ (.A1(_00658_),
    .A2(_00666_),
    .B1(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__a21o_1 _07585_ (.A1(_00667_),
    .A2(_00671_),
    .B1(_00669_),
    .X(_00676_));
 sky130_fd_sc_hd__a21oi_4 _07586_ (.A1(_00653_),
    .A2(_00657_),
    .B1(_00656_),
    .Y(_00677_));
 sky130_fd_sc_hd__a21oi_4 _07587_ (.A1(_00660_),
    .A2(_00661_),
    .B1(_00663_),
    .Y(_00678_));
 sky130_fd_sc_hd__nor2_1 _07588_ (.A(_00677_),
    .B(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hd__xor2_4 _07589_ (.A(_00677_),
    .B(_00678_),
    .X(_00680_));
 sky130_fd_sc_hd__xnor2_2 _07590_ (.A(_00676_),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__a21bo_1 _07591_ (.A1(_00418_),
    .A2(_00484_),
    .B1_N(_00483_),
    .X(_00682_));
 sky130_fd_sc_hd__nand2b_1 _07592_ (.A_N(_00681_),
    .B(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__xnor2_2 _07593_ (.A(_00681_),
    .B(_00682_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand2b_1 _07594_ (.A_N(_00675_),
    .B(_00684_),
    .Y(_00685_));
 sky130_fd_sc_hd__xnor2_2 _07595_ (.A(_00675_),
    .B(_00684_),
    .Y(_00686_));
 sky130_fd_sc_hd__and2_1 _07596_ (.A(_00651_),
    .B(_00686_),
    .X(_00687_));
 sky130_fd_sc_hd__xor2_4 _07597_ (.A(_00651_),
    .B(_00686_),
    .X(_00688_));
 sky130_fd_sc_hd__xnor2_4 _07598_ (.A(_00494_),
    .B(_00688_),
    .Y(_00689_));
 sky130_fd_sc_hd__xnor2_4 _07599_ (.A(_00672_),
    .B(_00673_),
    .Y(_00690_));
 sky130_fd_sc_hd__xnor2_2 _07600_ (.A(_00491_),
    .B(_00492_),
    .Y(_00691_));
 sky130_fd_sc_hd__and2_1 _07601_ (.A(_00690_),
    .B(_00691_),
    .X(_00692_));
 sky130_fd_sc_hd__xnor2_4 _07602_ (.A(_00399_),
    .B(_00400_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _07603_ (.A(_00267_),
    .B(_00271_),
    .Y(_00694_));
 sky130_fd_sc_hd__nand2_1 _07604_ (.A(_00272_),
    .B(_00694_),
    .Y(_00695_));
 sky130_fd_sc_hd__o22a_1 _07605_ (.A1(net98),
    .A2(net94),
    .B1(net135),
    .B2(net69),
    .X(_00696_));
 sky130_fd_sc_hd__xnor2_1 _07606_ (.A(net100),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__o32a_1 _07607_ (.A1(net146),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net66),
    .B2(net142),
    .X(_00698_));
 sky130_fd_sc_hd__xnor2_1 _07608_ (.A(net102),
    .B(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _07609_ (.A(_00697_),
    .B(_00699_),
    .Y(_00700_));
 sky130_fd_sc_hd__xor2_1 _07610_ (.A(_00697_),
    .B(_00699_),
    .X(_00701_));
 sky130_fd_sc_hd__o22a_1 _07611_ (.A1(net140),
    .A2(net20),
    .B1(net64),
    .B2(net137),
    .X(_00702_));
 sky130_fd_sc_hd__xnor2_1 _07612_ (.A(net91),
    .B(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _07613_ (.A(_00701_),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__a21oi_1 _07614_ (.A1(_00700_),
    .A2(_00704_),
    .B1(_00695_),
    .Y(_00705_));
 sky130_fd_sc_hd__o22a_1 _07615_ (.A1(net123),
    .A2(net88),
    .B1(net83),
    .B2(net119),
    .X(_00706_));
 sky130_fd_sc_hd__xnor2_1 _07616_ (.A(net186),
    .B(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__o22a_1 _07617_ (.A1(net74),
    .A2(net96),
    .B1(net89),
    .B2(net115),
    .X(_00708_));
 sky130_fd_sc_hd__xnor2_1 _07618_ (.A(net149),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__o22a_1 _07619_ (.A1(net125),
    .A2(net117),
    .B1(net113),
    .B2(net121),
    .X(_00710_));
 sky130_fd_sc_hd__xnor2_1 _07620_ (.A(net152),
    .B(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__xnor2_1 _07621_ (.A(_00707_),
    .B(_00709_),
    .Y(_00712_));
 sky130_fd_sc_hd__or2_1 _07622_ (.A(_00711_),
    .B(_00712_),
    .X(_00713_));
 sky130_fd_sc_hd__o21ai_1 _07623_ (.A1(_00707_),
    .A2(_00709_),
    .B1(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__and3_1 _07624_ (.A(_00695_),
    .B(_00700_),
    .C(_00704_),
    .X(_00715_));
 sky130_fd_sc_hd__or2_1 _07625_ (.A(_00705_),
    .B(_00715_),
    .X(_00716_));
 sky130_fd_sc_hd__and2b_1 _07626_ (.A_N(_00716_),
    .B(_00714_),
    .X(_00717_));
 sky130_fd_sc_hd__or2_1 _07627_ (.A(_00705_),
    .B(_00717_),
    .X(_00718_));
 sky130_fd_sc_hd__xnor2_2 _07628_ (.A(_00393_),
    .B(_00394_),
    .Y(_00719_));
 sky130_fd_sc_hd__xor2_2 _07629_ (.A(_06562_),
    .B(_00145_),
    .X(_00720_));
 sky130_fd_sc_hd__and2b_1 _07630_ (.A_N(_00719_),
    .B(_00720_),
    .X(_00721_));
 sky130_fd_sc_hd__xnor2_2 _07631_ (.A(_00719_),
    .B(_00720_),
    .Y(_00722_));
 sky130_fd_sc_hd__o21bai_1 _07632_ (.A1(_00378_),
    .A2(_00382_),
    .B1_N(_00373_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_1 _07633_ (.A(_00383_),
    .B(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__a21oi_1 _07634_ (.A1(_00722_),
    .A2(_00724_),
    .B1(_00721_),
    .Y(_00725_));
 sky130_fd_sc_hd__o21ba_1 _07635_ (.A1(_00705_),
    .A2(_00717_),
    .B1_N(_00725_),
    .X(_00726_));
 sky130_fd_sc_hd__or2_1 _07636_ (.A(_00184_),
    .B(_00194_),
    .X(_00727_));
 sky130_fd_sc_hd__and2_1 _07637_ (.A(_00195_),
    .B(_00727_),
    .X(_00728_));
 sky130_fd_sc_hd__o22a_1 _07638_ (.A1(net229),
    .A2(net30),
    .B1(net28),
    .B2(net185),
    .X(_00729_));
 sky130_fd_sc_hd__xnor2_1 _07639_ (.A(net112),
    .B(_00729_),
    .Y(_00730_));
 sky130_fd_sc_hd__o22a_1 _07640_ (.A1(net148),
    .A2(net73),
    .B1(net144),
    .B2(net26),
    .X(_00731_));
 sky130_fd_sc_hd__xnor2_1 _07641_ (.A(net106),
    .B(_00731_),
    .Y(_00732_));
 sky130_fd_sc_hd__xor2_1 _07642_ (.A(_00730_),
    .B(_00732_),
    .X(_00733_));
 sky130_fd_sc_hd__o22a_1 _07643_ (.A1(net183),
    .A2(net24),
    .B1(net71),
    .B2(net180),
    .X(_00734_));
 sky130_fd_sc_hd__xnor2_1 _07644_ (.A(net110),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__and2_1 _07645_ (.A(_00733_),
    .B(_00735_),
    .X(_00736_));
 sky130_fd_sc_hd__a21o_1 _07646_ (.A1(_00730_),
    .A2(_00732_),
    .B1(_00736_),
    .X(_00737_));
 sky130_fd_sc_hd__xnor2_1 _07647_ (.A(_00380_),
    .B(_00381_),
    .Y(_00738_));
 sky130_fd_sc_hd__o22a_1 _07648_ (.A1(net171),
    .A2(net47),
    .B1(net38),
    .B2(net133),
    .X(_00739_));
 sky130_fd_sc_hd__xnor2_1 _07649_ (.A(net210),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__o22a_1 _07650_ (.A1(net306),
    .A2(net62),
    .B1(net257),
    .B2(net50),
    .X(_00741_));
 sky130_fd_sc_hd__xnor2_1 _07651_ (.A(net258),
    .B(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__nor2_1 _07652_ (.A(_00740_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__o22a_1 _07653_ (.A1(net173),
    .A2(net53),
    .B1(net44),
    .B2(net176),
    .X(_00744_));
 sky130_fd_sc_hd__xnor2_1 _07654_ (.A(net212),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__inv_2 _07655_ (.A(_00745_),
    .Y(_00746_));
 sky130_fd_sc_hd__xor2_1 _07656_ (.A(_00740_),
    .B(_00742_),
    .X(_00747_));
 sky130_fd_sc_hd__a21oi_1 _07657_ (.A1(_00746_),
    .A2(_00747_),
    .B1(_00743_),
    .Y(_00748_));
 sky130_fd_sc_hd__nand2b_1 _07658_ (.A_N(_00748_),
    .B(_00738_),
    .Y(_00749_));
 sky130_fd_sc_hd__o22a_1 _07659_ (.A1(net132),
    .A2(net80),
    .B1(net41),
    .B2(net170),
    .X(_00750_));
 sky130_fd_sc_hd__xnor2_1 _07660_ (.A(net194),
    .B(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__o22a_1 _07661_ (.A1(net120),
    .A2(net130),
    .B1(net128),
    .B2(net85),
    .X(_00752_));
 sky130_fd_sc_hd__xnor2_1 _07662_ (.A(net167),
    .B(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__nor2_1 _07663_ (.A(_00751_),
    .B(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__xnor2_1 _07664_ (.A(_00738_),
    .B(_00748_),
    .Y(_00755_));
 sky130_fd_sc_hd__a21bo_1 _07665_ (.A1(_00754_),
    .A2(_00755_),
    .B1_N(_00749_),
    .X(_00756_));
 sky130_fd_sc_hd__xnor2_1 _07666_ (.A(_00728_),
    .B(_00737_),
    .Y(_00757_));
 sky130_fd_sc_hd__and2b_1 _07667_ (.A_N(_00757_),
    .B(_00756_),
    .X(_00758_));
 sky130_fd_sc_hd__a21o_1 _07668_ (.A1(_00728_),
    .A2(_00737_),
    .B1(_00758_),
    .X(_00759_));
 sky130_fd_sc_hd__xnor2_2 _07669_ (.A(_00718_),
    .B(_00725_),
    .Y(_00760_));
 sky130_fd_sc_hd__a21oi_4 _07670_ (.A1(_00759_),
    .A2(_00760_),
    .B1(_00726_),
    .Y(_00761_));
 sky130_fd_sc_hd__xor2_1 _07671_ (.A(_00148_),
    .B(_00196_),
    .X(_00762_));
 sky130_fd_sc_hd__xnor2_1 _07672_ (.A(_00360_),
    .B(_00361_),
    .Y(_00763_));
 sky130_fd_sc_hd__nor2_1 _07673_ (.A(_00762_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__xnor2_4 _07674_ (.A(_00395_),
    .B(_00397_),
    .Y(_00765_));
 sky130_fd_sc_hd__and2_1 _07675_ (.A(_00762_),
    .B(_00763_),
    .X(_00766_));
 sky130_fd_sc_hd__nor2_2 _07676_ (.A(_00764_),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__a21o_1 _07677_ (.A1(_00765_),
    .A2(_00767_),
    .B1(_00764_),
    .X(_00768_));
 sky130_fd_sc_hd__xnor2_2 _07678_ (.A(_00693_),
    .B(_00761_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2b_1 _07679_ (.A_N(_00769_),
    .B(_00768_),
    .Y(_00770_));
 sky130_fd_sc_hd__o21ai_4 _07680_ (.A1(_00693_),
    .A2(_00761_),
    .B1(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__xor2_4 _07681_ (.A(_00690_),
    .B(_00691_),
    .X(_00772_));
 sky130_fd_sc_hd__a21oi_4 _07682_ (.A1(_00771_),
    .A2(_00772_),
    .B1(_00692_),
    .Y(_00773_));
 sky130_fd_sc_hd__or2_1 _07683_ (.A(_00689_),
    .B(_00773_),
    .X(_00774_));
 sky130_fd_sc_hd__and2_1 _07684_ (.A(_00689_),
    .B(_00773_),
    .X(_00775_));
 sky130_fd_sc_hd__xnor2_4 _07685_ (.A(_00689_),
    .B(_00773_),
    .Y(_00776_));
 sky130_fd_sc_hd__o22a_1 _07686_ (.A1(net26),
    .A2(net179),
    .B1(net143),
    .B2(net73),
    .X(_00777_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(net106),
    .B(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__nor2_1 _07688_ (.A(net225),
    .B(net28),
    .Y(_00779_));
 sky130_fd_sc_hd__xnor2_1 _07689_ (.A(_06524_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__and2_1 _07690_ (.A(_00778_),
    .B(_00780_),
    .X(_00781_));
 sky130_fd_sc_hd__xnor2_1 _07691_ (.A(_00778_),
    .B(_00780_),
    .Y(_00782_));
 sky130_fd_sc_hd__o22a_1 _07692_ (.A1(net185),
    .A2(net24),
    .B1(net71),
    .B2(net181),
    .X(_00783_));
 sky130_fd_sc_hd__xnor2_1 _07693_ (.A(net110),
    .B(_00783_),
    .Y(_00784_));
 sky130_fd_sc_hd__and2b_1 _07694_ (.A_N(_00782_),
    .B(_00784_),
    .X(_00785_));
 sky130_fd_sc_hd__and2b_1 _07695_ (.A_N(_00784_),
    .B(_00782_),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _07696_ (.A(_00785_),
    .B(_00786_),
    .X(_00787_));
 sky130_fd_sc_hd__inv_2 _07697_ (.A(_00787_),
    .Y(_00788_));
 sky130_fd_sc_hd__o22a_1 _07698_ (.A1(net257),
    .A2(net53),
    .B1(net51),
    .B2(net306),
    .X(_00789_));
 sky130_fd_sc_hd__xnor2_1 _07699_ (.A(net258),
    .B(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__o22a_1 _07700_ (.A1(net176),
    .A2(net47),
    .B1(net44),
    .B2(net173),
    .X(_00791_));
 sky130_fd_sc_hd__xnor2_1 _07701_ (.A(net212),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__or2_2 _07702_ (.A(_00790_),
    .B(_00792_),
    .X(_00793_));
 sky130_fd_sc_hd__xnor2_1 _07703_ (.A(_00745_),
    .B(_00747_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _07704_ (.A(net111),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__xnor2_1 _07705_ (.A(net111),
    .B(_00794_),
    .Y(_00796_));
 sky130_fd_sc_hd__xnor2_1 _07706_ (.A(_00793_),
    .B(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__o22a_1 _07707_ (.A1(net69),
    .A2(net137),
    .B1(net135),
    .B2(net95),
    .X(_00798_));
 sky130_fd_sc_hd__xnor2_1 _07708_ (.A(net101),
    .B(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__o32a_1 _07709_ (.A1(net148),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net67),
    .B2(net146),
    .X(_00800_));
 sky130_fd_sc_hd__xnor2_1 _07710_ (.A(net104),
    .B(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__and2_1 _07711_ (.A(_00799_),
    .B(_00801_),
    .X(_00802_));
 sky130_fd_sc_hd__nor2_1 _07712_ (.A(_00799_),
    .B(_00801_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_1 _07713_ (.A(_00802_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hd__o22a_1 _07714_ (.A1(_00171_),
    .A2(net21),
    .B1(net65),
    .B2(_00180_),
    .X(_00805_));
 sky130_fd_sc_hd__xnor2_1 _07715_ (.A(_00174_),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__xor2_1 _07716_ (.A(_00804_),
    .B(_00806_),
    .X(_00807_));
 sky130_fd_sc_hd__and2b_1 _07717_ (.A_N(_00797_),
    .B(_00807_),
    .X(_00808_));
 sky130_fd_sc_hd__xnor2_1 _07718_ (.A(_00797_),
    .B(_00807_),
    .Y(_00809_));
 sky130_fd_sc_hd__xnor2_1 _07719_ (.A(_00787_),
    .B(_00809_),
    .Y(_00810_));
 sky130_fd_sc_hd__o22a_1 _07720_ (.A1(net133),
    .A2(net41),
    .B1(net38),
    .B2(net171),
    .X(_00811_));
 sky130_fd_sc_hd__xnor2_1 _07721_ (.A(net210),
    .B(_00811_),
    .Y(_00812_));
 sky130_fd_sc_hd__o22a_1 _07722_ (.A1(net124),
    .A2(net130),
    .B1(net128),
    .B2(net120),
    .X(_00813_));
 sky130_fd_sc_hd__xnor2_1 _07723_ (.A(net166),
    .B(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__or2_1 _07724_ (.A(_00812_),
    .B(_00814_),
    .X(_00815_));
 sky130_fd_sc_hd__o22a_1 _07725_ (.A1(net131),
    .A2(net84),
    .B1(net79),
    .B2(net169),
    .X(_00816_));
 sky130_fd_sc_hd__xnor2_1 _07726_ (.A(net193),
    .B(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hd__xnor2_1 _07727_ (.A(_00812_),
    .B(_00814_),
    .Y(_00818_));
 sky130_fd_sc_hd__o21ai_1 _07728_ (.A1(_00817_),
    .A2(_00818_),
    .B1(_00815_),
    .Y(_00819_));
 sky130_fd_sc_hd__and2_1 _07729_ (.A(_00751_),
    .B(_00753_),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _07730_ (.A(_00754_),
    .B(_00820_),
    .X(_00821_));
 sky130_fd_sc_hd__o22a_1 _07731_ (.A1(net118),
    .A2(net87),
    .B1(net82),
    .B2(net114),
    .X(_00822_));
 sky130_fd_sc_hd__xnor2_1 _07732_ (.A(net187),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__o22a_1 _07733_ (.A1(net116),
    .A2(net99),
    .B1(net136),
    .B2(net75),
    .X(_00824_));
 sky130_fd_sc_hd__xnor2_1 _07734_ (.A(net150),
    .B(_00824_),
    .Y(_00825_));
 sky130_fd_sc_hd__or2_1 _07735_ (.A(_00823_),
    .B(_00825_),
    .X(_00826_));
 sky130_fd_sc_hd__o22a_1 _07736_ (.A1(net126),
    .A2(net97),
    .B1(net90),
    .B2(net122),
    .X(_00827_));
 sky130_fd_sc_hd__xnor2_1 _07737_ (.A(net154),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__xnor2_1 _07738_ (.A(_00823_),
    .B(_00825_),
    .Y(_00829_));
 sky130_fd_sc_hd__or2_1 _07739_ (.A(_00828_),
    .B(_00829_),
    .X(_00830_));
 sky130_fd_sc_hd__a21oi_1 _07740_ (.A1(_00826_),
    .A2(_00830_),
    .B1(_00821_),
    .Y(_00831_));
 sky130_fd_sc_hd__and3_1 _07741_ (.A(_00821_),
    .B(_00826_),
    .C(_00830_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _07742_ (.A(_00831_),
    .B(_00832_),
    .X(_00833_));
 sky130_fd_sc_hd__and2b_1 _07743_ (.A_N(_00833_),
    .B(_00819_),
    .X(_00834_));
 sky130_fd_sc_hd__xnor2_1 _07744_ (.A(_00819_),
    .B(_00833_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(_00810_),
    .B(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__xnor2_1 _07746_ (.A(_00810_),
    .B(_00835_),
    .Y(_00837_));
 sky130_fd_sc_hd__o22a_1 _07747_ (.A1(_04428_),
    .A2(net53),
    .B1(net44),
    .B2(net257),
    .X(_00838_));
 sky130_fd_sc_hd__xnor2_2 _07748_ (.A(net258),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__o22a_1 _07749_ (.A1(net173),
    .A2(net47),
    .B1(net38),
    .B2(net176),
    .X(_00840_));
 sky130_fd_sc_hd__xnor2_2 _07750_ (.A(net212),
    .B(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__a21o_1 _07751_ (.A1(_06552_),
    .A2(_06553_),
    .B1(net181),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _07752_ (.A(net73),
    .B(net179),
    .X(_00843_));
 sky130_fd_sc_hd__nand3_1 _07753_ (.A(net106),
    .B(_00842_),
    .C(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__a21o_1 _07754_ (.A1(_00842_),
    .A2(_00843_),
    .B1(net106),
    .X(_00845_));
 sky130_fd_sc_hd__a211o_1 _07755_ (.A1(_00844_),
    .A2(_00845_),
    .B1(_00839_),
    .C1(_00841_),
    .X(_00846_));
 sky130_fd_sc_hd__o211ai_2 _07756_ (.A1(_00839_),
    .A2(_00841_),
    .B1(_00844_),
    .C1(_00845_),
    .Y(_00847_));
 sky130_fd_sc_hd__o22a_1 _07757_ (.A1(net225),
    .A2(net24),
    .B1(net71),
    .B2(net184),
    .X(_00848_));
 sky130_fd_sc_hd__xnor2_1 _07758_ (.A(net109),
    .B(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__and3_1 _07759_ (.A(_00846_),
    .B(_00847_),
    .C(_00849_),
    .X(_00850_));
 sky130_fd_sc_hd__a21bo_1 _07760_ (.A1(_00847_),
    .A2(_00849_),
    .B1_N(_00846_),
    .X(_00851_));
 sky130_fd_sc_hd__o22a_1 _07761_ (.A1(net122),
    .A2(net118),
    .B1(net90),
    .B2(net126),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_1 _07762_ (.A(net154),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__o22a_1 _07763_ (.A1(net114),
    .A2(net87),
    .B1(net82),
    .B2(net124),
    .X(_00854_));
 sky130_fd_sc_hd__xnor2_1 _07764_ (.A(net187),
    .B(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__o22a_1 _07765_ (.A1(net75),
    .A2(net99),
    .B1(net97),
    .B2(net116),
    .X(_00856_));
 sky130_fd_sc_hd__xnor2_1 _07766_ (.A(net150),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__or2_1 _07767_ (.A(_00855_),
    .B(_00857_),
    .X(_00858_));
 sky130_fd_sc_hd__nand2_1 _07768_ (.A(_00855_),
    .B(_00857_),
    .Y(_00859_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(_00858_),
    .B(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_00853_),
    .B(_00860_),
    .Y(_00861_));
 sky130_fd_sc_hd__o22a_1 _07771_ (.A1(net69),
    .A2(net139),
    .B1(net138),
    .B2(net95),
    .X(_00862_));
 sky130_fd_sc_hd__xnor2_1 _07772_ (.A(net101),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__o22a_1 _07773_ (.A1(net143),
    .A2(net22),
    .B1(net67),
    .B2(net147),
    .X(_00864_));
 sky130_fd_sc_hd__xnor2_1 _07774_ (.A(net104),
    .B(_00864_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _07775_ (.A(_00863_),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__xor2_1 _07776_ (.A(_00863_),
    .B(_00865_),
    .X(_00867_));
 sky130_fd_sc_hd__o22a_1 _07777_ (.A1(net145),
    .A2(net21),
    .B1(net65),
    .B2(net141),
    .X(_00868_));
 sky130_fd_sc_hd__xnor2_1 _07778_ (.A(_00174_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__nand2_1 _07779_ (.A(_00867_),
    .B(_00869_),
    .Y(_00870_));
 sky130_fd_sc_hd__a21oi_1 _07780_ (.A1(_00866_),
    .A2(_00870_),
    .B1(_00861_),
    .Y(_00871_));
 sky130_fd_sc_hd__and3_1 _07781_ (.A(_00861_),
    .B(_00866_),
    .C(_00870_),
    .X(_00872_));
 sky130_fd_sc_hd__nor2_1 _07782_ (.A(_00871_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__xnor2_1 _07783_ (.A(_00851_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__xor2_1 _07784_ (.A(_00837_),
    .B(_00874_),
    .X(_00875_));
 sky130_fd_sc_hd__o32a_1 _07785_ (.A1(net171),
    .A2(_00310_),
    .A3(_00311_),
    .B1(net79),
    .B2(net133),
    .X(_00876_));
 sky130_fd_sc_hd__xnor2_2 _07786_ (.A(net210),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__o22a_1 _07787_ (.A1(net114),
    .A2(net129),
    .B1(net127),
    .B2(net124),
    .X(_00878_));
 sky130_fd_sc_hd__xnor2_2 _07788_ (.A(net166),
    .B(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__or2_1 _07789_ (.A(_00877_),
    .B(_00879_),
    .X(_00880_));
 sky130_fd_sc_hd__xnor2_2 _07790_ (.A(_00877_),
    .B(_00879_),
    .Y(_00881_));
 sky130_fd_sc_hd__o22a_1 _07791_ (.A1(net120),
    .A2(net131),
    .B1(net169),
    .B2(net84),
    .X(_00882_));
 sky130_fd_sc_hd__xnor2_2 _07792_ (.A(net193),
    .B(_00882_),
    .Y(_00883_));
 sky130_fd_sc_hd__o21ai_2 _07793_ (.A1(_00881_),
    .A2(_00883_),
    .B1(_00880_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _07794_ (.A(_00790_),
    .B(_00792_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _07795_ (.A(_00793_),
    .B(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__o22a_1 _07796_ (.A1(net90),
    .A2(net87),
    .B1(net82),
    .B2(net118),
    .X(_00887_));
 sky130_fd_sc_hd__xnor2_1 _07797_ (.A(net187),
    .B(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__a21oi_2 _07798_ (.A1(_06504_),
    .A2(_06505_),
    .B1(net137),
    .Y(_00889_));
 sky130_fd_sc_hd__nor2_1 _07799_ (.A(net116),
    .B(net136),
    .Y(_00890_));
 sky130_fd_sc_hd__or3_1 _07800_ (.A(net150),
    .B(_00889_),
    .C(_00890_),
    .X(_00891_));
 sky130_fd_sc_hd__o21ai_1 _07801_ (.A1(_00889_),
    .A2(_00890_),
    .B1(net150),
    .Y(_00892_));
 sky130_fd_sc_hd__a21o_1 _07802_ (.A1(_00891_),
    .A2(_00892_),
    .B1(_00888_),
    .X(_00893_));
 sky130_fd_sc_hd__o22a_1 _07803_ (.A1(net126),
    .A2(net99),
    .B1(net97),
    .B2(net122),
    .X(_00894_));
 sky130_fd_sc_hd__xor2_1 _07804_ (.A(net154),
    .B(_00894_),
    .X(_00895_));
 sky130_fd_sc_hd__nand3_1 _07805_ (.A(_00888_),
    .B(_00891_),
    .C(_00892_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand3_2 _07806_ (.A(_00893_),
    .B(_00895_),
    .C(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__nand2_1 _07807_ (.A(_00893_),
    .B(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__and3_1 _07808_ (.A(_00793_),
    .B(_00885_),
    .C(_00898_),
    .X(_00899_));
 sky130_fd_sc_hd__xnor2_1 _07809_ (.A(_00886_),
    .B(_00898_),
    .Y(_00900_));
 sky130_fd_sc_hd__xnor2_1 _07810_ (.A(_00884_),
    .B(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__xor2_1 _07811_ (.A(_00867_),
    .B(_00869_),
    .X(_00902_));
 sky130_fd_sc_hd__a21oi_1 _07812_ (.A1(_00846_),
    .A2(_00847_),
    .B1(_00849_),
    .Y(_00903_));
 sky130_fd_sc_hd__xor2_1 _07813_ (.A(_00828_),
    .B(_00829_),
    .X(_00904_));
 sky130_fd_sc_hd__or3b_1 _07814_ (.A(_00850_),
    .B(_00903_),
    .C_N(_00904_),
    .X(_00905_));
 sky130_fd_sc_hd__o21bai_1 _07815_ (.A1(_00850_),
    .A2(_00903_),
    .B1_N(_00904_),
    .Y(_00906_));
 sky130_fd_sc_hd__and3_1 _07816_ (.A(_00902_),
    .B(_00905_),
    .C(_00906_),
    .X(_00907_));
 sky130_fd_sc_hd__a21oi_1 _07817_ (.A1(_00905_),
    .A2(_00906_),
    .B1(_00902_),
    .Y(_00908_));
 sky130_fd_sc_hd__or3_1 _07818_ (.A(_00901_),
    .B(_00907_),
    .C(_00908_),
    .X(_00909_));
 sky130_fd_sc_hd__nor2_1 _07819_ (.A(net225),
    .B(net71),
    .Y(_00910_));
 sky130_fd_sc_hd__a21o_1 _07820_ (.A1(_06552_),
    .A2(_06553_),
    .B1(net185),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _07821_ (.A(net181),
    .B(net73),
    .X(_00912_));
 sky130_fd_sc_hd__nand3_1 _07822_ (.A(net106),
    .B(_00911_),
    .C(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__a21o_1 _07823_ (.A1(_00911_),
    .A2(_00912_),
    .B1(net106),
    .X(_00914_));
 sky130_fd_sc_hd__and3_1 _07824_ (.A(_00910_),
    .B(_00913_),
    .C(_00914_),
    .X(_00915_));
 sky130_fd_sc_hd__o21bai_1 _07825_ (.A1(net109),
    .A2(_00910_),
    .B1_N(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hd__o22a_1 _07826_ (.A1(net69),
    .A2(net141),
    .B1(net139),
    .B2(net95),
    .X(_00917_));
 sky130_fd_sc_hd__xnor2_1 _07827_ (.A(net101),
    .B(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hd__o32a_1 _07828_ (.A1(net179),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net67),
    .B2(net143),
    .X(_00919_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(net104),
    .B(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__and2_1 _07830_ (.A(_00918_),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__xor2_1 _07831_ (.A(_00918_),
    .B(_00920_),
    .X(_00922_));
 sky130_fd_sc_hd__o22a_1 _07832_ (.A1(net147),
    .A2(net21),
    .B1(net65),
    .B2(net145),
    .X(_00923_));
 sky130_fd_sc_hd__xnor2_1 _07833_ (.A(_00174_),
    .B(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__a21o_1 _07834_ (.A1(_00922_),
    .A2(_00924_),
    .B1(_00921_),
    .X(_00925_));
 sky130_fd_sc_hd__xor2_1 _07835_ (.A(_00817_),
    .B(_00818_),
    .X(_00926_));
 sky130_fd_sc_hd__xor2_1 _07836_ (.A(_00925_),
    .B(_00926_),
    .X(_00927_));
 sky130_fd_sc_hd__and2b_1 _07837_ (.A_N(_00916_),
    .B(_00927_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_1 _07838_ (.A(_00916_),
    .B(_00927_),
    .Y(_00929_));
 sky130_fd_sc_hd__o21ai_1 _07839_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00901_),
    .Y(_00930_));
 sky130_fd_sc_hd__and3_1 _07840_ (.A(_00909_),
    .B(_00929_),
    .C(_00930_),
    .X(_00931_));
 sky130_fd_sc_hd__a21boi_1 _07841_ (.A1(_00929_),
    .A2(_00930_),
    .B1_N(_00909_),
    .Y(_00932_));
 sky130_fd_sc_hd__a21o_1 _07842_ (.A1(_00925_),
    .A2(_00926_),
    .B1(_00928_),
    .X(_00933_));
 sky130_fd_sc_hd__a21o_1 _07843_ (.A1(_00884_),
    .A2(_00900_),
    .B1(_00899_),
    .X(_00934_));
 sky130_fd_sc_hd__a21bo_1 _07844_ (.A1(_00902_),
    .A2(_00906_),
    .B1_N(_00905_),
    .X(_00935_));
 sky130_fd_sc_hd__nand2_1 _07845_ (.A(_00934_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__xor2_1 _07846_ (.A(_00934_),
    .B(_00935_),
    .X(_00937_));
 sky130_fd_sc_hd__xnor2_1 _07847_ (.A(_00933_),
    .B(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__a21o_1 _07848_ (.A1(_00893_),
    .A2(_00896_),
    .B1(_00895_),
    .X(_00939_));
 sky130_fd_sc_hd__a21oi_1 _07849_ (.A1(_00913_),
    .A2(_00914_),
    .B1(_00910_),
    .Y(_00940_));
 sky130_fd_sc_hd__o211a_1 _07850_ (.A1(_00915_),
    .A2(_00940_),
    .B1(_00939_),
    .C1(_00897_),
    .X(_00941_));
 sky130_fd_sc_hd__o211ai_1 _07851_ (.A1(_00915_),
    .A2(_00940_),
    .B1(_00939_),
    .C1(_00897_),
    .Y(_00942_));
 sky130_fd_sc_hd__a211o_1 _07852_ (.A1(_00897_),
    .A2(_00939_),
    .B1(_00940_),
    .C1(_00915_),
    .X(_00943_));
 sky130_fd_sc_hd__xor2_1 _07853_ (.A(_00922_),
    .B(_00924_),
    .X(_00944_));
 sky130_fd_sc_hd__and3_1 _07854_ (.A(_00942_),
    .B(_00943_),
    .C(_00944_),
    .X(_00945_));
 sky130_fd_sc_hd__a21o_1 _07855_ (.A1(_00943_),
    .A2(_00944_),
    .B1(_00941_),
    .X(_00946_));
 sky130_fd_sc_hd__xor2_1 _07856_ (.A(_00839_),
    .B(_00841_),
    .X(_00947_));
 sky130_fd_sc_hd__o22a_1 _07857_ (.A1(net124),
    .A2(net131),
    .B1(net169),
    .B2(net120),
    .X(_00948_));
 sky130_fd_sc_hd__xnor2_1 _07858_ (.A(net193),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__o22a_1 _07859_ (.A1(net97),
    .A2(net87),
    .B1(net82),
    .B2(net90),
    .X(_00950_));
 sky130_fd_sc_hd__xnor2_1 _07860_ (.A(net187),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nor2_1 _07861_ (.A(_00949_),
    .B(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__xor2_1 _07862_ (.A(_00949_),
    .B(_00951_),
    .X(_00953_));
 sky130_fd_sc_hd__o22a_1 _07863_ (.A1(net118),
    .A2(net129),
    .B1(net127),
    .B2(net114),
    .X(_00954_));
 sky130_fd_sc_hd__xnor2_1 _07864_ (.A(net166),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__inv_2 _07865_ (.A(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__a21o_1 _07866_ (.A1(_00953_),
    .A2(_00956_),
    .B1(_00952_),
    .X(_00957_));
 sky130_fd_sc_hd__nand2_1 _07867_ (.A(_00947_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__o22a_1 _07868_ (.A1(net133),
    .A2(net84),
    .B1(net79),
    .B2(net171),
    .X(_00959_));
 sky130_fd_sc_hd__xnor2_1 _07869_ (.A(net210),
    .B(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__o22a_1 _07870_ (.A1(net256),
    .A2(net47),
    .B1(net44),
    .B2(net305),
    .X(_00961_));
 sky130_fd_sc_hd__xnor2_1 _07871_ (.A(net258),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__or2_1 _07872_ (.A(_00960_),
    .B(_00962_),
    .X(_00963_));
 sky130_fd_sc_hd__o22a_1 _07873_ (.A1(net176),
    .A2(net41),
    .B1(net38),
    .B2(net173),
    .X(_00964_));
 sky130_fd_sc_hd__xnor2_2 _07874_ (.A(net212),
    .B(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__and2_1 _07875_ (.A(_00960_),
    .B(_00962_),
    .X(_00966_));
 sky130_fd_sc_hd__xor2_1 _07876_ (.A(_00960_),
    .B(_00962_),
    .X(_00967_));
 sky130_fd_sc_hd__o21ai_2 _07877_ (.A1(_00965_),
    .A2(_00966_),
    .B1(_00963_),
    .Y(_00968_));
 sky130_fd_sc_hd__xor2_1 _07878_ (.A(_00947_),
    .B(_00957_),
    .X(_00969_));
 sky130_fd_sc_hd__a21boi_2 _07879_ (.A1(_00968_),
    .A2(_00969_),
    .B1_N(_00958_),
    .Y(_00970_));
 sky130_fd_sc_hd__o21ba_1 _07880_ (.A1(_00941_),
    .A2(_00945_),
    .B1_N(_00970_),
    .X(_00971_));
 sky130_fd_sc_hd__xor2_1 _07881_ (.A(_00881_),
    .B(_00883_),
    .X(_00972_));
 sky130_fd_sc_hd__o22a_1 _07882_ (.A1(net122),
    .A2(net99),
    .B1(net136),
    .B2(net126),
    .X(_00973_));
 sky130_fd_sc_hd__xnor2_1 _07883_ (.A(net154),
    .B(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__a21o_2 _07884_ (.A1(_00161_),
    .A2(_00162_),
    .B1(net146),
    .X(_00975_));
 sky130_fd_sc_hd__or2_1 _07885_ (.A(net95),
    .B(net141),
    .X(_00976_));
 sky130_fd_sc_hd__nand3_1 _07886_ (.A(net101),
    .B(_00975_),
    .C(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__a21o_1 _07887_ (.A1(_00975_),
    .A2(_00976_),
    .B1(net101),
    .X(_00978_));
 sky130_fd_sc_hd__a21oi_1 _07888_ (.A1(_00977_),
    .A2(_00978_),
    .B1(_00974_),
    .Y(_00979_));
 sky130_fd_sc_hd__and3_1 _07889_ (.A(_00974_),
    .B(_00977_),
    .C(_00978_),
    .X(_00980_));
 sky130_fd_sc_hd__nor2_1 _07890_ (.A(_00979_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__o22a_1 _07891_ (.A1(net75),
    .A2(net139),
    .B1(net138),
    .B2(net116),
    .X(_00982_));
 sky130_fd_sc_hd__xnor2_1 _07892_ (.A(net150),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__o21bai_1 _07893_ (.A1(_00980_),
    .A2(_00983_),
    .B1_N(_00979_),
    .Y(_00984_));
 sky130_fd_sc_hd__and2_1 _07894_ (.A(_00972_),
    .B(_00984_),
    .X(_00985_));
 sky130_fd_sc_hd__a21o_1 _07895_ (.A1(_00188_),
    .A2(_00189_),
    .B1(net143),
    .X(_00986_));
 sky130_fd_sc_hd__or2_1 _07896_ (.A(net147),
    .B(net65),
    .X(_00987_));
 sky130_fd_sc_hd__nand3_1 _07897_ (.A(net92),
    .B(_00986_),
    .C(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__a21o_1 _07898_ (.A1(_00986_),
    .A2(_00987_),
    .B1(net92),
    .X(_00989_));
 sky130_fd_sc_hd__o32a_1 _07899_ (.A1(net181),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net67),
    .B2(net179),
    .X(_00990_));
 sky130_fd_sc_hd__xor2_1 _07900_ (.A(net104),
    .B(_00990_),
    .X(_00991_));
 sky130_fd_sc_hd__a21o_1 _07901_ (.A1(_00988_),
    .A2(_00989_),
    .B1(_00991_),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_1 _07902_ (.A(_00972_),
    .B(_00984_),
    .Y(_00993_));
 sky130_fd_sc_hd__or3_1 _07903_ (.A(_00985_),
    .B(_00992_),
    .C(_00993_),
    .X(_00994_));
 sky130_fd_sc_hd__nand2b_1 _07904_ (.A_N(_00985_),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__xnor2_2 _07905_ (.A(_00946_),
    .B(_00970_),
    .Y(_00996_));
 sky130_fd_sc_hd__a21o_1 _07906_ (.A1(_00995_),
    .A2(_00996_),
    .B1(_00971_),
    .X(_00997_));
 sky130_fd_sc_hd__nand2b_1 _07907_ (.A_N(_00938_),
    .B(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__xnor2_1 _07908_ (.A(_00938_),
    .B(_00997_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2b_1 _07909_ (.A_N(_00932_),
    .B(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__xnor2_1 _07910_ (.A(_00932_),
    .B(_00999_),
    .Y(_01001_));
 sky130_fd_sc_hd__nand3_1 _07911_ (.A(_00988_),
    .B(_00989_),
    .C(_00991_),
    .Y(_01002_));
 sky130_fd_sc_hd__xnor2_1 _07912_ (.A(_00953_),
    .B(_00955_),
    .Y(_01003_));
 sky130_fd_sc_hd__and3_1 _07913_ (.A(_00992_),
    .B(_01002_),
    .C(_01003_),
    .X(_01004_));
 sky130_fd_sc_hd__a21oi_1 _07914_ (.A1(_00992_),
    .A2(_01002_),
    .B1(_01003_),
    .Y(_01005_));
 sky130_fd_sc_hd__xor2_1 _07915_ (.A(_00981_),
    .B(_00983_),
    .X(_01006_));
 sky130_fd_sc_hd__or3_1 _07916_ (.A(_01004_),
    .B(_01005_),
    .C(_01006_),
    .X(_01007_));
 sky130_fd_sc_hd__o21ba_1 _07917_ (.A1(_01005_),
    .A2(_01006_),
    .B1_N(_01004_),
    .X(_01008_));
 sky130_fd_sc_hd__o22a_1 _07918_ (.A1(net114),
    .A2(net131),
    .B1(net169),
    .B2(net124),
    .X(_01009_));
 sky130_fd_sc_hd__xnor2_2 _07919_ (.A(net193),
    .B(_01009_),
    .Y(_01010_));
 sky130_fd_sc_hd__o22a_1 _07920_ (.A1(net99),
    .A2(net87),
    .B1(net82),
    .B2(net97),
    .X(_01011_));
 sky130_fd_sc_hd__xnor2_2 _07921_ (.A(net187),
    .B(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__nor2_1 _07922_ (.A(_01010_),
    .B(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__xor2_2 _07923_ (.A(_01010_),
    .B(_01012_),
    .X(_01014_));
 sky130_fd_sc_hd__o22a_1 _07924_ (.A1(net90),
    .A2(net129),
    .B1(net127),
    .B2(net118),
    .X(_01015_));
 sky130_fd_sc_hd__xnor2_1 _07925_ (.A(net166),
    .B(_01015_),
    .Y(_01016_));
 sky130_fd_sc_hd__inv_2 _07926_ (.A(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__a21oi_2 _07927_ (.A1(_01014_),
    .A2(_01017_),
    .B1(_01013_),
    .Y(_01018_));
 sky130_fd_sc_hd__o22a_1 _07928_ (.A1(net225),
    .A2(net26),
    .B1(net73),
    .B2(net184),
    .X(_01019_));
 sky130_fd_sc_hd__xnor2_2 _07929_ (.A(net106),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__and2b_1 _07930_ (.A_N(_01018_),
    .B(_01020_),
    .X(_01021_));
 sky130_fd_sc_hd__o22a_2 _07931_ (.A1(net305),
    .A2(net47),
    .B1(net38),
    .B2(net256),
    .X(_01022_));
 sky130_fd_sc_hd__xnor2_4 _07932_ (.A(net258),
    .B(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__o22a_2 _07933_ (.A1(net120),
    .A2(net133),
    .B1(net171),
    .B2(net84),
    .X(_01024_));
 sky130_fd_sc_hd__xnor2_4 _07934_ (.A(net210),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__nor2_1 _07935_ (.A(_01023_),
    .B(_01025_),
    .Y(_01026_));
 sky130_fd_sc_hd__o22a_2 _07936_ (.A1(net176),
    .A2(net79),
    .B1(net41),
    .B2(net173),
    .X(_01027_));
 sky130_fd_sc_hd__xnor2_4 _07937_ (.A(net214),
    .B(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__xor2_4 _07938_ (.A(_01023_),
    .B(_01025_),
    .X(_01029_));
 sky130_fd_sc_hd__a21o_1 _07939_ (.A1(_01028_),
    .A2(_01029_),
    .B1(_01026_),
    .X(_01030_));
 sky130_fd_sc_hd__xnor2_2 _07940_ (.A(_01018_),
    .B(_01020_),
    .Y(_01031_));
 sky130_fd_sc_hd__a21oi_2 _07941_ (.A1(_01030_),
    .A2(_01031_),
    .B1(_01021_),
    .Y(_01032_));
 sky130_fd_sc_hd__nor2_1 _07942_ (.A(_01008_),
    .B(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__xnor2_2 _07943_ (.A(_00965_),
    .B(_00967_),
    .Y(_01034_));
 sky130_fd_sc_hd__o22a_1 _07944_ (.A1(net126),
    .A2(net138),
    .B1(net136),
    .B2(net122),
    .X(_01035_));
 sky130_fd_sc_hd__xnor2_1 _07945_ (.A(net154),
    .B(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__o22a_1 _07946_ (.A1(net147),
    .A2(net69),
    .B1(net95),
    .B2(net145),
    .X(_01037_));
 sky130_fd_sc_hd__xnor2_1 _07947_ (.A(_00153_),
    .B(_01037_),
    .Y(_01038_));
 sky130_fd_sc_hd__nor2_1 _07948_ (.A(_01036_),
    .B(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__xnor2_1 _07949_ (.A(_01036_),
    .B(_01038_),
    .Y(_01040_));
 sky130_fd_sc_hd__o22a_1 _07950_ (.A1(net75),
    .A2(net141),
    .B1(net139),
    .B2(net116),
    .X(_01041_));
 sky130_fd_sc_hd__xnor2_1 _07951_ (.A(net150),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__o21ba_1 _07952_ (.A1(_01040_),
    .A2(_01042_),
    .B1_N(_01039_),
    .X(_01043_));
 sky130_fd_sc_hd__and2b_1 _07953_ (.A_N(_01043_),
    .B(_01034_),
    .X(_01044_));
 sky130_fd_sc_hd__a21o_1 _07954_ (.A1(_00188_),
    .A2(_00189_),
    .B1(net179),
    .X(_01045_));
 sky130_fd_sc_hd__or2_1 _07955_ (.A(net143),
    .B(net65),
    .X(_01046_));
 sky130_fd_sc_hd__nand3_1 _07956_ (.A(net92),
    .B(_01045_),
    .C(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__a21o_1 _07957_ (.A1(_01045_),
    .A2(_01046_),
    .B1(net92),
    .X(_01048_));
 sky130_fd_sc_hd__o32a_1 _07958_ (.A1(net184),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net67),
    .B2(net181),
    .X(_01049_));
 sky130_fd_sc_hd__xor2_1 _07959_ (.A(net104),
    .B(_01049_),
    .X(_01050_));
 sky130_fd_sc_hd__a21o_1 _07960_ (.A1(_01047_),
    .A2(_01048_),
    .B1(_01050_),
    .X(_01051_));
 sky130_fd_sc_hd__inv_2 _07961_ (.A(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__xnor2_2 _07962_ (.A(_01034_),
    .B(_01043_),
    .Y(_01053_));
 sky130_fd_sc_hd__a21o_1 _07963_ (.A1(_01052_),
    .A2(_01053_),
    .B1(_01044_),
    .X(_01054_));
 sky130_fd_sc_hd__xor2_2 _07964_ (.A(_01008_),
    .B(_01032_),
    .X(_01055_));
 sky130_fd_sc_hd__a21oi_2 _07965_ (.A1(_01054_),
    .A2(_01055_),
    .B1(_01033_),
    .Y(_01056_));
 sky130_fd_sc_hd__xnor2_2 _07966_ (.A(_00995_),
    .B(_00996_),
    .Y(_01057_));
 sky130_fd_sc_hd__a21oi_1 _07967_ (.A1(_00942_),
    .A2(_00943_),
    .B1(_00944_),
    .Y(_01058_));
 sky130_fd_sc_hd__xnor2_1 _07968_ (.A(_00968_),
    .B(_00969_),
    .Y(_01059_));
 sky130_fd_sc_hd__or3_1 _07969_ (.A(_00945_),
    .B(_01058_),
    .C(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__o21ai_1 _07970_ (.A1(_00945_),
    .A2(_01058_),
    .B1(_01059_),
    .Y(_01061_));
 sky130_fd_sc_hd__o21ai_1 _07971_ (.A1(_00985_),
    .A2(_00993_),
    .B1(_00992_),
    .Y(_01062_));
 sky130_fd_sc_hd__and2_1 _07972_ (.A(_00994_),
    .B(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__nand3_1 _07973_ (.A(_01060_),
    .B(_01061_),
    .C(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(_01060_),
    .B(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__xnor2_2 _07975_ (.A(_01056_),
    .B(_01057_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2b_1 _07976_ (.A_N(_01066_),
    .B(_01065_),
    .Y(_01067_));
 sky130_fd_sc_hd__o21ai_2 _07977_ (.A1(_01056_),
    .A2(_01057_),
    .B1(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__xnor2_1 _07978_ (.A(_00875_),
    .B(_01001_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2b_1 _07979_ (.A_N(_01069_),
    .B(_01068_),
    .Y(_01070_));
 sky130_fd_sc_hd__a21bo_2 _07980_ (.A1(_00875_),
    .A2(_01001_),
    .B1_N(_01070_),
    .X(_01071_));
 sky130_fd_sc_hd__nand2_2 _07981_ (.A(_00998_),
    .B(_01000_),
    .Y(_01072_));
 sky130_fd_sc_hd__o21a_1 _07982_ (.A1(_00793_),
    .A2(_00796_),
    .B1(_00795_),
    .X(_01073_));
 sky130_fd_sc_hd__nand2_1 _07983_ (.A(_00711_),
    .B(_00712_),
    .Y(_01074_));
 sky130_fd_sc_hd__and2_1 _07984_ (.A(_00713_),
    .B(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__o21ai_1 _07985_ (.A1(_00781_),
    .A2(_00785_),
    .B1(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__or3_1 _07986_ (.A(_00781_),
    .B(_00785_),
    .C(_01075_),
    .X(_01077_));
 sky130_fd_sc_hd__and2_1 _07987_ (.A(_01076_),
    .B(_01077_),
    .X(_01078_));
 sky130_fd_sc_hd__nand2b_1 _07988_ (.A_N(_01073_),
    .B(_01078_),
    .Y(_01079_));
 sky130_fd_sc_hd__xnor2_2 _07989_ (.A(_01073_),
    .B(_01078_),
    .Y(_01080_));
 sky130_fd_sc_hd__nor2_1 _07990_ (.A(_00733_),
    .B(_00735_),
    .Y(_01081_));
 sky130_fd_sc_hd__or2_1 _07991_ (.A(_00736_),
    .B(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__or2_1 _07992_ (.A(_00701_),
    .B(_00703_),
    .X(_01083_));
 sky130_fd_sc_hd__and2_1 _07993_ (.A(_00704_),
    .B(_01083_),
    .X(_01084_));
 sky130_fd_sc_hd__inv_2 _07994_ (.A(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__xnor2_1 _07995_ (.A(_00754_),
    .B(_00755_),
    .Y(_01086_));
 sky130_fd_sc_hd__xnor2_1 _07996_ (.A(_01085_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__xnor2_1 _07997_ (.A(_01082_),
    .B(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__o21ai_1 _07998_ (.A1(_00853_),
    .A2(_00860_),
    .B1(_00858_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(_00387_),
    .B(_00389_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _08000_ (.A(_00390_),
    .B(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__a21o_1 _08001_ (.A1(_00804_),
    .A2(_00806_),
    .B1(_00802_),
    .X(_01092_));
 sky130_fd_sc_hd__xor2_1 _08002_ (.A(_01091_),
    .B(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__and2b_1 _08003_ (.A_N(_01093_),
    .B(_01089_),
    .X(_01094_));
 sky130_fd_sc_hd__xor2_1 _08004_ (.A(_01089_),
    .B(_01093_),
    .X(_01095_));
 sky130_fd_sc_hd__nor2_1 _08005_ (.A(_01088_),
    .B(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__and2_1 _08006_ (.A(_01088_),
    .B(_01095_),
    .X(_01097_));
 sky130_fd_sc_hd__nor2_1 _08007_ (.A(_01096_),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__xor2_2 _08008_ (.A(_01080_),
    .B(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__o21ai_2 _08009_ (.A1(_00837_),
    .A2(_00874_),
    .B1(_00836_),
    .Y(_01100_));
 sky130_fd_sc_hd__a21bo_1 _08010_ (.A1(_00933_),
    .A2(_00937_),
    .B1_N(_00936_),
    .X(_01101_));
 sky130_fd_sc_hd__a21o_2 _08011_ (.A1(_00851_),
    .A2(_00873_),
    .B1(_00871_),
    .X(_01102_));
 sky130_fd_sc_hd__a21o_2 _08012_ (.A1(_00788_),
    .A2(_00809_),
    .B1(_00808_),
    .X(_01103_));
 sky130_fd_sc_hd__nor2_2 _08013_ (.A(_00831_),
    .B(_00834_),
    .Y(_01104_));
 sky130_fd_sc_hd__o21a_1 _08014_ (.A1(_00831_),
    .A2(_00834_),
    .B1(_01103_),
    .X(_01105_));
 sky130_fd_sc_hd__xnor2_4 _08015_ (.A(_01103_),
    .B(_01104_),
    .Y(_01106_));
 sky130_fd_sc_hd__xor2_2 _08016_ (.A(_01102_),
    .B(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__xnor2_2 _08017_ (.A(_01101_),
    .B(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand2b_1 _08018_ (.A_N(_01108_),
    .B(_01100_),
    .Y(_01109_));
 sky130_fd_sc_hd__xnor2_2 _08019_ (.A(_01100_),
    .B(_01108_),
    .Y(_01110_));
 sky130_fd_sc_hd__and2_1 _08020_ (.A(_01099_),
    .B(_01110_),
    .X(_01111_));
 sky130_fd_sc_hd__xor2_2 _08021_ (.A(_01099_),
    .B(_01110_),
    .X(_01112_));
 sky130_fd_sc_hd__xor2_2 _08022_ (.A(_01072_),
    .B(_01112_),
    .X(_01113_));
 sky130_fd_sc_hd__or2_1 _08023_ (.A(_01071_),
    .B(_01113_),
    .X(_01114_));
 sky130_fd_sc_hd__xor2_1 _08024_ (.A(_01068_),
    .B(_01069_),
    .X(_01115_));
 sky130_fd_sc_hd__a21oi_1 _08025_ (.A1(_00909_),
    .A2(_00930_),
    .B1(_00929_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_1 _08026_ (.A(_00931_),
    .B(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__xnor2_2 _08027_ (.A(_01065_),
    .B(_01066_),
    .Y(_01118_));
 sky130_fd_sc_hd__xnor2_1 _08028_ (.A(_01054_),
    .B(_01055_),
    .Y(_01119_));
 sky130_fd_sc_hd__xnor2_1 _08029_ (.A(_01014_),
    .B(_01016_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand3_1 _08030_ (.A(_01047_),
    .B(_01048_),
    .C(_01050_),
    .Y(_01121_));
 sky130_fd_sc_hd__and3_1 _08031_ (.A(_01051_),
    .B(_01120_),
    .C(_01121_),
    .X(_01122_));
 sky130_fd_sc_hd__a21oi_1 _08032_ (.A1(_01051_),
    .A2(_01121_),
    .B1(_01120_),
    .Y(_01123_));
 sky130_fd_sc_hd__xnor2_1 _08033_ (.A(_01040_),
    .B(_01042_),
    .Y(_01124_));
 sky130_fd_sc_hd__or3_1 _08034_ (.A(_01122_),
    .B(_01123_),
    .C(_01124_),
    .X(_01125_));
 sky130_fd_sc_hd__o21ba_1 _08035_ (.A1(_01123_),
    .A2(_01124_),
    .B1_N(_01122_),
    .X(_01126_));
 sky130_fd_sc_hd__o22a_1 _08036_ (.A1(net124),
    .A2(net133),
    .B1(net171),
    .B2(net120),
    .X(_01127_));
 sky130_fd_sc_hd__xnor2_1 _08037_ (.A(net210),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__or3_1 _08038_ (.A(net256),
    .B(_00310_),
    .C(_00311_),
    .X(_01129_));
 sky130_fd_sc_hd__a21o_2 _08039_ (.A1(_00315_),
    .A2(_00316_),
    .B1(net306),
    .X(_01130_));
 sky130_fd_sc_hd__a21oi_1 _08040_ (.A1(_01129_),
    .A2(_01130_),
    .B1(net258),
    .Y(_01131_));
 sky130_fd_sc_hd__and3_1 _08041_ (.A(net258),
    .B(_01129_),
    .C(_01130_),
    .X(_01132_));
 sky130_fd_sc_hd__or3_2 _08042_ (.A(_01128_),
    .B(_01131_),
    .C(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__o22a_1 _08043_ (.A1(net176),
    .A2(net84),
    .B1(net79),
    .B2(net173),
    .X(_01134_));
 sky130_fd_sc_hd__xnor2_1 _08044_ (.A(net214),
    .B(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__o21ai_1 _08045_ (.A1(_01131_),
    .A2(_01132_),
    .B1(_01128_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand3_2 _08046_ (.A(_01133_),
    .B(_01135_),
    .C(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__a211o_1 _08047_ (.A1(_01133_),
    .A2(_01137_),
    .B1(net225),
    .C1(net73),
    .X(_01138_));
 sky130_fd_sc_hd__o21ai_1 _08048_ (.A1(net225),
    .A2(net73),
    .B1(net106),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_01138_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2b_1 _08050_ (.A_N(_01126_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__o22a_1 _08051_ (.A1(net118),
    .A2(net131),
    .B1(net169),
    .B2(net114),
    .X(_01142_));
 sky130_fd_sc_hd__xnor2_1 _08052_ (.A(net193),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__o22a_1 _08053_ (.A1(net136),
    .A2(net87),
    .B1(net82),
    .B2(net99),
    .X(_01144_));
 sky130_fd_sc_hd__xnor2_1 _08054_ (.A(net187),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__xor2_1 _08055_ (.A(_01143_),
    .B(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__o22a_1 _08056_ (.A1(net97),
    .A2(net129),
    .B1(net127),
    .B2(net90),
    .X(_01147_));
 sky130_fd_sc_hd__xnor2_1 _08057_ (.A(net166),
    .B(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__and2b_1 _08058_ (.A_N(_01148_),
    .B(_01146_),
    .X(_01149_));
 sky130_fd_sc_hd__o21ba_2 _08059_ (.A1(_01143_),
    .A2(_01145_),
    .B1_N(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__xor2_4 _08060_ (.A(_01028_),
    .B(_01029_),
    .X(_01151_));
 sky130_fd_sc_hd__and2b_1 _08061_ (.A_N(_01150_),
    .B(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__o22a_1 _08062_ (.A1(net126),
    .A2(net139),
    .B1(net138),
    .B2(net122),
    .X(_01153_));
 sky130_fd_sc_hd__xnor2_2 _08063_ (.A(net154),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__o22a_1 _08064_ (.A1(net75),
    .A2(net145),
    .B1(net141),
    .B2(net116),
    .X(_01155_));
 sky130_fd_sc_hd__xnor2_1 _08065_ (.A(net150),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__nor2_2 _08066_ (.A(_01154_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__xnor2_4 _08067_ (.A(_01150_),
    .B(_01151_),
    .Y(_01158_));
 sky130_fd_sc_hd__a21o_1 _08068_ (.A1(_01157_),
    .A2(_01158_),
    .B1(_01152_),
    .X(_01159_));
 sky130_fd_sc_hd__xnor2_2 _08069_ (.A(_01126_),
    .B(_01140_),
    .Y(_01160_));
 sky130_fd_sc_hd__a21boi_1 _08070_ (.A1(_01159_),
    .A2(_01160_),
    .B1_N(_01141_),
    .Y(_01161_));
 sky130_fd_sc_hd__o21ai_1 _08071_ (.A1(_01004_),
    .A2(_01005_),
    .B1(_01006_),
    .Y(_01162_));
 sky130_fd_sc_hd__xor2_1 _08072_ (.A(_01030_),
    .B(_01031_),
    .X(_01163_));
 sky130_fd_sc_hd__and3_1 _08073_ (.A(_01007_),
    .B(_01162_),
    .C(_01163_),
    .X(_01164_));
 sky130_fd_sc_hd__a21oi_1 _08074_ (.A1(_01007_),
    .A2(_01162_),
    .B1(_01163_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _08075_ (.A(_01164_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__xnor2_2 _08076_ (.A(_01052_),
    .B(_01053_),
    .Y(_01167_));
 sky130_fd_sc_hd__o21ba_1 _08077_ (.A1(_01165_),
    .A2(_01167_),
    .B1_N(_01164_),
    .X(_01168_));
 sky130_fd_sc_hd__xor2_1 _08078_ (.A(_01119_),
    .B(_01161_),
    .X(_01169_));
 sky130_fd_sc_hd__nand2b_1 _08079_ (.A_N(_01168_),
    .B(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__o21ai_1 _08080_ (.A1(_01119_),
    .A2(_01161_),
    .B1(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__xnor2_1 _08081_ (.A(_01117_),
    .B(_01118_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2b_1 _08082_ (.A_N(_01172_),
    .B(_01171_),
    .Y(_01173_));
 sky130_fd_sc_hd__a21boi_2 _08083_ (.A1(_01117_),
    .A2(_01118_),
    .B1_N(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__or2_1 _08084_ (.A(_01115_),
    .B(_01174_),
    .X(_01175_));
 sky130_fd_sc_hd__a21bo_1 _08085_ (.A1(_01071_),
    .A2(_01113_),
    .B1_N(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__o22a_1 _08086_ (.A1(net99),
    .A2(net131),
    .B1(net169),
    .B2(net97),
    .X(_01177_));
 sky130_fd_sc_hd__xnor2_1 _08087_ (.A(net193),
    .B(_01177_),
    .Y(_01178_));
 sky130_fd_sc_hd__o22a_1 _08088_ (.A1(net138),
    .A2(net129),
    .B1(net127),
    .B2(net136),
    .X(_01179_));
 sky130_fd_sc_hd__xnor2_1 _08089_ (.A(net166),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__or2_2 _08090_ (.A(_01178_),
    .B(_01180_),
    .X(_01181_));
 sky130_fd_sc_hd__o22a_1 _08091_ (.A1(net97),
    .A2(net131),
    .B1(net169),
    .B2(net90),
    .X(_01182_));
 sky130_fd_sc_hd__xnor2_2 _08092_ (.A(net193),
    .B(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__o22a_1 _08093_ (.A1(net136),
    .A2(net129),
    .B1(net127),
    .B2(net99),
    .X(_01184_));
 sky130_fd_sc_hd__xnor2_2 _08094_ (.A(net166),
    .B(_01184_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _08095_ (.A(_01183_),
    .B(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__xnor2_2 _08096_ (.A(_01183_),
    .B(_01185_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _08097_ (.A(_01181_),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__xor2_2 _08098_ (.A(_01181_),
    .B(_01187_),
    .X(_01189_));
 sky130_fd_sc_hd__o22a_1 _08099_ (.A1(net124),
    .A2(net176),
    .B1(net173),
    .B2(net120),
    .X(_01190_));
 sky130_fd_sc_hd__xnor2_2 _08100_ (.A(net212),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__o22a_1 _08101_ (.A1(net118),
    .A2(net133),
    .B1(net171),
    .B2(net114),
    .X(_01192_));
 sky130_fd_sc_hd__xnor2_2 _08102_ (.A(net210),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__o22a_1 _08103_ (.A1(net256),
    .A2(net84),
    .B1(net79),
    .B2(net305),
    .X(_01194_));
 sky130_fd_sc_hd__xnor2_2 _08104_ (.A(net258),
    .B(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__or2_1 _08105_ (.A(_01193_),
    .B(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__xor2_2 _08106_ (.A(_01193_),
    .B(_01195_),
    .X(_01197_));
 sky130_fd_sc_hd__nand2b_1 _08107_ (.A_N(_01191_),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__xnor2_2 _08108_ (.A(_01191_),
    .B(_01197_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _08109_ (.A(_01189_),
    .B(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__or2_1 _08110_ (.A(_01189_),
    .B(_01199_),
    .X(_01201_));
 sky130_fd_sc_hd__nand2_1 _08111_ (.A(_01200_),
    .B(_01201_),
    .Y(_01202_));
 sky130_fd_sc_hd__o22a_1 _08112_ (.A1(net126),
    .A2(net145),
    .B1(net141),
    .B2(net122),
    .X(_01203_));
 sky130_fd_sc_hd__xnor2_1 _08113_ (.A(net154),
    .B(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__o22a_1 _08114_ (.A1(net139),
    .A2(net87),
    .B1(net82),
    .B2(net138),
    .X(_01205_));
 sky130_fd_sc_hd__xnor2_1 _08115_ (.A(net187),
    .B(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__o22a_1 _08116_ (.A1(net116),
    .A2(net147),
    .B1(net143),
    .B2(net75),
    .X(_01207_));
 sky130_fd_sc_hd__xnor2_1 _08117_ (.A(net150),
    .B(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__or2_1 _08118_ (.A(_01206_),
    .B(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__xnor2_1 _08119_ (.A(_01206_),
    .B(_01208_),
    .Y(_01210_));
 sky130_fd_sc_hd__xor2_1 _08120_ (.A(_01204_),
    .B(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__xnor2_1 _08121_ (.A(_01202_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__o22a_1 _08122_ (.A1(net118),
    .A2(net171),
    .B1(net90),
    .B2(net133),
    .X(_01213_));
 sky130_fd_sc_hd__xnor2_2 _08123_ (.A(net210),
    .B(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__o22a_1 _08124_ (.A1(net120),
    .A2(net256),
    .B1(net84),
    .B2(net305),
    .X(_01215_));
 sky130_fd_sc_hd__xnor2_2 _08125_ (.A(net258),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _08126_ (.A(_01214_),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__o22a_1 _08127_ (.A1(net114),
    .A2(net176),
    .B1(net173),
    .B2(net124),
    .X(_01218_));
 sky130_fd_sc_hd__xnor2_2 _08128_ (.A(net212),
    .B(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__inv_2 _08129_ (.A(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__xor2_2 _08130_ (.A(_01214_),
    .B(_01216_),
    .X(_01221_));
 sky130_fd_sc_hd__a21oi_1 _08131_ (.A1(_01220_),
    .A2(_01221_),
    .B1(_01217_),
    .Y(_01222_));
 sky130_fd_sc_hd__o22a_1 _08132_ (.A1(net181),
    .A2(net69),
    .B1(net95),
    .B2(net179),
    .X(_01223_));
 sky130_fd_sc_hd__xnor2_1 _08133_ (.A(net101),
    .B(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2b_1 _08134_ (.A_N(_01222_),
    .B(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__xnor2_1 _08135_ (.A(_01222_),
    .B(_01224_),
    .Y(_01226_));
 sky130_fd_sc_hd__o22a_1 _08136_ (.A1(net225),
    .A2(net21),
    .B1(net65),
    .B2(net184),
    .X(_01227_));
 sky130_fd_sc_hd__xnor2_2 _08137_ (.A(net92),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__xor2_1 _08138_ (.A(_01226_),
    .B(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__xnor2_1 _08139_ (.A(_01212_),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__xnor2_2 _08140_ (.A(_01219_),
    .B(_01221_),
    .Y(_01231_));
 sky130_fd_sc_hd__o22a_1 _08141_ (.A1(net305),
    .A2(net120),
    .B1(net256),
    .B2(net124),
    .X(_01232_));
 sky130_fd_sc_hd__xnor2_1 _08142_ (.A(net258),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__o22a_1 _08143_ (.A1(net118),
    .A2(net176),
    .B1(net173),
    .B2(net114),
    .X(_01234_));
 sky130_fd_sc_hd__xnor2_1 _08144_ (.A(net212),
    .B(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__or2_1 _08145_ (.A(_01233_),
    .B(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__xnor2_1 _08146_ (.A(_01178_),
    .B(_01180_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _08147_ (.A(_01236_),
    .B(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(_01236_),
    .B(_01237_),
    .Y(_01239_));
 sky130_fd_sc_hd__and2b_1 _08149_ (.A_N(_01238_),
    .B(_01239_),
    .X(_01240_));
 sky130_fd_sc_hd__xnor2_2 _08150_ (.A(_01231_),
    .B(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__o22a_1 _08151_ (.A1(net126),
    .A2(net147),
    .B1(net145),
    .B2(net122),
    .X(_01242_));
 sky130_fd_sc_hd__xnor2_2 _08152_ (.A(net154),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__o22a_1 _08153_ (.A1(net141),
    .A2(net87),
    .B1(net82),
    .B2(net139),
    .X(_01244_));
 sky130_fd_sc_hd__xnor2_2 _08154_ (.A(net187),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__o22a_1 _08155_ (.A1(net75),
    .A2(net179),
    .B1(net143),
    .B2(net116),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_2 _08156_ (.A(net150),
    .B(_01246_),
    .Y(_01247_));
 sky130_fd_sc_hd__or2_1 _08157_ (.A(_01245_),
    .B(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__xnor2_2 _08158_ (.A(_01245_),
    .B(_01247_),
    .Y(_01249_));
 sky130_fd_sc_hd__xor2_2 _08159_ (.A(_01243_),
    .B(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__nand2b_1 _08160_ (.A_N(_01241_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__xnor2_2 _08161_ (.A(_01241_),
    .B(_01250_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _08162_ (.A(net225),
    .B(net65),
    .Y(_01253_));
 sky130_fd_sc_hd__o22a_1 _08163_ (.A1(net184),
    .A2(net69),
    .B1(net95),
    .B2(net181),
    .X(_01254_));
 sky130_fd_sc_hd__xnor2_1 _08164_ (.A(net101),
    .B(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__or3_1 _08165_ (.A(net225),
    .B(net65),
    .C(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__nand2b_1 _08166_ (.A_N(_01253_),
    .B(_01255_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_2 _08167_ (.A(_01256_),
    .B(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__a21bo_1 _08168_ (.A1(_01252_),
    .A2(_01258_),
    .B1_N(_01251_),
    .X(_01259_));
 sky130_fd_sc_hd__xor2_1 _08169_ (.A(_01233_),
    .B(_01235_),
    .X(_01260_));
 sky130_fd_sc_hd__o22a_1 _08170_ (.A1(net225),
    .A2(net69),
    .B1(net95),
    .B2(net184),
    .X(_01261_));
 sky130_fd_sc_hd__xnor2_1 _08171_ (.A(net101),
    .B(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__and2_1 _08172_ (.A(_01260_),
    .B(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__o22a_1 _08173_ (.A1(net118),
    .A2(net173),
    .B1(net90),
    .B2(net176),
    .X(_01264_));
 sky130_fd_sc_hd__xnor2_1 _08174_ (.A(net212),
    .B(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__o22a_1 _08175_ (.A1(net305),
    .A2(net124),
    .B1(net114),
    .B2(net256),
    .X(_01266_));
 sky130_fd_sc_hd__xnor2_1 _08176_ (.A(net258),
    .B(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__nor2_1 _08177_ (.A(_01265_),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__xor2_1 _08178_ (.A(_01260_),
    .B(_01262_),
    .X(_01269_));
 sky130_fd_sc_hd__a21o_1 _08179_ (.A1(_01268_),
    .A2(_01269_),
    .B1(_01263_),
    .X(_01270_));
 sky130_fd_sc_hd__o22a_1 _08180_ (.A1(net97),
    .A2(net133),
    .B1(net171),
    .B2(net90),
    .X(_01271_));
 sky130_fd_sc_hd__xnor2_1 _08181_ (.A(net210),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__o22a_1 _08182_ (.A1(net139),
    .A2(net129),
    .B1(net127),
    .B2(net138),
    .X(_01273_));
 sky130_fd_sc_hd__xnor2_1 _08183_ (.A(net166),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__or2_1 _08184_ (.A(_01272_),
    .B(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__o22a_1 _08185_ (.A1(net136),
    .A2(net131),
    .B1(net169),
    .B2(net99),
    .X(_01276_));
 sky130_fd_sc_hd__xnor2_1 _08186_ (.A(net193),
    .B(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__xnor2_1 _08187_ (.A(_01272_),
    .B(_01274_),
    .Y(_01278_));
 sky130_fd_sc_hd__or2_1 _08188_ (.A(_01277_),
    .B(_01278_),
    .X(_01279_));
 sky130_fd_sc_hd__and2_1 _08189_ (.A(_01275_),
    .B(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__a21boi_1 _08190_ (.A1(_01275_),
    .A2(_01279_),
    .B1_N(_01270_),
    .Y(_01281_));
 sky130_fd_sc_hd__o22a_1 _08191_ (.A1(net145),
    .A2(net87),
    .B1(net82),
    .B2(net141),
    .X(_01282_));
 sky130_fd_sc_hd__xnor2_2 _08192_ (.A(net187),
    .B(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__o22a_1 _08193_ (.A1(net75),
    .A2(net181),
    .B1(net179),
    .B2(net116),
    .X(_01284_));
 sky130_fd_sc_hd__xnor2_1 _08194_ (.A(net150),
    .B(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__o22a_1 _08195_ (.A1(net122),
    .A2(net147),
    .B1(net143),
    .B2(net126),
    .X(_01286_));
 sky130_fd_sc_hd__xnor2_1 _08196_ (.A(net154),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__xnor2_1 _08197_ (.A(_01283_),
    .B(_01285_),
    .Y(_01288_));
 sky130_fd_sc_hd__or2_1 _08198_ (.A(_01287_),
    .B(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__o21ai_2 _08199_ (.A1(_01283_),
    .A2(_01285_),
    .B1(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__xnor2_2 _08200_ (.A(_01270_),
    .B(_01280_),
    .Y(_01291_));
 sky130_fd_sc_hd__a21o_1 _08201_ (.A1(_01290_),
    .A2(_01291_),
    .B1(_01281_),
    .X(_01292_));
 sky130_fd_sc_hd__o21ai_2 _08202_ (.A1(net92),
    .A2(_01253_),
    .B1(_01256_),
    .Y(_01293_));
 sky130_fd_sc_hd__a21o_1 _08203_ (.A1(_01231_),
    .A2(_01239_),
    .B1(_01238_),
    .X(_01294_));
 sky130_fd_sc_hd__o21ai_2 _08204_ (.A1(_01243_),
    .A2(_01249_),
    .B1(_01248_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _08205_ (.A(_01294_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__nor2_1 _08206_ (.A(_01294_),
    .B(_01295_),
    .Y(_01297_));
 sky130_fd_sc_hd__xor2_1 _08207_ (.A(_01294_),
    .B(_01295_),
    .X(_01298_));
 sky130_fd_sc_hd__xnor2_1 _08208_ (.A(_01293_),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__and2_1 _08209_ (.A(_01292_),
    .B(_01299_),
    .X(_01300_));
 sky130_fd_sc_hd__xor2_1 _08210_ (.A(_01292_),
    .B(_01299_),
    .X(_01301_));
 sky130_fd_sc_hd__xnor2_1 _08211_ (.A(_01259_),
    .B(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__nor2_1 _08212_ (.A(_01230_),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__xor2_1 _08213_ (.A(_01230_),
    .B(_01302_),
    .X(_01304_));
 sky130_fd_sc_hd__xnor2_2 _08214_ (.A(_01290_),
    .B(_01291_),
    .Y(_01305_));
 sky130_fd_sc_hd__xor2_1 _08215_ (.A(_01265_),
    .B(_01267_),
    .X(_01306_));
 sky130_fd_sc_hd__nor2_1 _08216_ (.A(net225),
    .B(net95),
    .Y(_01307_));
 sky130_fd_sc_hd__mux2_1 _08217_ (.A0(net101),
    .A1(_01306_),
    .S(_01307_),
    .X(_01308_));
 sky130_fd_sc_hd__o22a_1 _08218_ (.A1(net99),
    .A2(net133),
    .B1(net171),
    .B2(net97),
    .X(_01309_));
 sky130_fd_sc_hd__xnor2_2 _08219_ (.A(net210),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__o22a_1 _08220_ (.A1(net141),
    .A2(net129),
    .B1(net127),
    .B2(net139),
    .X(_01311_));
 sky130_fd_sc_hd__xnor2_2 _08221_ (.A(net166),
    .B(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__or2_1 _08222_ (.A(_01310_),
    .B(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__o22a_1 _08223_ (.A1(net138),
    .A2(net131),
    .B1(net169),
    .B2(net136),
    .X(_01314_));
 sky130_fd_sc_hd__xnor2_2 _08224_ (.A(net193),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__xnor2_2 _08225_ (.A(_01310_),
    .B(_01312_),
    .Y(_01316_));
 sky130_fd_sc_hd__o21ai_2 _08226_ (.A1(_01315_),
    .A2(_01316_),
    .B1(_01313_),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _08227_ (.A(_01308_),
    .B(_01317_),
    .Y(_01318_));
 sky130_fd_sc_hd__o22a_1 _08228_ (.A1(net147),
    .A2(net87),
    .B1(net82),
    .B2(net145),
    .X(_01319_));
 sky130_fd_sc_hd__xnor2_1 _08229_ (.A(net187),
    .B(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__o22a_1 _08230_ (.A1(net75),
    .A2(net184),
    .B1(net181),
    .B2(net116),
    .X(_01321_));
 sky130_fd_sc_hd__xnor2_1 _08231_ (.A(net150),
    .B(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__or2_1 _08232_ (.A(_01320_),
    .B(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__o22a_1 _08233_ (.A1(net126),
    .A2(net179),
    .B1(net143),
    .B2(net122),
    .X(_01324_));
 sky130_fd_sc_hd__xnor2_1 _08234_ (.A(net154),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__xnor2_1 _08235_ (.A(_01320_),
    .B(_01322_),
    .Y(_01326_));
 sky130_fd_sc_hd__o21a_1 _08236_ (.A1(_01325_),
    .A2(_01326_),
    .B1(_01323_),
    .X(_01327_));
 sky130_fd_sc_hd__nor2_1 _08237_ (.A(_01308_),
    .B(_01317_),
    .Y(_01328_));
 sky130_fd_sc_hd__xor2_1 _08238_ (.A(_01308_),
    .B(_01317_),
    .X(_01329_));
 sky130_fd_sc_hd__o21a_1 _08239_ (.A1(_01327_),
    .A2(_01328_),
    .B1(_01318_),
    .X(_01330_));
 sky130_fd_sc_hd__xnor2_1 _08240_ (.A(_01268_),
    .B(_01269_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _08241_ (.A(_01277_),
    .B(_01278_),
    .Y(_01332_));
 sky130_fd_sc_hd__and2_1 _08242_ (.A(_01279_),
    .B(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__nand2b_1 _08243_ (.A_N(_01331_),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__xnor2_1 _08244_ (.A(_01331_),
    .B(_01333_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(_01287_),
    .B(_01288_),
    .Y(_01336_));
 sky130_fd_sc_hd__and2_1 _08246_ (.A(_01289_),
    .B(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(_01335_),
    .B(_01337_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _08248_ (.A(_01334_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__xnor2_1 _08249_ (.A(_01305_),
    .B(_01330_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2b_1 _08250_ (.A_N(_01340_),
    .B(_01339_),
    .Y(_01341_));
 sky130_fd_sc_hd__o21ai_2 _08251_ (.A1(_01305_),
    .A2(_01330_),
    .B1(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__xor2_1 _08252_ (.A(_01304_),
    .B(_01342_),
    .X(_01343_));
 sky130_fd_sc_hd__xor2_2 _08253_ (.A(_01252_),
    .B(_01258_),
    .X(_01344_));
 sky130_fd_sc_hd__xnor2_1 _08254_ (.A(_01339_),
    .B(_01340_),
    .Y(_01345_));
 sky130_fd_sc_hd__and2_1 _08255_ (.A(_01344_),
    .B(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__o22a_1 _08256_ (.A1(net126),
    .A2(net181),
    .B1(net179),
    .B2(net122),
    .X(_01347_));
 sky130_fd_sc_hd__xnor2_2 _08257_ (.A(net154),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__o22a_1 _08258_ (.A1(net225),
    .A2(net75),
    .B1(net116),
    .B2(net184),
    .X(_01349_));
 sky130_fd_sc_hd__xnor2_2 _08259_ (.A(net150),
    .B(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_1 _08260_ (.A(_01348_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__o22a_1 _08261_ (.A1(net136),
    .A2(net133),
    .B1(net171),
    .B2(net99),
    .X(_01352_));
 sky130_fd_sc_hd__xnor2_2 _08262_ (.A(net210),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__o22a_1 _08263_ (.A1(net305),
    .A2(net114),
    .B1(net256),
    .B2(net118),
    .X(_01354_));
 sky130_fd_sc_hd__xnor2_2 _08264_ (.A(net258),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__or2_1 _08265_ (.A(_01353_),
    .B(_01355_),
    .X(_01356_));
 sky130_fd_sc_hd__xnor2_2 _08266_ (.A(_01353_),
    .B(_01355_),
    .Y(_01357_));
 sky130_fd_sc_hd__o22a_1 _08267_ (.A1(net97),
    .A2(net176),
    .B1(net173),
    .B2(net90),
    .X(_01358_));
 sky130_fd_sc_hd__xnor2_2 _08268_ (.A(net212),
    .B(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__o21a_1 _08269_ (.A1(_01357_),
    .A2(_01359_),
    .B1(_01356_),
    .X(_01360_));
 sky130_fd_sc_hd__or3_1 _08270_ (.A(_01348_),
    .B(_01350_),
    .C(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__o22a_1 _08271_ (.A1(net143),
    .A2(net87),
    .B1(net82),
    .B2(net147),
    .X(_01362_));
 sky130_fd_sc_hd__xnor2_2 _08272_ (.A(net187),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__o22a_1 _08273_ (.A1(net139),
    .A2(net131),
    .B1(net169),
    .B2(net138),
    .X(_01364_));
 sky130_fd_sc_hd__xnor2_2 _08274_ (.A(net193),
    .B(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__xor2_1 _08275_ (.A(_01363_),
    .B(_01365_),
    .X(_01366_));
 sky130_fd_sc_hd__o22a_1 _08276_ (.A1(net145),
    .A2(net129),
    .B1(net127),
    .B2(net141),
    .X(_01367_));
 sky130_fd_sc_hd__xnor2_1 _08277_ (.A(net166),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__nand2b_1 _08278_ (.A_N(_01368_),
    .B(_01366_),
    .Y(_01369_));
 sky130_fd_sc_hd__o21ai_2 _08279_ (.A1(_01363_),
    .A2(_01365_),
    .B1(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__xnor2_2 _08280_ (.A(_01351_),
    .B(_01360_),
    .Y(_01371_));
 sky130_fd_sc_hd__a21boi_1 _08281_ (.A1(_01370_),
    .A2(_01371_),
    .B1_N(_01361_),
    .Y(_01372_));
 sky130_fd_sc_hd__xnor2_1 _08282_ (.A(_01327_),
    .B(_01329_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2b_1 _08283_ (.A_N(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__xor2_1 _08284_ (.A(_01315_),
    .B(_01316_),
    .X(_01375_));
 sky130_fd_sc_hd__xnor2_1 _08285_ (.A(_01306_),
    .B(_01307_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2b_1 _08286_ (.A_N(_01376_),
    .B(_01375_),
    .Y(_01377_));
 sky130_fd_sc_hd__xor2_1 _08287_ (.A(_01325_),
    .B(_01326_),
    .X(_01378_));
 sky130_fd_sc_hd__xnor2_1 _08288_ (.A(_01375_),
    .B(_01376_),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _08289_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__and2_1 _08290_ (.A(_01377_),
    .B(_01380_),
    .X(_01381_));
 sky130_fd_sc_hd__xor2_1 _08291_ (.A(_01372_),
    .B(_01373_),
    .X(_01382_));
 sky130_fd_sc_hd__o21ai_1 _08292_ (.A1(_01381_),
    .A2(_01382_),
    .B1(_01374_),
    .Y(_01383_));
 sky130_fd_sc_hd__xnor2_1 _08293_ (.A(_01344_),
    .B(_01345_),
    .Y(_01384_));
 sky130_fd_sc_hd__and2b_1 _08294_ (.A_N(_01384_),
    .B(_01383_),
    .X(_01385_));
 sky130_fd_sc_hd__nor3_1 _08295_ (.A(_01343_),
    .B(_01346_),
    .C(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__or2_1 _08296_ (.A(_01335_),
    .B(_01337_),
    .X(_01387_));
 sky130_fd_sc_hd__nand2_1 _08297_ (.A(_01338_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__xnor2_1 _08298_ (.A(_01381_),
    .B(_01382_),
    .Y(_01389_));
 sky130_fd_sc_hd__or2_1 _08299_ (.A(_01388_),
    .B(_01389_),
    .X(_01390_));
 sky130_fd_sc_hd__xor2_1 _08300_ (.A(_01388_),
    .B(_01389_),
    .X(_01391_));
 sky130_fd_sc_hd__xnor2_2 _08301_ (.A(_01370_),
    .B(_01371_),
    .Y(_01392_));
 sky130_fd_sc_hd__o22a_1 _08302_ (.A1(net126),
    .A2(net185),
    .B1(net181),
    .B2(net122),
    .X(_01393_));
 sky130_fd_sc_hd__xnor2_1 _08303_ (.A(net154),
    .B(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_1 _08304_ (.A(net225),
    .B(net116),
    .Y(_01395_));
 sky130_fd_sc_hd__xnor2_1 _08305_ (.A(net150),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2b_1 _08306_ (.A_N(_01394_),
    .B(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__o22a_1 _08307_ (.A1(net138),
    .A2(net133),
    .B1(net171),
    .B2(net136),
    .X(_01398_));
 sky130_fd_sc_hd__xnor2_2 _08308_ (.A(net210),
    .B(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__o22a_1 _08309_ (.A1(net305),
    .A2(net118),
    .B1(net256),
    .B2(net90),
    .X(_01400_));
 sky130_fd_sc_hd__xnor2_2 _08310_ (.A(net258),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_1 _08311_ (.A(_01399_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__o22a_1 _08312_ (.A1(net99),
    .A2(net176),
    .B1(net173),
    .B2(net97),
    .X(_01403_));
 sky130_fd_sc_hd__xnor2_2 _08313_ (.A(net212),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__inv_2 _08314_ (.A(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__xor2_2 _08315_ (.A(_01399_),
    .B(_01401_),
    .X(_01406_));
 sky130_fd_sc_hd__a21oi_2 _08316_ (.A1(_01405_),
    .A2(_01406_),
    .B1(_01402_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _08317_ (.A(_01397_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__o22a_1 _08318_ (.A1(net141),
    .A2(net131),
    .B1(net169),
    .B2(net139),
    .X(_01409_));
 sky130_fd_sc_hd__xnor2_2 _08319_ (.A(net193),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__o22a_1 _08320_ (.A1(net179),
    .A2(net87),
    .B1(net82),
    .B2(net143),
    .X(_01411_));
 sky130_fd_sc_hd__xnor2_2 _08321_ (.A(net187),
    .B(_01411_),
    .Y(_01412_));
 sky130_fd_sc_hd__xor2_1 _08322_ (.A(_01410_),
    .B(_01412_),
    .X(_01413_));
 sky130_fd_sc_hd__o22a_1 _08323_ (.A1(net147),
    .A2(net129),
    .B1(net128),
    .B2(net145),
    .X(_01414_));
 sky130_fd_sc_hd__xnor2_1 _08324_ (.A(net166),
    .B(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2b_1 _08325_ (.A_N(_01415_),
    .B(_01413_),
    .Y(_01416_));
 sky130_fd_sc_hd__o21ai_2 _08326_ (.A1(_01410_),
    .A2(_01412_),
    .B1(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__xor2_2 _08327_ (.A(_01397_),
    .B(_01407_),
    .X(_01418_));
 sky130_fd_sc_hd__a21oi_2 _08328_ (.A1(_01417_),
    .A2(_01418_),
    .B1(_01408_),
    .Y(_01419_));
 sky130_fd_sc_hd__xnor2_2 _08329_ (.A(_01357_),
    .B(_01359_),
    .Y(_01420_));
 sky130_fd_sc_hd__xnor2_2 _08330_ (.A(_01348_),
    .B(_01350_),
    .Y(_01421_));
 sky130_fd_sc_hd__xor2_1 _08331_ (.A(_01420_),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__xnor2_1 _08332_ (.A(_01366_),
    .B(_01368_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _08333_ (.A(_01422_),
    .B(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__o21ai_2 _08334_ (.A1(_01420_),
    .A2(_01421_),
    .B1(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__xnor2_2 _08335_ (.A(_01392_),
    .B(_01419_),
    .Y(_01426_));
 sky130_fd_sc_hd__and2b_1 _08336_ (.A_N(_01426_),
    .B(_01425_),
    .X(_01427_));
 sky130_fd_sc_hd__o21ba_1 _08337_ (.A1(_01392_),
    .A2(_01419_),
    .B1_N(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__nand2b_1 _08338_ (.A_N(_01428_),
    .B(_01391_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_1 _08339_ (.A(_01390_),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__xor2_1 _08340_ (.A(_01383_),
    .B(_01384_),
    .X(_01431_));
 sky130_fd_sc_hd__nand2b_1 _08341_ (.A_N(_01431_),
    .B(_01430_),
    .Y(_01432_));
 sky130_fd_sc_hd__and3_1 _08342_ (.A(_01390_),
    .B(_01429_),
    .C(_01431_),
    .X(_01433_));
 sky130_fd_sc_hd__xor2_1 _08343_ (.A(_01430_),
    .B(_01431_),
    .X(_01434_));
 sky130_fd_sc_hd__inv_2 _08344_ (.A(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__or2_1 _08345_ (.A(_01378_),
    .B(_01379_),
    .X(_01436_));
 sky130_fd_sc_hd__nand2_1 _08346_ (.A(_01380_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__xor2_2 _08347_ (.A(_01425_),
    .B(_01426_),
    .X(_01438_));
 sky130_fd_sc_hd__nor2_1 _08348_ (.A(_01437_),
    .B(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__xnor2_2 _08349_ (.A(_01417_),
    .B(_01418_),
    .Y(_01440_));
 sky130_fd_sc_hd__o22a_1 _08350_ (.A1(net146),
    .A2(net132),
    .B1(net170),
    .B2(net141),
    .X(_01441_));
 sky130_fd_sc_hd__xnor2_1 _08351_ (.A(net193),
    .B(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__o22a_1 _08352_ (.A1(net143),
    .A2(net129),
    .B1(net127),
    .B2(net147),
    .X(_01443_));
 sky130_fd_sc_hd__xnor2_1 _08353_ (.A(net166),
    .B(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _08354_ (.A(_01442_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _08355_ (.A(net151),
    .B(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__o22a_1 _08356_ (.A1(net140),
    .A2(net134),
    .B1(net172),
    .B2(net138),
    .X(_01447_));
 sky130_fd_sc_hd__xnor2_1 _08357_ (.A(net211),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__o22a_1 _08358_ (.A1(net97),
    .A2(net257),
    .B1(net90),
    .B2(net306),
    .X(_01449_));
 sky130_fd_sc_hd__xnor2_1 _08359_ (.A(net259),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _08360_ (.A(_01448_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__o22a_1 _08361_ (.A1(net136),
    .A2(net176),
    .B1(net174),
    .B2(net99),
    .X(_01452_));
 sky130_fd_sc_hd__xnor2_1 _08362_ (.A(net213),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__inv_2 _08363_ (.A(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__xor2_1 _08364_ (.A(_01448_),
    .B(_01450_),
    .X(_01455_));
 sky130_fd_sc_hd__a21oi_1 _08365_ (.A1(_01454_),
    .A2(_01455_),
    .B1(_01451_),
    .Y(_01456_));
 sky130_fd_sc_hd__nor2_1 _08366_ (.A(net151),
    .B(_01445_),
    .Y(_01457_));
 sky130_fd_sc_hd__or2_1 _08367_ (.A(net151),
    .B(_01445_),
    .X(_01458_));
 sky130_fd_sc_hd__and2_1 _08368_ (.A(_01446_),
    .B(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__o21a_1 _08369_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01446_),
    .X(_01460_));
 sky130_fd_sc_hd__xnor2_1 _08370_ (.A(_01394_),
    .B(_01396_),
    .Y(_01461_));
 sky130_fd_sc_hd__xnor2_1 _08371_ (.A(_01404_),
    .B(_01406_),
    .Y(_01462_));
 sky130_fd_sc_hd__xnor2_1 _08372_ (.A(_01461_),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__xnor2_1 _08373_ (.A(_01413_),
    .B(_01415_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2b_1 _08374_ (.A_N(_01463_),
    .B(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__a21bo_1 _08375_ (.A1(_01461_),
    .A2(_01462_),
    .B1_N(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__xnor2_2 _08376_ (.A(_01440_),
    .B(_01460_),
    .Y(_01467_));
 sky130_fd_sc_hd__and2b_1 _08377_ (.A_N(_01467_),
    .B(_01466_),
    .X(_01468_));
 sky130_fd_sc_hd__o21bai_2 _08378_ (.A1(_01440_),
    .A2(_01460_),
    .B1_N(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__xor2_2 _08379_ (.A(_01437_),
    .B(_01438_),
    .X(_01470_));
 sky130_fd_sc_hd__and2_1 _08380_ (.A(_01469_),
    .B(_01470_),
    .X(_01471_));
 sky130_fd_sc_hd__xnor2_1 _08381_ (.A(_01391_),
    .B(_01428_),
    .Y(_01472_));
 sky130_fd_sc_hd__nor3_1 _08382_ (.A(_01439_),
    .B(_01471_),
    .C(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__or2_1 _08383_ (.A(_01422_),
    .B(_01423_),
    .X(_01474_));
 sky130_fd_sc_hd__nand2_1 _08384_ (.A(_01424_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__xor2_2 _08385_ (.A(_01466_),
    .B(_01467_),
    .X(_01476_));
 sky130_fd_sc_hd__nor2_1 _08386_ (.A(_01475_),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__xnor2_1 _08387_ (.A(_01456_),
    .B(_01459_),
    .Y(_01478_));
 sky130_fd_sc_hd__o22a_1 _08388_ (.A1(net141),
    .A2(net133),
    .B1(net172),
    .B2(net139),
    .X(_01479_));
 sky130_fd_sc_hd__xnor2_1 _08389_ (.A(_00249_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__a21oi_1 _08390_ (.A1(_00156_),
    .A2(_00157_),
    .B1(net256),
    .Y(_01481_));
 sky130_fd_sc_hd__and3_1 _08391_ (.A(net308),
    .B(_00164_),
    .C(_00165_),
    .X(_01482_));
 sky130_fd_sc_hd__o21ai_1 _08392_ (.A1(_01481_),
    .A2(_01482_),
    .B1(net261),
    .Y(_01483_));
 sky130_fd_sc_hd__or3_1 _08393_ (.A(net261),
    .B(_01481_),
    .C(_01482_),
    .X(_01484_));
 sky130_fd_sc_hd__and3_1 _08394_ (.A(_01480_),
    .B(_01483_),
    .C(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__o22a_1 _08395_ (.A1(net138),
    .A2(net176),
    .B1(net173),
    .B2(net136),
    .X(_01486_));
 sky130_fd_sc_hd__xnor2_2 _08396_ (.A(net214),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__a21o_1 _08397_ (.A1(_01483_),
    .A2(_01484_),
    .B1(_01480_),
    .X(_01488_));
 sky130_fd_sc_hd__nand2b_1 _08398_ (.A_N(_01485_),
    .B(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__a21o_1 _08399_ (.A1(_01487_),
    .A2(_01488_),
    .B1(_01485_),
    .X(_01490_));
 sky130_fd_sc_hd__o22a_1 _08400_ (.A1(net181),
    .A2(net87),
    .B1(net82),
    .B2(net180),
    .X(_01491_));
 sky130_fd_sc_hd__xnor2_1 _08401_ (.A(_06470_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(_01490_),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__o22a_1 _08403_ (.A1(net226),
    .A2(net126),
    .B1(net122),
    .B2(net184),
    .X(_01494_));
 sky130_fd_sc_hd__xnor2_1 _08404_ (.A(net154),
    .B(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__xnor2_1 _08405_ (.A(_01490_),
    .B(_01492_),
    .Y(_01496_));
 sky130_fd_sc_hd__o21a_1 _08406_ (.A1(_01495_),
    .A2(_01496_),
    .B1(_01493_),
    .X(_01497_));
 sky130_fd_sc_hd__and2b_1 _08407_ (.A_N(_01497_),
    .B(_01478_),
    .X(_01498_));
 sky130_fd_sc_hd__o22a_1 _08408_ (.A1(net148),
    .A2(net131),
    .B1(net169),
    .B2(net145),
    .X(_01499_));
 sky130_fd_sc_hd__xnor2_1 _08409_ (.A(net195),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__o22a_1 _08410_ (.A1(net180),
    .A2(net129),
    .B1(net127),
    .B2(net143),
    .X(_01501_));
 sky130_fd_sc_hd__xnor2_1 _08411_ (.A(net166),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__or2_1 _08412_ (.A(_01500_),
    .B(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__and2_1 _08413_ (.A(_01442_),
    .B(_01444_),
    .X(_01504_));
 sky130_fd_sc_hd__or2_1 _08414_ (.A(_01445_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__xnor2_1 _08415_ (.A(_01503_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__xnor2_1 _08416_ (.A(_01453_),
    .B(_01455_),
    .Y(_01507_));
 sky130_fd_sc_hd__and2b_1 _08417_ (.A_N(_01506_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__o21ba_1 _08418_ (.A1(_01503_),
    .A2(_01505_),
    .B1_N(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__xnor2_1 _08419_ (.A(_01478_),
    .B(_01497_),
    .Y(_01510_));
 sky130_fd_sc_hd__and2b_1 _08420_ (.A_N(_01509_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__or2_1 _08421_ (.A(_01498_),
    .B(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__xor2_2 _08422_ (.A(_01475_),
    .B(_01476_),
    .X(_01513_));
 sky130_fd_sc_hd__a21oi_2 _08423_ (.A1(_01512_),
    .A2(_01513_),
    .B1(_01477_),
    .Y(_01514_));
 sky130_fd_sc_hd__xnor2_2 _08424_ (.A(_01469_),
    .B(_01470_),
    .Y(_01515_));
 sky130_fd_sc_hd__or2_1 _08425_ (.A(_01514_),
    .B(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__xnor2_1 _08426_ (.A(_01514_),
    .B(_01515_),
    .Y(_01517_));
 sky130_fd_sc_hd__inv_2 _08427_ (.A(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__xnor2_1 _08428_ (.A(_01463_),
    .B(_01464_),
    .Y(_01519_));
 sky130_fd_sc_hd__xnor2_1 _08429_ (.A(_01509_),
    .B(_01510_),
    .Y(_01520_));
 sky130_fd_sc_hd__o22a_1 _08430_ (.A1(net184),
    .A2(net87),
    .B1(net82),
    .B2(net182),
    .X(_01521_));
 sky130_fd_sc_hd__xnor2_1 _08431_ (.A(net187),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__or2_1 _08432_ (.A(net226),
    .B(net122),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _08433_ (.A0(_01522_),
    .A1(net154),
    .S(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__xor2_1 _08434_ (.A(_01495_),
    .B(_01496_),
    .X(_01525_));
 sky130_fd_sc_hd__nand2b_1 _08435_ (.A_N(_01524_),
    .B(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__or2_1 _08436_ (.A(net136),
    .B(net257),
    .X(_01527_));
 sky130_fd_sc_hd__a21o_1 _08437_ (.A1(_00156_),
    .A2(_00157_),
    .B1(net305),
    .X(_01528_));
 sky130_fd_sc_hd__a21oi_1 _08438_ (.A1(_01527_),
    .A2(_01528_),
    .B1(net258),
    .Y(_01529_));
 sky130_fd_sc_hd__and3_1 _08439_ (.A(net259),
    .B(_01527_),
    .C(_01528_),
    .X(_01530_));
 sky130_fd_sc_hd__o22a_1 _08440_ (.A1(net139),
    .A2(net177),
    .B1(net173),
    .B2(net138),
    .X(_01531_));
 sky130_fd_sc_hd__xnor2_1 _08441_ (.A(net213),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__or3_2 _08442_ (.A(_01529_),
    .B(_01530_),
    .C(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__nand2_1 _08443_ (.A(_01500_),
    .B(_01502_),
    .Y(_01534_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_01503_),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _08445_ (.A(_01533_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__xor2_1 _08446_ (.A(_01533_),
    .B(_01535_),
    .X(_01537_));
 sky130_fd_sc_hd__xnor2_2 _08447_ (.A(_01487_),
    .B(_01489_),
    .Y(_01538_));
 sky130_fd_sc_hd__a21o_1 _08448_ (.A1(_01537_),
    .A2(_01538_),
    .B1(_01536_),
    .X(_01539_));
 sky130_fd_sc_hd__xnor2_1 _08449_ (.A(_01524_),
    .B(_01525_),
    .Y(_01540_));
 sky130_fd_sc_hd__a21bo_1 _08450_ (.A1(_01539_),
    .A2(_01540_),
    .B1_N(_01526_),
    .X(_01541_));
 sky130_fd_sc_hd__xnor2_1 _08451_ (.A(_01519_),
    .B(_01520_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2b_1 _08452_ (.A_N(_01542_),
    .B(_01541_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21bo_1 _08453_ (.A1(_01519_),
    .A2(_01520_),
    .B1_N(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__xor2_1 _08454_ (.A(_01512_),
    .B(_01513_),
    .X(_01545_));
 sky130_fd_sc_hd__or2_1 _08455_ (.A(_01544_),
    .B(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__xor2_1 _08456_ (.A(_01506_),
    .B(_01507_),
    .X(_01547_));
 sky130_fd_sc_hd__xnor2_1 _08457_ (.A(_01539_),
    .B(_01540_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _08458_ (.A(_01547_),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__xnor2_1 _08459_ (.A(_01547_),
    .B(_01548_),
    .Y(_01550_));
 sky130_fd_sc_hd__o22a_1 _08460_ (.A1(net145),
    .A2(net133),
    .B1(net171),
    .B2(net141),
    .X(_01551_));
 sky130_fd_sc_hd__xnor2_1 _08461_ (.A(net211),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__o22a_1 _08462_ (.A1(net182),
    .A2(net129),
    .B1(net127),
    .B2(net180),
    .X(_01553_));
 sky130_fd_sc_hd__xnor2_1 _08463_ (.A(net166),
    .B(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__or2_1 _08464_ (.A(_01552_),
    .B(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__o22a_1 _08465_ (.A1(net144),
    .A2(net131),
    .B1(net170),
    .B2(net147),
    .X(_01556_));
 sky130_fd_sc_hd__xnor2_1 _08466_ (.A(net193),
    .B(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__xnor2_1 _08467_ (.A(_01552_),
    .B(_01554_),
    .Y(_01558_));
 sky130_fd_sc_hd__o21a_1 _08468_ (.A1(_01557_),
    .A2(_01558_),
    .B1(_01555_),
    .X(_01559_));
 sky130_fd_sc_hd__xor2_1 _08469_ (.A(_01522_),
    .B(_01523_),
    .X(_01560_));
 sky130_fd_sc_hd__nand2b_1 _08470_ (.A_N(_01559_),
    .B(_01560_),
    .Y(_01561_));
 sky130_fd_sc_hd__o21ai_1 _08471_ (.A1(_01529_),
    .A2(_01530_),
    .B1(_01532_),
    .Y(_01562_));
 sky130_fd_sc_hd__o22a_1 _08472_ (.A1(net226),
    .A2(net87),
    .B1(net82),
    .B2(net184),
    .X(_01563_));
 sky130_fd_sc_hd__xnor2_1 _08473_ (.A(_06470_),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__and3_1 _08474_ (.A(_01533_),
    .B(_01562_),
    .C(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__o22a_1 _08475_ (.A1(net306),
    .A2(net136),
    .B1(net256),
    .B2(net138),
    .X(_01566_));
 sky130_fd_sc_hd__xnor2_1 _08476_ (.A(net259),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__o22a_1 _08477_ (.A1(net141),
    .A2(net177),
    .B1(net174),
    .B2(net139),
    .X(_01568_));
 sky130_fd_sc_hd__xnor2_1 _08478_ (.A(net213),
    .B(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__nor2_1 _08479_ (.A(_01567_),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__a21o_1 _08480_ (.A1(_01533_),
    .A2(_01562_),
    .B1(_01564_),
    .X(_01571_));
 sky130_fd_sc_hd__nand2b_1 _08481_ (.A_N(_01565_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__a21oi_1 _08482_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01565_),
    .Y(_01573_));
 sky130_fd_sc_hd__xnor2_1 _08483_ (.A(_01559_),
    .B(_01560_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2b_1 _08484_ (.A_N(_01573_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _08485_ (.A(_01561_),
    .B(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__and2b_1 _08486_ (.A_N(_01550_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__xnor2_1 _08487_ (.A(_01541_),
    .B(_01542_),
    .Y(_01578_));
 sky130_fd_sc_hd__o21a_1 _08488_ (.A1(_01549_),
    .A2(_01577_),
    .B1(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__nor3_1 _08489_ (.A(_01549_),
    .B(_01577_),
    .C(_01578_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_1 _08490_ (.A(_01579_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__or2_1 _08491_ (.A(_01579_),
    .B(_01580_),
    .X(_01582_));
 sky130_fd_sc_hd__xor2_1 _08492_ (.A(_01537_),
    .B(_01538_),
    .X(_01583_));
 sky130_fd_sc_hd__xnor2_1 _08493_ (.A(_01573_),
    .B(_01574_),
    .Y(_01584_));
 sky130_fd_sc_hd__xnor2_1 _08494_ (.A(_01583_),
    .B(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__xor2_1 _08495_ (.A(_01557_),
    .B(_01558_),
    .X(_01586_));
 sky130_fd_sc_hd__o22a_1 _08496_ (.A1(net147),
    .A2(net134),
    .B1(net171),
    .B2(net145),
    .X(_01587_));
 sky130_fd_sc_hd__xnor2_1 _08497_ (.A(net211),
    .B(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__o22a_1 _08498_ (.A1(net184),
    .A2(net129),
    .B1(net127),
    .B2(net182),
    .X(_01589_));
 sky130_fd_sc_hd__xnor2_1 _08499_ (.A(net168),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__or2_1 _08500_ (.A(_01588_),
    .B(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _08501_ (.A(_01588_),
    .B(_01590_),
    .Y(_01592_));
 sky130_fd_sc_hd__o22a_1 _08502_ (.A1(net180),
    .A2(net131),
    .B1(net169),
    .B2(net144),
    .X(_01593_));
 sky130_fd_sc_hd__xnor2_1 _08503_ (.A(net195),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__o21ai_1 _08504_ (.A1(_01592_),
    .A2(_01594_),
    .B1(_01591_),
    .Y(_01595_));
 sky130_fd_sc_hd__and2_1 _08505_ (.A(_01586_),
    .B(_01595_),
    .X(_01596_));
 sky130_fd_sc_hd__xor2_1 _08506_ (.A(_01586_),
    .B(_01595_),
    .X(_01597_));
 sky130_fd_sc_hd__or2_1 _08507_ (.A(net226),
    .B(net83),
    .X(_01598_));
 sky130_fd_sc_hd__xor2_1 _08508_ (.A(_01567_),
    .B(_01569_),
    .X(_01599_));
 sky130_fd_sc_hd__nor2_1 _08509_ (.A(_01598_),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__a21oi_1 _08510_ (.A1(net187),
    .A2(_01598_),
    .B1(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__a21o_1 _08511_ (.A1(_01597_),
    .A2(_01601_),
    .B1(_01596_),
    .X(_01602_));
 sky130_fd_sc_hd__nand2b_1 _08512_ (.A_N(_01585_),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21bo_1 _08513_ (.A1(_01583_),
    .A2(_01584_),
    .B1_N(_01603_),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _08514_ (.A(_01550_),
    .B(_01576_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _08515_ (.A(_01604_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__inv_2 _08516_ (.A(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__xor2_1 _08517_ (.A(_01585_),
    .B(_01602_),
    .X(_01608_));
 sky130_fd_sc_hd__xor2_1 _08518_ (.A(_01570_),
    .B(_01572_),
    .X(_01609_));
 sky130_fd_sc_hd__xnor2_1 _08519_ (.A(_01597_),
    .B(_01601_),
    .Y(_01610_));
 sky130_fd_sc_hd__or2_1 _08520_ (.A(_01609_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__xor2_1 _08521_ (.A(_01592_),
    .B(_01594_),
    .X(_01612_));
 sky130_fd_sc_hd__o22a_1 _08522_ (.A1(net144),
    .A2(net134),
    .B1(net172),
    .B2(net147),
    .X(_01613_));
 sky130_fd_sc_hd__xnor2_1 _08523_ (.A(net210),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__o22a_1 _08524_ (.A1(net305),
    .A2(net138),
    .B1(net256),
    .B2(net139),
    .X(_01615_));
 sky130_fd_sc_hd__xnor2_1 _08525_ (.A(net259),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _08526_ (.A(_01614_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__o22a_1 _08527_ (.A1(net145),
    .A2(net177),
    .B1(net173),
    .B2(net142),
    .X(_01618_));
 sky130_fd_sc_hd__xnor2_1 _08528_ (.A(net214),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_01614_),
    .B(_01616_),
    .Y(_01620_));
 sky130_fd_sc_hd__xnor2_1 _08530_ (.A(_01614_),
    .B(_01616_),
    .Y(_01621_));
 sky130_fd_sc_hd__a21o_1 _08531_ (.A1(_01619_),
    .A2(_01620_),
    .B1(_01617_),
    .X(_01622_));
 sky130_fd_sc_hd__and2_1 _08532_ (.A(_01612_),
    .B(_01622_),
    .X(_01623_));
 sky130_fd_sc_hd__o22a_1 _08533_ (.A1(net182),
    .A2(net132),
    .B1(net169),
    .B2(net180),
    .X(_01624_));
 sky130_fd_sc_hd__xnor2_1 _08534_ (.A(net193),
    .B(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__o22a_1 _08535_ (.A1(net226),
    .A2(net129),
    .B1(net127),
    .B2(net184),
    .X(_01626_));
 sky130_fd_sc_hd__xnor2_1 _08536_ (.A(net166),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _08537_ (.A(_01625_),
    .B(_01627_),
    .Y(_01628_));
 sky130_fd_sc_hd__xor2_1 _08538_ (.A(_01612_),
    .B(_01622_),
    .X(_01629_));
 sky130_fd_sc_hd__a21o_1 _08539_ (.A1(_01628_),
    .A2(_01629_),
    .B1(_01623_),
    .X(_01630_));
 sky130_fd_sc_hd__xnor2_1 _08540_ (.A(_01609_),
    .B(_01610_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand2b_1 _08541_ (.A_N(_01631_),
    .B(_01630_),
    .Y(_01632_));
 sky130_fd_sc_hd__a21oi_1 _08542_ (.A1(_01611_),
    .A2(_01632_),
    .B1(_01608_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand3_1 _08543_ (.A(_01608_),
    .B(_01611_),
    .C(_01632_),
    .Y(_01634_));
 sky130_fd_sc_hd__and2b_1 _08544_ (.A_N(_01633_),
    .B(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__xnor2_1 _08545_ (.A(_01628_),
    .B(_01629_),
    .Y(_01636_));
 sky130_fd_sc_hd__and2_1 _08546_ (.A(_01598_),
    .B(_01599_),
    .X(_01637_));
 sky130_fd_sc_hd__nor2_1 _08547_ (.A(_01600_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _08548_ (.A(_01636_),
    .B(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__xnor2_1 _08549_ (.A(_01636_),
    .B(_01638_),
    .Y(_01640_));
 sky130_fd_sc_hd__o22a_1 _08550_ (.A1(net180),
    .A2(net134),
    .B1(net172),
    .B2(net143),
    .X(_01641_));
 sky130_fd_sc_hd__xnor2_2 _08551_ (.A(net211),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__o22a_1 _08552_ (.A1(net305),
    .A2(net140),
    .B1(net256),
    .B2(net142),
    .X(_01643_));
 sky130_fd_sc_hd__xnor2_2 _08553_ (.A(net259),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _08554_ (.A(_01642_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__o22a_1 _08555_ (.A1(net148),
    .A2(net177),
    .B1(net174),
    .B2(net146),
    .X(_01646_));
 sky130_fd_sc_hd__xnor2_2 _08556_ (.A(net212),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__inv_2 _08557_ (.A(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__xor2_2 _08558_ (.A(_01642_),
    .B(_01644_),
    .X(_01649_));
 sky130_fd_sc_hd__a21oi_1 _08559_ (.A1(_01648_),
    .A2(_01649_),
    .B1(_01645_),
    .Y(_01650_));
 sky130_fd_sc_hd__xnor2_1 _08560_ (.A(_01619_),
    .B(_01621_),
    .Y(_01651_));
 sky130_fd_sc_hd__and2b_1 _08561_ (.A_N(_01650_),
    .B(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__o22a_1 _08562_ (.A1(net184),
    .A2(net132),
    .B1(net170),
    .B2(net182),
    .X(_01653_));
 sky130_fd_sc_hd__xnor2_2 _08563_ (.A(net193),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _08564_ (.A(net226),
    .B(net127),
    .Y(_01655_));
 sky130_fd_sc_hd__xnor2_2 _08565_ (.A(net168),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__and2b_1 _08566_ (.A_N(_01654_),
    .B(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__xnor2_1 _08567_ (.A(_01650_),
    .B(_01651_),
    .Y(_01658_));
 sky130_fd_sc_hd__a21oi_1 _08568_ (.A1(_01657_),
    .A2(_01658_),
    .B1(_01652_),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_1 _08569_ (.A(_01640_),
    .B(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__xnor2_1 _08570_ (.A(_01630_),
    .B(_01631_),
    .Y(_01661_));
 sky130_fd_sc_hd__nor3_1 _08571_ (.A(_01639_),
    .B(_01660_),
    .C(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__xnor2_1 _08572_ (.A(_01640_),
    .B(_01659_),
    .Y(_01663_));
 sky130_fd_sc_hd__and2_1 _08573_ (.A(_01625_),
    .B(_01627_),
    .X(_01664_));
 sky130_fd_sc_hd__or2_1 _08574_ (.A(_01628_),
    .B(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__xnor2_1 _08575_ (.A(_01657_),
    .B(_01658_),
    .Y(_01666_));
 sky130_fd_sc_hd__or2_1 _08576_ (.A(_01665_),
    .B(_01666_),
    .X(_01667_));
 sky130_fd_sc_hd__xnor2_2 _08577_ (.A(_01647_),
    .B(_01649_),
    .Y(_01668_));
 sky130_fd_sc_hd__and2b_1 _08578_ (.A_N(net168),
    .B(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__o22a_1 _08579_ (.A1(net144),
    .A2(net177),
    .B1(net174),
    .B2(net148),
    .X(_01670_));
 sky130_fd_sc_hd__xnor2_1 _08580_ (.A(net212),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__o22a_1 _08581_ (.A1(net305),
    .A2(net142),
    .B1(net256),
    .B2(net146),
    .X(_01672_));
 sky130_fd_sc_hd__xnor2_1 _08582_ (.A(net259),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__nor2_2 _08583_ (.A(_01671_),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__xnor2_2 _08584_ (.A(net168),
    .B(_01668_),
    .Y(_01675_));
 sky130_fd_sc_hd__a21o_1 _08585_ (.A1(_01674_),
    .A2(_01675_),
    .B1(_01669_),
    .X(_01676_));
 sky130_fd_sc_hd__xor2_1 _08586_ (.A(_01665_),
    .B(_01666_),
    .X(_01677_));
 sky130_fd_sc_hd__nand2_1 _08587_ (.A(_01676_),
    .B(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__a21o_1 _08588_ (.A1(_01667_),
    .A2(_01678_),
    .B1(_01663_),
    .X(_01679_));
 sky130_fd_sc_hd__nand3_1 _08589_ (.A(_01663_),
    .B(_01667_),
    .C(_01678_),
    .Y(_01680_));
 sky130_fd_sc_hd__and2_1 _08590_ (.A(_01679_),
    .B(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__xnor2_2 _08591_ (.A(_01654_),
    .B(_01656_),
    .Y(_01682_));
 sky130_fd_sc_hd__xor2_2 _08592_ (.A(_01674_),
    .B(_01675_),
    .X(_01683_));
 sky130_fd_sc_hd__nand2_1 _08593_ (.A(_01682_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__xnor2_2 _08594_ (.A(_01682_),
    .B(_01683_),
    .Y(_01685_));
 sky130_fd_sc_hd__o22a_1 _08595_ (.A1(net305),
    .A2(net145),
    .B1(net256),
    .B2(net148),
    .X(_01686_));
 sky130_fd_sc_hd__xnor2_2 _08596_ (.A(net261),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__o22a_1 _08597_ (.A1(net179),
    .A2(net176),
    .B1(net174),
    .B2(net144),
    .X(_01688_));
 sky130_fd_sc_hd__xnor2_2 _08598_ (.A(net214),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__o22a_1 _08599_ (.A1(net182),
    .A2(net133),
    .B1(net172),
    .B2(net180),
    .X(_01690_));
 sky130_fd_sc_hd__xnor2_1 _08600_ (.A(_00249_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand3_1 _08601_ (.A(_01687_),
    .B(_01689_),
    .C(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__o22a_1 _08602_ (.A1(net226),
    .A2(net131),
    .B1(net170),
    .B2(net185),
    .X(_01693_));
 sky130_fd_sc_hd__xor2_1 _08603_ (.A(net195),
    .B(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__a21o_1 _08604_ (.A1(_01687_),
    .A2(_01689_),
    .B1(_01691_),
    .X(_01695_));
 sky130_fd_sc_hd__nand3_1 _08605_ (.A(_01692_),
    .B(_01694_),
    .C(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _08606_ (.A(_01692_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__inv_2 _08607_ (.A(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__o21ai_1 _08608_ (.A1(_01685_),
    .A2(_01698_),
    .B1(_01684_),
    .Y(_01699_));
 sky130_fd_sc_hd__xor2_1 _08609_ (.A(_01676_),
    .B(_01677_),
    .X(_01700_));
 sky130_fd_sc_hd__or2_1 _08610_ (.A(_01699_),
    .B(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__xnor2_2 _08611_ (.A(_01685_),
    .B(_01698_),
    .Y(_01702_));
 sky130_fd_sc_hd__and2_1 _08612_ (.A(_01671_),
    .B(_01673_),
    .X(_01703_));
 sky130_fd_sc_hd__nor2_1 _08613_ (.A(_01674_),
    .B(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__a21o_1 _08614_ (.A1(_01692_),
    .A2(_01695_),
    .B1(_01694_),
    .X(_01705_));
 sky130_fd_sc_hd__and3_1 _08615_ (.A(_01696_),
    .B(_01704_),
    .C(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__a21oi_1 _08616_ (.A1(_01696_),
    .A2(_01705_),
    .B1(_01704_),
    .Y(_01707_));
 sky130_fd_sc_hd__nor2_1 _08617_ (.A(net226),
    .B(net169),
    .Y(_01708_));
 sky130_fd_sc_hd__o22a_1 _08618_ (.A1(net185),
    .A2(net134),
    .B1(net172),
    .B2(net182),
    .X(_01709_));
 sky130_fd_sc_hd__xnor2_2 _08619_ (.A(net210),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__mux2_1 _08620_ (.A0(net195),
    .A1(_01710_),
    .S(_01708_),
    .X(_01711_));
 sky130_fd_sc_hd__or3_1 _08621_ (.A(_01706_),
    .B(_01707_),
    .C(_01711_),
    .X(_01712_));
 sky130_fd_sc_hd__and2b_1 _08622_ (.A_N(_01706_),
    .B(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__nor2_1 _08623_ (.A(_01702_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__or2_1 _08624_ (.A(_01702_),
    .B(_01713_),
    .X(_01715_));
 sky130_fd_sc_hd__xnor2_2 _08625_ (.A(_01702_),
    .B(_01713_),
    .Y(_01716_));
 sky130_fd_sc_hd__o21ai_1 _08626_ (.A1(_01706_),
    .A2(_01707_),
    .B1(_01711_),
    .Y(_01717_));
 sky130_fd_sc_hd__xor2_2 _08627_ (.A(_01687_),
    .B(_01689_),
    .X(_01718_));
 sky130_fd_sc_hd__xor2_2 _08628_ (.A(_01708_),
    .B(_01710_),
    .X(_01719_));
 sky130_fd_sc_hd__and2b_1 _08629_ (.A_N(_01719_),
    .B(_01718_),
    .X(_01720_));
 sky130_fd_sc_hd__o22a_1 _08630_ (.A1(net182),
    .A2(net177),
    .B1(net174),
    .B2(net179),
    .X(_01721_));
 sky130_fd_sc_hd__xnor2_1 _08631_ (.A(net213),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand3_1 _08632_ (.A(_00140_),
    .B(_00141_),
    .C(_00239_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21o_1 _08633_ (.A1(_06545_),
    .A2(_06546_),
    .B1(_04428_),
    .X(_01724_));
 sky130_fd_sc_hd__a21oi_2 _08634_ (.A1(_01723_),
    .A2(_01724_),
    .B1(net260),
    .Y(_01725_));
 sky130_fd_sc_hd__and3_1 _08635_ (.A(net260),
    .B(_01723_),
    .C(_01724_),
    .X(_01726_));
 sky130_fd_sc_hd__or3_4 _08636_ (.A(_01722_),
    .B(_01725_),
    .C(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__xor2_2 _08637_ (.A(_01718_),
    .B(_01719_),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_1 _08638_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__a211oi_1 _08639_ (.A1(_01712_),
    .A2(_01717_),
    .B1(_01720_),
    .C1(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__o21ai_1 _08640_ (.A1(_01725_),
    .A2(_01726_),
    .B1(_01722_),
    .Y(_01731_));
 sky130_fd_sc_hd__o22a_1 _08641_ (.A1(net226),
    .A2(net134),
    .B1(net172),
    .B2(net185),
    .X(_01732_));
 sky130_fd_sc_hd__xnor2_1 _08642_ (.A(_00249_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand3_1 _08643_ (.A(_01727_),
    .B(_01731_),
    .C(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__a32o_1 _08644_ (.A1(net308),
    .A2(_00140_),
    .A3(_00141_),
    .B1(_00239_),
    .B2(_06565_),
    .X(_01735_));
 sky130_fd_sc_hd__xnor2_2 _08645_ (.A(net261),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__o22a_1 _08646_ (.A1(net185),
    .A2(net177),
    .B1(net174),
    .B2(net182),
    .X(_01737_));
 sky130_fd_sc_hd__xnor2_1 _08647_ (.A(net212),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _08648_ (.A(_01736_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__a21o_1 _08649_ (.A1(_01727_),
    .A2(_01731_),
    .B1(_01733_),
    .X(_01740_));
 sky130_fd_sc_hd__and3_1 _08650_ (.A(_01734_),
    .B(_01739_),
    .C(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__a31o_1 _08651_ (.A1(_01727_),
    .A2(_01731_),
    .A3(_01733_),
    .B1(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__xor2_2 _08652_ (.A(_01727_),
    .B(_01728_),
    .X(_01743_));
 sky130_fd_sc_hd__xnor2_1 _08653_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__a21oi_1 _08654_ (.A1(_01734_),
    .A2(_01740_),
    .B1(_01739_),
    .Y(_01745_));
 sky130_fd_sc_hd__xor2_1 _08655_ (.A(_01736_),
    .B(_01738_),
    .X(_01746_));
 sky130_fd_sc_hd__or2_1 _08656_ (.A(net226),
    .B(net171),
    .X(_01747_));
 sky130_fd_sc_hd__nor2_1 _08657_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__a21o_1 _08658_ (.A1(net210),
    .A2(_01747_),
    .B1(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__o21a_1 _08659_ (.A1(_01741_),
    .A2(_01745_),
    .B1(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__o21ai_1 _08660_ (.A1(_01741_),
    .A2(_01745_),
    .B1(_01749_),
    .Y(_01751_));
 sky130_fd_sc_hd__o22a_1 _08661_ (.A1(net226),
    .A2(net177),
    .B1(net174),
    .B2(net185),
    .X(_01752_));
 sky130_fd_sc_hd__xnor2_1 _08662_ (.A(net212),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__o22a_1 _08663_ (.A1(net305),
    .A2(net179),
    .B1(net257),
    .B2(net181),
    .X(_01754_));
 sky130_fd_sc_hd__xnor2_1 _08664_ (.A(net258),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_1 _08665_ (.A(_01753_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__xor2_1 _08666_ (.A(_01746_),
    .B(_01747_),
    .X(_01757_));
 sky130_fd_sc_hd__and2b_1 _08667_ (.A_N(_01757_),
    .B(_01756_),
    .X(_01758_));
 sky130_fd_sc_hd__or3_1 _08668_ (.A(_01753_),
    .B(_01755_),
    .C(_01757_),
    .X(_01759_));
 sky130_fd_sc_hd__and2b_1 _08669_ (.A_N(_01756_),
    .B(_01757_),
    .X(_01760_));
 sky130_fd_sc_hd__nor2_1 _08670_ (.A(_01758_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__o22a_1 _08671_ (.A1(net305),
    .A2(net181),
    .B1(net257),
    .B2(net185),
    .X(_01762_));
 sky130_fd_sc_hd__xnor2_1 _08672_ (.A(net259),
    .B(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _08673_ (.A(net226),
    .B(net174),
    .Y(_01764_));
 sky130_fd_sc_hd__or2_1 _08674_ (.A(net213),
    .B(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__nand2_1 _08675_ (.A(net212),
    .B(_01764_),
    .Y(_01766_));
 sky130_fd_sc_hd__a21oi_1 _08676_ (.A1(_01765_),
    .A2(_01766_),
    .B1(_01763_),
    .Y(_01767_));
 sky130_fd_sc_hd__and3_1 _08677_ (.A(_01763_),
    .B(_01765_),
    .C(_01766_),
    .X(_01768_));
 sky130_fd_sc_hd__xnor2_1 _08678_ (.A(_01763_),
    .B(_01764_),
    .Y(_01769_));
 sky130_fd_sc_hd__a22o_1 _08679_ (.A1(net308),
    .A2(_06526_),
    .B1(_00239_),
    .B2(net224),
    .X(_01770_));
 sky130_fd_sc_hd__or2_2 _08680_ (.A(_06408_),
    .B(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__nor2_1 _08681_ (.A(net259),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _08682_ (.A(_01769_),
    .B(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__xor2_1 _08683_ (.A(_01753_),
    .B(_01755_),
    .X(_01774_));
 sky130_fd_sc_hd__inv_2 _08684_ (.A(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__xnor2_1 _08685_ (.A(_01767_),
    .B(_01774_),
    .Y(_01776_));
 sky130_fd_sc_hd__o21ba_1 _08686_ (.A1(net213),
    .A2(_01768_),
    .B1_N(_01767_),
    .X(_01777_));
 sky130_fd_sc_hd__o22a_1 _08687_ (.A1(_01773_),
    .A2(_01776_),
    .B1(_01777_),
    .B2(_01775_),
    .X(_01778_));
 sky130_fd_sc_hd__o21ai_2 _08688_ (.A1(_01760_),
    .A2(_01778_),
    .B1(_01759_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor3_1 _08689_ (.A(_01741_),
    .B(_01745_),
    .C(_01749_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _08690_ (.A(_01750_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__a21oi_1 _08691_ (.A1(_01751_),
    .A2(_01779_),
    .B1(_01780_),
    .Y(_01782_));
 sky130_fd_sc_hd__o211a_1 _08692_ (.A1(_01720_),
    .A2(_01729_),
    .B1(_01712_),
    .C1(_01717_),
    .X(_01783_));
 sky130_fd_sc_hd__a221o_1 _08693_ (.A1(_01742_),
    .A2(_01743_),
    .B1(_01751_),
    .B2(_01779_),
    .C1(_01780_),
    .X(_01784_));
 sky130_fd_sc_hd__o21ai_1 _08694_ (.A1(_01742_),
    .A2(_01743_),
    .B1(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _08695_ (.A(_01730_),
    .B(_01783_),
    .Y(_01786_));
 sky130_fd_sc_hd__o21ba_2 _08696_ (.A1(_01730_),
    .A2(_01785_),
    .B1_N(_01783_),
    .X(_01787_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_01699_),
    .B(_01700_),
    .Y(_01788_));
 sky130_fd_sc_hd__o211ai_2 _08698_ (.A1(_01716_),
    .A2(_01787_),
    .B1(_01788_),
    .C1(_01715_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(_01701_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__o21a_1 _08700_ (.A1(_01639_),
    .A2(_01660_),
    .B1(_01661_),
    .X(_01791_));
 sky130_fd_sc_hd__o21ai_1 _08701_ (.A1(_01639_),
    .A2(_01660_),
    .B1(_01661_),
    .Y(_01792_));
 sky130_fd_sc_hd__a21oi_1 _08702_ (.A1(_01679_),
    .A2(_01792_),
    .B1(_01662_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _08703_ (.A(_01662_),
    .B(_01791_),
    .Y(_01794_));
 sky130_fd_sc_hd__a41o_1 _08704_ (.A1(_01681_),
    .A2(_01701_),
    .A3(_01789_),
    .A4(_01794_),
    .B1(_01793_),
    .X(_01795_));
 sky130_fd_sc_hd__and2_1 _08705_ (.A(_01604_),
    .B(_01605_),
    .X(_01796_));
 sky130_fd_sc_hd__a211o_1 _08706_ (.A1(_01635_),
    .A2(_01795_),
    .B1(_01796_),
    .C1(_01633_),
    .X(_01797_));
 sky130_fd_sc_hd__nand2_1 _08707_ (.A(_01607_),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__and2_1 _08708_ (.A(_01544_),
    .B(_01545_),
    .X(_01799_));
 sky130_fd_sc_hd__a311o_1 _08709_ (.A1(_01581_),
    .A2(_01607_),
    .A3(_01797_),
    .B1(_01799_),
    .C1(_01579_),
    .X(_01800_));
 sky130_fd_sc_hd__xnor2_1 _08710_ (.A(_01544_),
    .B(_01545_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(_01546_),
    .B(_01800_),
    .Y(_01802_));
 sky130_fd_sc_hd__o21ai_2 _08712_ (.A1(_01439_),
    .A2(_01471_),
    .B1(_01472_),
    .Y(_01803_));
 sky130_fd_sc_hd__a21oi_1 _08713_ (.A1(_01516_),
    .A2(_01803_),
    .B1(_01473_),
    .Y(_01804_));
 sky130_fd_sc_hd__and2b_1 _08714_ (.A_N(_01473_),
    .B(_01803_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2b_1 _08715_ (.A_N(_01473_),
    .B(_01803_),
    .Y(_01806_));
 sky130_fd_sc_hd__a41o_1 _08716_ (.A1(_01518_),
    .A2(_01546_),
    .A3(_01800_),
    .A4(_01805_),
    .B1(_01804_),
    .X(_01807_));
 sky130_fd_sc_hd__o21ai_1 _08717_ (.A1(_01346_),
    .A2(_01385_),
    .B1(_01343_),
    .Y(_01808_));
 sky130_fd_sc_hd__a21oi_1 _08718_ (.A1(_01432_),
    .A2(_01808_),
    .B1(_01386_),
    .Y(_01809_));
 sky130_fd_sc_hd__and2b_1 _08719_ (.A_N(_01386_),
    .B(_01808_),
    .X(_01810_));
 sky130_fd_sc_hd__a31o_1 _08720_ (.A1(_01435_),
    .A2(_01807_),
    .A3(_01810_),
    .B1(_01809_),
    .X(_01811_));
 sky130_fd_sc_hd__o22a_1 _08721_ (.A1(net126),
    .A2(net141),
    .B1(net139),
    .B2(net122),
    .X(_01812_));
 sky130_fd_sc_hd__xnor2_2 _08722_ (.A(net154),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__o22a_1 _08723_ (.A1(net75),
    .A2(net147),
    .B1(net145),
    .B2(net116),
    .X(_01814_));
 sky130_fd_sc_hd__xnor2_2 _08724_ (.A(net150),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _08725_ (.A(_01813_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__xnor2_1 _08726_ (.A(_01813_),
    .B(_01815_),
    .Y(_01817_));
 sky130_fd_sc_hd__o22a_1 _08727_ (.A1(net120),
    .A2(net176),
    .B1(net173),
    .B2(net84),
    .X(_01818_));
 sky130_fd_sc_hd__xnor2_1 _08728_ (.A(net212),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__inv_2 _08729_ (.A(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__o32a_1 _08730_ (.A1(net305),
    .A2(_00310_),
    .A3(_00311_),
    .B1(net256),
    .B2(net79),
    .X(_01821_));
 sky130_fd_sc_hd__xnor2_2 _08731_ (.A(net258),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__o22a_1 _08732_ (.A1(net114),
    .A2(net133),
    .B1(net171),
    .B2(net124),
    .X(_01823_));
 sky130_fd_sc_hd__xnor2_2 _08733_ (.A(net210),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _08734_ (.A(_01822_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__xor2_2 _08735_ (.A(_01822_),
    .B(_01824_),
    .X(_01826_));
 sky130_fd_sc_hd__xnor2_1 _08736_ (.A(_01819_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__and2b_1 _08737_ (.A_N(_01817_),
    .B(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__xnor2_1 _08738_ (.A(_01817_),
    .B(_01827_),
    .Y(_01829_));
 sky130_fd_sc_hd__o22a_1 _08739_ (.A1(net138),
    .A2(net87),
    .B1(net82),
    .B2(net136),
    .X(_01830_));
 sky130_fd_sc_hd__xnor2_1 _08740_ (.A(net187),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__o22a_1 _08741_ (.A1(net90),
    .A2(net131),
    .B1(net169),
    .B2(net118),
    .X(_01832_));
 sky130_fd_sc_hd__xnor2_1 _08742_ (.A(net193),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__xor2_1 _08743_ (.A(_01831_),
    .B(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__o22a_1 _08744_ (.A1(net99),
    .A2(net129),
    .B1(net127),
    .B2(net97),
    .X(_01835_));
 sky130_fd_sc_hd__xnor2_1 _08745_ (.A(net166),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__and2b_1 _08746_ (.A_N(_01836_),
    .B(_01834_),
    .X(_01837_));
 sky130_fd_sc_hd__and2b_1 _08747_ (.A_N(_01834_),
    .B(_01836_),
    .X(_01838_));
 sky130_fd_sc_hd__nor2_1 _08748_ (.A(_01837_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__xnor2_1 _08749_ (.A(_01829_),
    .B(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__o22a_1 _08750_ (.A1(net179),
    .A2(net69),
    .B1(net95),
    .B2(net143),
    .X(_01841_));
 sky130_fd_sc_hd__xnor2_1 _08751_ (.A(net101),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _08752_ (.A(net225),
    .B(net67),
    .Y(_01843_));
 sky130_fd_sc_hd__xnor2_1 _08753_ (.A(net104),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__and2b_1 _08754_ (.A_N(_01844_),
    .B(_01842_),
    .X(_01845_));
 sky130_fd_sc_hd__and2b_1 _08755_ (.A_N(_01842_),
    .B(_01844_),
    .X(_01846_));
 sky130_fd_sc_hd__nor2_1 _08756_ (.A(_01845_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__o22a_1 _08757_ (.A1(net184),
    .A2(net21),
    .B1(net65),
    .B2(net181),
    .X(_01848_));
 sky130_fd_sc_hd__xnor2_1 _08758_ (.A(net92),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__xnor2_1 _08759_ (.A(_01847_),
    .B(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _08760_ (.A(_01840_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(_01840_),
    .B(_01850_),
    .Y(_01852_));
 sky130_fd_sc_hd__and2b_1 _08762_ (.A_N(_01851_),
    .B(_01852_),
    .X(_01853_));
 sky130_fd_sc_hd__xnor2_1 _08763_ (.A(net104),
    .B(_01186_),
    .Y(_01854_));
 sky130_fd_sc_hd__a21oi_1 _08764_ (.A1(_01196_),
    .A2(_01198_),
    .B1(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__and3_1 _08765_ (.A(_01196_),
    .B(_01198_),
    .C(_01854_),
    .X(_01856_));
 sky130_fd_sc_hd__nor2_2 _08766_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__xnor2_4 _08767_ (.A(_01853_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__a32o_1 _08768_ (.A1(_01200_),
    .A2(_01201_),
    .A3(_01211_),
    .B1(_01212_),
    .B2(_01229_),
    .X(_01859_));
 sky130_fd_sc_hd__a21bo_1 _08769_ (.A1(_01226_),
    .A2(_01228_),
    .B1_N(_01225_),
    .X(_01860_));
 sky130_fd_sc_hd__a21oi_2 _08770_ (.A1(_01189_),
    .A2(_01199_),
    .B1(_01188_),
    .Y(_01861_));
 sky130_fd_sc_hd__o21a_1 _08771_ (.A1(_01204_),
    .A2(_01210_),
    .B1(_01209_),
    .X(_01862_));
 sky130_fd_sc_hd__nor2_1 _08772_ (.A(_01861_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__nand2_1 _08773_ (.A(_01861_),
    .B(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__xnor2_1 _08774_ (.A(_01861_),
    .B(_01862_),
    .Y(_01865_));
 sky130_fd_sc_hd__xnor2_2 _08775_ (.A(_01860_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__o21a_1 _08776_ (.A1(_01293_),
    .A2(_01297_),
    .B1(_01296_),
    .X(_01867_));
 sky130_fd_sc_hd__and2b_1 _08777_ (.A_N(_01867_),
    .B(_01866_),
    .X(_01868_));
 sky130_fd_sc_hd__xnor2_2 _08778_ (.A(_01866_),
    .B(_01867_),
    .Y(_01869_));
 sky130_fd_sc_hd__xnor2_2 _08779_ (.A(_01859_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__xnor2_2 _08780_ (.A(_01858_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21o_1 _08781_ (.A1(_01259_),
    .A2(_01301_),
    .B1(_01300_),
    .X(_01872_));
 sky130_fd_sc_hd__nand2b_1 _08782_ (.A_N(_01871_),
    .B(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__xnor2_2 _08783_ (.A(_01871_),
    .B(_01872_),
    .Y(_01874_));
 sky130_fd_sc_hd__a21oi_1 _08784_ (.A1(_01304_),
    .A2(_01342_),
    .B1(_01303_),
    .Y(_01875_));
 sky130_fd_sc_hd__and2b_1 _08785_ (.A_N(_01875_),
    .B(_01874_),
    .X(_01876_));
 sky130_fd_sc_hd__nand2b_1 _08786_ (.A_N(_01875_),
    .B(_01874_),
    .Y(_01877_));
 sky130_fd_sc_hd__and2b_1 _08787_ (.A_N(_01874_),
    .B(_01875_),
    .X(_01878_));
 sky130_fd_sc_hd__nor2_1 _08788_ (.A(_01876_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__o21ai_4 _08789_ (.A1(_01858_),
    .A2(_01870_),
    .B1(_01873_),
    .Y(_01880_));
 sky130_fd_sc_hd__a21o_2 _08790_ (.A1(_01859_),
    .A2(_01869_),
    .B1(_01868_),
    .X(_01881_));
 sky130_fd_sc_hd__o21ba_1 _08791_ (.A1(_01831_),
    .A2(_01833_),
    .B1_N(_01837_),
    .X(_01882_));
 sky130_fd_sc_hd__a21oi_2 _08792_ (.A1(_01820_),
    .A2(_01826_),
    .B1(_01825_),
    .Y(_01883_));
 sky130_fd_sc_hd__xnor2_1 _08793_ (.A(_01816_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2b_1 _08794_ (.A_N(_01882_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__xnor2_1 _08795_ (.A(_01882_),
    .B(_01884_),
    .Y(_01886_));
 sky130_fd_sc_hd__o22a_1 _08796_ (.A1(net143),
    .A2(net69),
    .B1(net95),
    .B2(net147),
    .X(_01887_));
 sky130_fd_sc_hd__xnor2_1 _08797_ (.A(net101),
    .B(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__o32a_1 _08798_ (.A1(net225),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net67),
    .B2(net184),
    .X(_01889_));
 sky130_fd_sc_hd__xnor2_1 _08799_ (.A(net104),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__and2_1 _08800_ (.A(_01888_),
    .B(_01890_),
    .X(_01891_));
 sky130_fd_sc_hd__xor2_1 _08801_ (.A(_01888_),
    .B(_01890_),
    .X(_01892_));
 sky130_fd_sc_hd__o22a_1 _08802_ (.A1(net181),
    .A2(net21),
    .B1(net65),
    .B2(net179),
    .X(_01893_));
 sky130_fd_sc_hd__xnor2_1 _08803_ (.A(net92),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__and2_1 _08804_ (.A(_01892_),
    .B(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__nor2_1 _08805_ (.A(_01892_),
    .B(_01894_),
    .Y(_01896_));
 sky130_fd_sc_hd__or2_1 _08806_ (.A(_01895_),
    .B(_01896_),
    .X(_01897_));
 sky130_fd_sc_hd__and2b_1 _08807_ (.A_N(_01146_),
    .B(_01148_),
    .X(_01898_));
 sky130_fd_sc_hd__nor2_1 _08808_ (.A(_01149_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__xor2_1 _08809_ (.A(_01154_),
    .B(_01156_),
    .X(_01900_));
 sky130_fd_sc_hd__a21o_1 _08810_ (.A1(_01133_),
    .A2(_01136_),
    .B1(_01135_),
    .X(_01901_));
 sky130_fd_sc_hd__nand3_1 _08811_ (.A(_01137_),
    .B(_01900_),
    .C(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__a21o_1 _08812_ (.A1(_01137_),
    .A2(_01901_),
    .B1(_01900_),
    .X(_01903_));
 sky130_fd_sc_hd__and3_1 _08813_ (.A(_01899_),
    .B(_01902_),
    .C(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__a21oi_1 _08814_ (.A1(_01902_),
    .A2(_01903_),
    .B1(_01899_),
    .Y(_01905_));
 sky130_fd_sc_hd__or3_1 _08815_ (.A(_01897_),
    .B(_01904_),
    .C(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__o21ai_1 _08816_ (.A1(_01904_),
    .A2(_01905_),
    .B1(_01897_),
    .Y(_01907_));
 sky130_fd_sc_hd__and3_1 _08817_ (.A(_01886_),
    .B(_01906_),
    .C(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__a21oi_1 _08818_ (.A1(_01906_),
    .A2(_01907_),
    .B1(_01886_),
    .Y(_01909_));
 sky130_fd_sc_hd__nor2_1 _08819_ (.A(_01908_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__a21oi_2 _08820_ (.A1(_01852_),
    .A2(_01857_),
    .B1(_01851_),
    .Y(_01911_));
 sky130_fd_sc_hd__a21o_1 _08821_ (.A1(net104),
    .A2(_01186_),
    .B1(_01855_),
    .X(_01912_));
 sky130_fd_sc_hd__a21oi_2 _08822_ (.A1(_01829_),
    .A2(_01839_),
    .B1(_01828_),
    .Y(_01913_));
 sky130_fd_sc_hd__a21oi_2 _08823_ (.A1(_01847_),
    .A2(_01849_),
    .B1(_01845_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _08824_ (.A(_01913_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__xor2_2 _08825_ (.A(_01913_),
    .B(_01914_),
    .X(_01916_));
 sky130_fd_sc_hd__xnor2_2 _08826_ (.A(_01912_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a21o_1 _08827_ (.A1(_01860_),
    .A2(_01864_),
    .B1(_01863_),
    .X(_01918_));
 sky130_fd_sc_hd__and2b_1 _08828_ (.A_N(_01917_),
    .B(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__xnor2_2 _08829_ (.A(_01917_),
    .B(_01918_),
    .Y(_01920_));
 sky130_fd_sc_hd__and2b_1 _08830_ (.A_N(_01911_),
    .B(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__xnor2_2 _08831_ (.A(_01911_),
    .B(_01920_),
    .Y(_01922_));
 sky130_fd_sc_hd__and2_1 _08832_ (.A(_01910_),
    .B(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__or2_1 _08833_ (.A(_01910_),
    .B(_01922_),
    .X(_01924_));
 sky130_fd_sc_hd__xnor2_2 _08834_ (.A(_01910_),
    .B(_01922_),
    .Y(_01925_));
 sky130_fd_sc_hd__xnor2_4 _08835_ (.A(_01881_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _08836_ (.A(_01880_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_01880_),
    .B(_01926_),
    .Y(_01928_));
 sky130_fd_sc_hd__xor2_2 _08838_ (.A(_01880_),
    .B(_01926_),
    .X(_01929_));
 sky130_fd_sc_hd__and2_1 _08839_ (.A(_01879_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__a21boi_1 _08840_ (.A1(_01880_),
    .A2(_01926_),
    .B1_N(_01877_),
    .Y(_01931_));
 sky130_fd_sc_hd__o2bb2a_1 _08841_ (.A1_N(_01811_),
    .A2_N(_01930_),
    .B1(_01931_),
    .B2(_01928_),
    .X(_01932_));
 sky130_fd_sc_hd__o21ai_1 _08842_ (.A1(_01122_),
    .A2(_01123_),
    .B1(_01124_),
    .Y(_01933_));
 sky130_fd_sc_hd__o211ai_1 _08843_ (.A1(net225),
    .A2(net73),
    .B1(_01133_),
    .C1(_01137_),
    .Y(_01934_));
 sky130_fd_sc_hd__and2_1 _08844_ (.A(_01138_),
    .B(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__and3_1 _08845_ (.A(_01125_),
    .B(_01933_),
    .C(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__a21oi_1 _08846_ (.A1(_01125_),
    .A2(_01933_),
    .B1(_01935_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_2 _08847_ (.A(_01936_),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__xnor2_4 _08848_ (.A(_01157_),
    .B(_01158_),
    .Y(_01939_));
 sky130_fd_sc_hd__xnor2_4 _08849_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__a21bo_2 _08850_ (.A1(_01886_),
    .A2(_01907_),
    .B1_N(_01906_),
    .X(_01941_));
 sky130_fd_sc_hd__a21o_1 _08851_ (.A1(_01912_),
    .A2(_01916_),
    .B1(_01915_),
    .X(_01942_));
 sky130_fd_sc_hd__o31ai_4 _08852_ (.A1(_01813_),
    .A2(_01815_),
    .A3(_01883_),
    .B1(_01885_),
    .Y(_01943_));
 sky130_fd_sc_hd__or2_1 _08853_ (.A(_01891_),
    .B(_01895_),
    .X(_01944_));
 sky130_fd_sc_hd__a21boi_2 _08854_ (.A1(_01899_),
    .A2(_01903_),
    .B1_N(_01902_),
    .Y(_01945_));
 sky130_fd_sc_hd__o21ba_1 _08855_ (.A1(_01891_),
    .A2(_01895_),
    .B1_N(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__nand2b_1 _08856_ (.A_N(_01944_),
    .B(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__xor2_1 _08857_ (.A(_01944_),
    .B(_01945_),
    .X(_01948_));
 sky130_fd_sc_hd__xnor2_2 _08858_ (.A(_01943_),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__xnor2_2 _08859_ (.A(_01942_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__and2b_1 _08860_ (.A_N(_01950_),
    .B(_01941_),
    .X(_01951_));
 sky130_fd_sc_hd__xnor2_4 _08861_ (.A(_01941_),
    .B(_01950_),
    .Y(_01952_));
 sky130_fd_sc_hd__and2_1 _08862_ (.A(_01940_),
    .B(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__xor2_4 _08863_ (.A(_01940_),
    .B(_01952_),
    .X(_01954_));
 sky130_fd_sc_hd__or2_2 _08864_ (.A(_01919_),
    .B(_01921_),
    .X(_01955_));
 sky130_fd_sc_hd__xnor2_4 _08865_ (.A(_01954_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__a21oi_4 _08866_ (.A1(_01881_),
    .A2(_01924_),
    .B1(_01923_),
    .Y(_01957_));
 sky130_fd_sc_hd__or2_1 _08867_ (.A(_01956_),
    .B(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__and2_1 _08868_ (.A(_01956_),
    .B(_01957_),
    .X(_01959_));
 sky130_fd_sc_hd__xor2_4 _08869_ (.A(_01956_),
    .B(_01957_),
    .X(_01960_));
 sky130_fd_sc_hd__a21o_1 _08870_ (.A1(_01954_),
    .A2(_01955_),
    .B1(_01953_),
    .X(_01961_));
 sky130_fd_sc_hd__a21o_1 _08871_ (.A1(_01942_),
    .A2(_01949_),
    .B1(_01951_),
    .X(_01962_));
 sky130_fd_sc_hd__xnor2_2 _08872_ (.A(_01166_),
    .B(_01167_),
    .Y(_01963_));
 sky130_fd_sc_hd__o21ba_1 _08873_ (.A1(_01937_),
    .A2(_01939_),
    .B1_N(_01936_),
    .X(_01964_));
 sky130_fd_sc_hd__xnor2_2 _08874_ (.A(_01159_),
    .B(_01160_),
    .Y(_01965_));
 sky130_fd_sc_hd__a21oi_2 _08875_ (.A1(_01943_),
    .A2(_01947_),
    .B1(_01946_),
    .Y(_01966_));
 sky130_fd_sc_hd__xor2_2 _08876_ (.A(_01965_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__nand2b_1 _08877_ (.A_N(_01964_),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__xnor2_2 _08878_ (.A(_01964_),
    .B(_01967_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(_01963_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__xor2_2 _08880_ (.A(_01963_),
    .B(_01969_),
    .X(_01971_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(_01962_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__xnor2_2 _08882_ (.A(_01962_),
    .B(_01971_),
    .Y(_01973_));
 sky130_fd_sc_hd__and2b_1 _08883_ (.A_N(_01961_),
    .B(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__nand2b_1 _08884_ (.A_N(_01973_),
    .B(_01961_),
    .Y(_01975_));
 sky130_fd_sc_hd__xnor2_2 _08885_ (.A(_01961_),
    .B(_01973_),
    .Y(_01976_));
 sky130_fd_sc_hd__and2_1 _08886_ (.A(_01960_),
    .B(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__and4bb_1 _08887_ (.A_N(_01928_),
    .B_N(_01931_),
    .C(_01960_),
    .D(_01976_),
    .X(_01978_));
 sky130_fd_sc_hd__o21ai_2 _08888_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01968_),
    .Y(_01979_));
 sky130_fd_sc_hd__a21o_1 _08889_ (.A1(_01060_),
    .A2(_01061_),
    .B1(_01063_),
    .X(_01980_));
 sky130_fd_sc_hd__and2_1 _08890_ (.A(_01064_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__xnor2_1 _08891_ (.A(_01168_),
    .B(_01169_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_01981_),
    .B(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_1 _08893_ (.A(_01981_),
    .B(_01982_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2b_1 _08894_ (.A_N(_01984_),
    .B(_01979_),
    .Y(_01985_));
 sky130_fd_sc_hd__xor2_1 _08895_ (.A(_01979_),
    .B(_01984_),
    .X(_01986_));
 sky130_fd_sc_hd__a21oi_1 _08896_ (.A1(_01970_),
    .A2(_01972_),
    .B1(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__a21o_1 _08897_ (.A1(_01970_),
    .A2(_01972_),
    .B1(_01986_),
    .X(_01988_));
 sky130_fd_sc_hd__and3_1 _08898_ (.A(_01970_),
    .B(_01972_),
    .C(_01986_),
    .X(_01989_));
 sky130_fd_sc_hd__nor2_2 _08899_ (.A(_01987_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__xor2_1 _08900_ (.A(_01171_),
    .B(_01172_),
    .X(_01991_));
 sky130_fd_sc_hd__and3_1 _08901_ (.A(_01983_),
    .B(_01985_),
    .C(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__a21o_1 _08902_ (.A1(_01983_),
    .A2(_01985_),
    .B1(_01991_),
    .X(_01993_));
 sky130_fd_sc_hd__and2b_1 _08903_ (.A_N(_01992_),
    .B(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__nand2_1 _08904_ (.A(_01990_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__a21o_1 _08905_ (.A1(_01988_),
    .A2(_01993_),
    .B1(_01992_),
    .X(_01996_));
 sky130_fd_sc_hd__a21oi_1 _08906_ (.A1(_01958_),
    .A2(_01975_),
    .B1(_01974_),
    .Y(_01997_));
 sky130_fd_sc_hd__a311oi_4 _08907_ (.A1(_01811_),
    .A2(_01930_),
    .A3(_01977_),
    .B1(_01978_),
    .C1(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__o21ai_4 _08908_ (.A1(_01995_),
    .A2(_01998_),
    .B1(_01996_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_1 _08909_ (.A(_01115_),
    .B(_01174_),
    .Y(_02000_));
 sky130_fd_sc_hd__and2_1 _08910_ (.A(_01175_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__xor2_1 _08911_ (.A(_01071_),
    .B(_01113_),
    .X(_02002_));
 sky130_fd_sc_hd__xnor2_1 _08912_ (.A(_01071_),
    .B(_01113_),
    .Y(_02003_));
 sky130_fd_sc_hd__a32o_2 _08913_ (.A1(_01999_),
    .A2(_02001_),
    .A3(_02002_),
    .B1(_01176_),
    .B2(_01114_),
    .X(_02004_));
 sky130_fd_sc_hd__a21o_2 _08914_ (.A1(_01072_),
    .A2(_01112_),
    .B1(_01111_),
    .X(_02005_));
 sky130_fd_sc_hd__a21bo_2 _08915_ (.A1(_01101_),
    .A2(_01107_),
    .B1_N(_01109_),
    .X(_02006_));
 sky130_fd_sc_hd__xnor2_1 _08916_ (.A(_00756_),
    .B(_00757_),
    .Y(_02007_));
 sky130_fd_sc_hd__and2b_1 _08917_ (.A_N(_00714_),
    .B(_00716_),
    .X(_02008_));
 sky130_fd_sc_hd__or2_1 _08918_ (.A(_00717_),
    .B(_02008_),
    .X(_02009_));
 sky130_fd_sc_hd__xnor2_2 _08919_ (.A(_00722_),
    .B(_00724_),
    .Y(_02010_));
 sky130_fd_sc_hd__xor2_1 _08920_ (.A(_02009_),
    .B(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__nand2_1 _08921_ (.A(_02007_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__or2_1 _08922_ (.A(_02007_),
    .B(_02011_),
    .X(_02013_));
 sky130_fd_sc_hd__and2_2 _08923_ (.A(_02012_),
    .B(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__a21o_1 _08924_ (.A1(_01080_),
    .A2(_01098_),
    .B1(_01096_),
    .X(_02015_));
 sky130_fd_sc_hd__nand2_2 _08925_ (.A(_01076_),
    .B(_01079_),
    .Y(_02016_));
 sky130_fd_sc_hd__o32a_2 _08926_ (.A1(_00736_),
    .A2(_01081_),
    .A3(_01087_),
    .B1(_01086_),
    .B2(_01085_),
    .X(_02017_));
 sky130_fd_sc_hd__a31oi_4 _08927_ (.A1(_00390_),
    .A2(_01090_),
    .A3(_01092_),
    .B1(_01094_),
    .Y(_02018_));
 sky130_fd_sc_hd__nor2_1 _08928_ (.A(_02017_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__xor2_4 _08929_ (.A(_02017_),
    .B(_02018_),
    .X(_02020_));
 sky130_fd_sc_hd__xnor2_4 _08930_ (.A(_02016_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__a21oi_4 _08931_ (.A1(_01102_),
    .A2(_01106_),
    .B1(_01105_),
    .Y(_02022_));
 sky130_fd_sc_hd__xnor2_2 _08932_ (.A(_02021_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__nand2b_1 _08933_ (.A_N(_02023_),
    .B(_02015_),
    .Y(_02024_));
 sky130_fd_sc_hd__xnor2_2 _08934_ (.A(_02015_),
    .B(_02023_),
    .Y(_02025_));
 sky130_fd_sc_hd__and2_1 _08935_ (.A(_02014_),
    .B(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__xor2_4 _08936_ (.A(_02014_),
    .B(_02025_),
    .X(_02027_));
 sky130_fd_sc_hd__xor2_4 _08937_ (.A(_02006_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__nor2_1 _08938_ (.A(_02005_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__xnor2_4 _08939_ (.A(_02005_),
    .B(_02028_),
    .Y(_02030_));
 sky130_fd_sc_hd__a21o_2 _08940_ (.A1(_02006_),
    .A2(_02027_),
    .B1(_02026_),
    .X(_02031_));
 sky130_fd_sc_hd__o21ai_4 _08941_ (.A1(_02021_),
    .A2(_02022_),
    .B1(_02024_),
    .Y(_02032_));
 sky130_fd_sc_hd__xor2_4 _08942_ (.A(_00765_),
    .B(_00767_),
    .X(_02033_));
 sky130_fd_sc_hd__o21ai_2 _08943_ (.A1(_02009_),
    .A2(_02010_),
    .B1(_02012_),
    .Y(_02034_));
 sky130_fd_sc_hd__xnor2_2 _08944_ (.A(_00759_),
    .B(_00760_),
    .Y(_02035_));
 sky130_fd_sc_hd__a21oi_2 _08945_ (.A1(_02016_),
    .A2(_02020_),
    .B1(_02019_),
    .Y(_02036_));
 sky130_fd_sc_hd__xnor2_2 _08946_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__nand2b_1 _08947_ (.A_N(_02037_),
    .B(_02034_),
    .Y(_02038_));
 sky130_fd_sc_hd__xnor2_2 _08948_ (.A(_02034_),
    .B(_02037_),
    .Y(_02039_));
 sky130_fd_sc_hd__and2_1 _08949_ (.A(_02033_),
    .B(_02039_),
    .X(_02040_));
 sky130_fd_sc_hd__xor2_4 _08950_ (.A(_02033_),
    .B(_02039_),
    .X(_02041_));
 sky130_fd_sc_hd__xor2_4 _08951_ (.A(_02032_),
    .B(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_02031_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__xor2_2 _08953_ (.A(_02031_),
    .B(_02042_),
    .X(_02044_));
 sky130_fd_sc_hd__xnor2_1 _08954_ (.A(_02031_),
    .B(_02042_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_1 _08955_ (.A(_02030_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__a21oi_2 _08956_ (.A1(_02032_),
    .A2(_02041_),
    .B1(_02040_),
    .Y(_02047_));
 sky130_fd_sc_hd__o21ai_2 _08957_ (.A1(_02035_),
    .A2(_02036_),
    .B1(_02038_),
    .Y(_02048_));
 sky130_fd_sc_hd__xor2_2 _08958_ (.A(_00489_),
    .B(_00490_),
    .X(_02049_));
 sky130_fd_sc_hd__xnor2_2 _08959_ (.A(_00768_),
    .B(_00769_),
    .Y(_02050_));
 sky130_fd_sc_hd__xnor2_2 _08960_ (.A(_02049_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__and2b_1 _08961_ (.A_N(_02051_),
    .B(_02048_),
    .X(_02052_));
 sky130_fd_sc_hd__xor2_2 _08962_ (.A(_02048_),
    .B(_02051_),
    .X(_02053_));
 sky130_fd_sc_hd__or2_1 _08963_ (.A(_02047_),
    .B(_02053_),
    .X(_02054_));
 sky130_fd_sc_hd__and2_1 _08964_ (.A(_02047_),
    .B(_02053_),
    .X(_02055_));
 sky130_fd_sc_hd__xor2_2 _08965_ (.A(_02047_),
    .B(_02053_),
    .X(_02056_));
 sky130_fd_sc_hd__inv_2 _08966_ (.A(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__a21o_2 _08967_ (.A1(_02049_),
    .A2(_02050_),
    .B1(_02052_),
    .X(_02058_));
 sky130_fd_sc_hd__xor2_4 _08968_ (.A(_00771_),
    .B(_00772_),
    .X(_02059_));
 sky130_fd_sc_hd__nor2_1 _08969_ (.A(_02058_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__xor2_2 _08970_ (.A(_02058_),
    .B(_02059_),
    .X(_02061_));
 sky130_fd_sc_hd__xnor2_2 _08971_ (.A(_02058_),
    .B(_02059_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand4_2 _08972_ (.A(_02004_),
    .B(_02046_),
    .C(_02056_),
    .D(_02061_),
    .Y(_02063_));
 sky130_fd_sc_hd__a21boi_1 _08973_ (.A1(_02058_),
    .A2(_02059_),
    .B1_N(_02054_),
    .Y(_02064_));
 sky130_fd_sc_hd__a22o_1 _08974_ (.A1(_02005_),
    .A2(_02028_),
    .B1(_02031_),
    .B2(_02042_),
    .X(_02065_));
 sky130_fd_sc_hd__o21ai_1 _08975_ (.A1(_02031_),
    .A2(_02042_),
    .B1(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__o32a_1 _08976_ (.A1(_02057_),
    .A2(_02062_),
    .A3(_02066_),
    .B1(_02064_),
    .B2(_02060_),
    .X(_02067_));
 sky130_fd_sc_hd__nand2_1 _08977_ (.A(_02063_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__xor2_2 _08978_ (.A(_00776_),
    .B(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__and2_2 _08979_ (.A(net309),
    .B(_04698_),
    .X(_02070_));
 sky130_fd_sc_hd__nand2_2 _08980_ (.A(net309),
    .B(_04698_),
    .Y(_02071_));
 sky130_fd_sc_hd__o31a_1 _08981_ (.A1(net213),
    .A2(_01767_),
    .A3(_01768_),
    .B1(_01773_),
    .X(_02072_));
 sky130_fd_sc_hd__xnor2_1 _08982_ (.A(_01776_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__or2_1 _08983_ (.A(_01769_),
    .B(_01772_),
    .X(_02074_));
 sky130_fd_sc_hd__and2_1 _08984_ (.A(_01773_),
    .B(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__nor2_1 _08985_ (.A(_01771_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _08986_ (.A(_02073_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__xnor2_1 _08987_ (.A(_01761_),
    .B(_01778_),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _08988_ (.A(_02077_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _08989_ (.A(_01779_),
    .B(_01781_),
    .Y(_02080_));
 sky130_fd_sc_hd__and2_1 _08990_ (.A(_02079_),
    .B(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__xnor2_1 _08991_ (.A(_01744_),
    .B(_01782_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _08992_ (.A(_02081_),
    .B(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__xnor2_1 _08993_ (.A(_01785_),
    .B(_01786_),
    .Y(_02084_));
 sky130_fd_sc_hd__or2_1 _08994_ (.A(_02083_),
    .B(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__xor2_2 _08995_ (.A(_01716_),
    .B(_01787_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_1 _08996_ (.A(_02085_),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__a21oi_1 _08997_ (.A1(_01702_),
    .A2(_01713_),
    .B1(_01787_),
    .Y(_02088_));
 sky130_fd_sc_hd__o211a_1 _08998_ (.A1(_01714_),
    .A2(_02088_),
    .B1(_01788_),
    .C1(_01701_),
    .X(_02089_));
 sky130_fd_sc_hd__a211oi_1 _08999_ (.A1(_01701_),
    .A2(_01788_),
    .B1(_02088_),
    .C1(_01714_),
    .Y(_02090_));
 sky130_fd_sc_hd__or2_1 _09000_ (.A(_02089_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__and2_1 _09001_ (.A(_02087_),
    .B(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__xor2_2 _09002_ (.A(_01681_),
    .B(_01790_),
    .X(_02093_));
 sky130_fd_sc_hd__and2_1 _09003_ (.A(_02092_),
    .B(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(_01679_),
    .B(_01788_),
    .Y(_02095_));
 sky130_fd_sc_hd__o21a_1 _09005_ (.A1(_02089_),
    .A2(_02095_),
    .B1(_01680_),
    .X(_02096_));
 sky130_fd_sc_hd__xnor2_1 _09006_ (.A(_01794_),
    .B(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__and3_1 _09007_ (.A(_02092_),
    .B(_02093_),
    .C(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__xnor2_1 _09008_ (.A(_01635_),
    .B(_01795_),
    .Y(_02099_));
 sky130_fd_sc_hd__and4_1 _09009_ (.A(_02092_),
    .B(_02093_),
    .C(_02097_),
    .D(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__xnor2_1 _09010_ (.A(_01604_),
    .B(_01605_),
    .Y(_02101_));
 sky130_fd_sc_hd__o21a_1 _09011_ (.A1(_01633_),
    .A2(_01791_),
    .B1(_01634_),
    .X(_02102_));
 sky130_fd_sc_hd__o2111a_1 _09012_ (.A1(_02089_),
    .A2(_02095_),
    .B1(_01635_),
    .C1(_01680_),
    .D1(_01794_),
    .X(_02103_));
 sky130_fd_sc_hd__nor2_1 _09013_ (.A(_02102_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__o21bai_1 _09014_ (.A1(_02102_),
    .A2(_02103_),
    .B1_N(_02101_),
    .Y(_02105_));
 sky130_fd_sc_hd__xnor2_1 _09015_ (.A(_02101_),
    .B(_02104_),
    .Y(_02106_));
 sky130_fd_sc_hd__and2_1 _09016_ (.A(_02100_),
    .B(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__xnor2_1 _09017_ (.A(_01582_),
    .B(_01798_),
    .Y(_02108_));
 sky130_fd_sc_hd__nor2_1 _09018_ (.A(_01579_),
    .B(_01796_),
    .Y(_02109_));
 sky130_fd_sc_hd__a21o_1 _09019_ (.A1(_02105_),
    .A2(_02109_),
    .B1(_01580_),
    .X(_02110_));
 sky130_fd_sc_hd__a211o_1 _09020_ (.A1(_02105_),
    .A2(_02109_),
    .B1(_01580_),
    .C1(_01801_),
    .X(_02111_));
 sky130_fd_sc_hd__xnor2_1 _09021_ (.A(_01801_),
    .B(_02110_),
    .Y(_02112_));
 sky130_fd_sc_hd__and3_1 _09022_ (.A(_02107_),
    .B(_02108_),
    .C(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__xnor2_1 _09023_ (.A(_01517_),
    .B(_01802_),
    .Y(_02114_));
 sky130_fd_sc_hd__o21ba_1 _09024_ (.A1(_01514_),
    .A2(_01515_),
    .B1_N(_01799_),
    .X(_02115_));
 sky130_fd_sc_hd__a22o_1 _09025_ (.A1(_01514_),
    .A2(_01515_),
    .B1(_02111_),
    .B2(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__xnor2_1 _09026_ (.A(_01806_),
    .B(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__and3_1 _09027_ (.A(_02113_),
    .B(_02114_),
    .C(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__xnor2_1 _09028_ (.A(_01435_),
    .B(_01807_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _09029_ (.A(_02118_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21o_1 _09030_ (.A1(_01432_),
    .A2(_01803_),
    .B1(_01433_),
    .X(_02121_));
 sky130_fd_sc_hd__o31a_1 _09031_ (.A1(_01434_),
    .A2(_01806_),
    .A3(_02116_),
    .B1(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__xnor2_2 _09032_ (.A(_01810_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__xnor2_1 _09033_ (.A(_01811_),
    .B(_01879_),
    .Y(_02124_));
 sky130_fd_sc_hd__and4b_1 _09034_ (.A_N(_02123_),
    .B(_02118_),
    .C(_02119_),
    .D(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__a21o_1 _09035_ (.A1(_01808_),
    .A2(_01877_),
    .B1(_01878_),
    .X(_02126_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(_01810_),
    .B(_01879_),
    .Y(_02127_));
 sky130_fd_sc_hd__o21ai_1 _09037_ (.A1(_02122_),
    .A2(_02127_),
    .B1(_02126_),
    .Y(_02128_));
 sky130_fd_sc_hd__xor2_2 _09038_ (.A(_01929_),
    .B(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nand2b_1 _09039_ (.A_N(_02129_),
    .B(_02125_),
    .Y(_02130_));
 sky130_fd_sc_hd__xnor2_2 _09040_ (.A(_01932_),
    .B(_01960_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21o_1 _09041_ (.A1(_01927_),
    .A2(_01958_),
    .B1(_01959_),
    .X(_02132_));
 sky130_fd_sc_hd__nand2_1 _09042_ (.A(_01929_),
    .B(_01960_),
    .Y(_02133_));
 sky130_fd_sc_hd__or4bb_1 _09043_ (.A(_02126_),
    .B(_01928_),
    .C_N(_01927_),
    .D_N(_01960_),
    .X(_02134_));
 sky130_fd_sc_hd__o311a_1 _09044_ (.A1(_02122_),
    .A2(_02127_),
    .A3(_02133_),
    .B1(_02134_),
    .C1(_02132_),
    .X(_02135_));
 sky130_fd_sc_hd__xor2_1 _09045_ (.A(_01976_),
    .B(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__and4bb_2 _09046_ (.A_N(_02129_),
    .B_N(_02131_),
    .C(_02136_),
    .D(_02125_),
    .X(_02137_));
 sky130_fd_sc_hd__xor2_2 _09047_ (.A(_01990_),
    .B(_01998_),
    .X(_02138_));
 sky130_fd_sc_hd__a21o_1 _09048_ (.A1(_01975_),
    .A2(_01988_),
    .B1(_01989_),
    .X(_02139_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(_01976_),
    .B(_01990_),
    .Y(_02140_));
 sky130_fd_sc_hd__o21a_1 _09050_ (.A1(_02135_),
    .A2(_02140_),
    .B1(_02139_),
    .X(_02141_));
 sky130_fd_sc_hd__xnor2_1 _09051_ (.A(_01994_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand3b_2 _09052_ (.A_N(_02142_),
    .B(_02137_),
    .C(_02138_),
    .Y(_02143_));
 sky130_fd_sc_hd__xor2_2 _09053_ (.A(_01999_),
    .B(_02001_),
    .X(_02144_));
 sky130_fd_sc_hd__a21boi_1 _09054_ (.A1(_01175_),
    .A2(_01993_),
    .B1_N(_02000_),
    .Y(_02145_));
 sky130_fd_sc_hd__inv_2 _09055_ (.A(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_1 _09056_ (.A(_01994_),
    .B(_02001_),
    .Y(_02147_));
 sky130_fd_sc_hd__o21a_1 _09057_ (.A1(_02141_),
    .A2(_02147_),
    .B1(_02146_),
    .X(_02148_));
 sky130_fd_sc_hd__xnor2_1 _09058_ (.A(_02002_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__or3_2 _09059_ (.A(_02143_),
    .B(_02144_),
    .C(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__xnor2_2 _09060_ (.A(_02004_),
    .B(_02030_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_2 _09061_ (.A(_02150_),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__a22oi_1 _09062_ (.A1(_01071_),
    .A2(_01113_),
    .B1(_02005_),
    .B2(_02028_),
    .Y(_02153_));
 sky130_fd_sc_hd__or2_1 _09063_ (.A(_02003_),
    .B(_02030_),
    .X(_02154_));
 sky130_fd_sc_hd__o32a_1 _09064_ (.A1(_02003_),
    .A2(_02030_),
    .A3(_02146_),
    .B1(_02153_),
    .B2(_02029_),
    .X(_02155_));
 sky130_fd_sc_hd__or4_1 _09065_ (.A(_02003_),
    .B(_02030_),
    .C(_02141_),
    .D(_02147_),
    .X(_02156_));
 sky130_fd_sc_hd__nand2_1 _09066_ (.A(_02155_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_2 _09067_ (.A(_02044_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21boi_2 _09068_ (.A1(_02004_),
    .A2(_02046_),
    .B1_N(_02066_),
    .Y(_02159_));
 sky130_fd_sc_hd__xnor2_2 _09069_ (.A(_02057_),
    .B(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hd__and3_1 _09070_ (.A(_02152_),
    .B(_02158_),
    .C(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__a21o_1 _09071_ (.A1(_02043_),
    .A2(_02054_),
    .B1(_02055_),
    .X(_02162_));
 sky130_fd_sc_hd__nand2_1 _09072_ (.A(_02044_),
    .B(_02056_),
    .Y(_02163_));
 sky130_fd_sc_hd__or4b_2 _09073_ (.A(_02029_),
    .B(_02045_),
    .C(_02153_),
    .D_N(_02056_),
    .X(_02164_));
 sky130_fd_sc_hd__o311ai_4 _09074_ (.A1(_02148_),
    .A2(_02154_),
    .A3(_02163_),
    .B1(_02164_),
    .C1(_02162_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_2 _09075_ (.A(_02061_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__and2_1 _09076_ (.A(_02161_),
    .B(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__nand4_2 _09077_ (.A(_02152_),
    .B(_02158_),
    .C(_02160_),
    .D(_02166_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _09078_ (.A(net161),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__nand2_1 _09079_ (.A(_02069_),
    .B(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_4 _09080_ (.A(_06422_),
    .B(_06428_),
    .Y(_02171_));
 sky130_fd_sc_hd__or2_1 _09081_ (.A(_06422_),
    .B(_06428_),
    .X(_02172_));
 sky130_fd_sc_hd__o211a_1 _09082_ (.A1(_02069_),
    .A2(_02169_),
    .B1(_02170_),
    .C1(_02171_),
    .X(_02173_));
 sky130_fd_sc_hd__nor2_1 _09083_ (.A(net304),
    .B(_06451_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand2_4 _09084_ (.A(net309),
    .B(_06450_),
    .Y(_02175_));
 sky130_fd_sc_hd__mux2_1 _09085_ (.A0(reg1_val[1]),
    .A1(reg1_val[30]),
    .S(net191),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(net308),
    .A1(reg1_val[31]),
    .S(net191),
    .X(_02177_));
 sky130_fd_sc_hd__mux2_1 _09087_ (.A0(_02176_),
    .A1(_02177_),
    .S(net228),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _09088_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net191),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net191),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_1 _09090_ (.A0(_02179_),
    .A1(_02180_),
    .S(net228),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_1 _09091_ (.A0(_02178_),
    .A1(_02181_),
    .S(net230),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_1 _09092_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net191),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _09093_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net191),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _09094_ (.A0(_02183_),
    .A1(_02184_),
    .S(net227),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _09095_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net191),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _09096_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net191),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(_02186_),
    .A1(_02187_),
    .S(net227),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _09098_ (.A0(_02185_),
    .A1(_02188_),
    .S(net231),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _09099_ (.A0(_02182_),
    .A1(_02189_),
    .S(net234),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _09100_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(net191),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _09101_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(net191),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _09102_ (.A0(_02191_),
    .A1(_02192_),
    .S(net227),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _09103_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net191),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net191),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _09105_ (.A0(_02194_),
    .A1(_02195_),
    .S(net227),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _09106_ (.A0(_02193_),
    .A1(_02196_),
    .S(net231),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _09107_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net191),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _09108_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net191),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _09109_ (.A0(_02198_),
    .A1(_02199_),
    .S(net227),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _09110_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net192),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _09111_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net192),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _09112_ (.A0(_02201_),
    .A1(_02202_),
    .S(net227),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _09113_ (.A0(_02200_),
    .A1(_02203_),
    .S(net231),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _09114_ (.A0(_02197_),
    .A1(_02204_),
    .S(net235),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _09115_ (.A0(_02190_),
    .A1(_02205_),
    .S(net237),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net189),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _09117_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net189),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(_02207_),
    .A1(_02208_),
    .S(net227),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net189),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net189),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _09121_ (.A0(_02210_),
    .A1(_02211_),
    .S(net227),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(_02209_),
    .A1(_02212_),
    .S(net231),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _09123_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net189),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net189),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _09125_ (.A0(_02214_),
    .A1(_02215_),
    .S(net227),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _09126_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(_02175_),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(_02175_),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _09128_ (.A0(_02217_),
    .A1(_02218_),
    .S(net227),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _09129_ (.A0(_02216_),
    .A1(_02219_),
    .S(net232),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(_02213_),
    .A1(_02220_),
    .S(net235),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _09131_ (.A0(reg1_val[0]),
    .A1(reg1_val[31]),
    .S(net189),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(net307),
    .A1(reg1_val[30]),
    .S(net189),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _09133_ (.A0(_02222_),
    .A1(_02223_),
    .S(net228),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net189),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _09135_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net189),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(_02225_),
    .A1(_02226_),
    .S(net228),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _09137_ (.A0(_02224_),
    .A1(_02227_),
    .S(net231),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _09138_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net189),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _09139_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net189),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(_02229_),
    .A1(_02230_),
    .S(net228),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _09141_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net189),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _09142_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net189),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(_02232_),
    .A1(_02233_),
    .S(net228),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _09144_ (.A0(_02231_),
    .A1(_02234_),
    .S(net231),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _09145_ (.A0(_02228_),
    .A1(_02235_),
    .S(net235),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(_02221_),
    .A1(_02236_),
    .S(net237),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(_02206_),
    .A1(_02237_),
    .S(net242),
    .X(_02238_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(net308),
    .B(curr_PC[0]),
    .Y(_02239_));
 sky130_fd_sc_hd__or2_1 _09149_ (.A(net308),
    .B(curr_PC[0]),
    .X(_02240_));
 sky130_fd_sc_hd__a21o_1 _09150_ (.A1(_02239_),
    .A2(_02240_),
    .B1(net243),
    .X(_02241_));
 sky130_fd_sc_hd__o211a_1 _09151_ (.A1(net269),
    .A2(_02238_),
    .B1(_02241_),
    .C1(_06446_),
    .X(_02242_));
 sky130_fd_sc_hd__nor2_4 _09152_ (.A(net309),
    .B(_06451_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_1 _09153_ (.A(net303),
    .B(_06450_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_4 _09154_ (.A(_06449_),
    .B(_06457_),
    .Y(_02245_));
 sky130_fd_sc_hd__or2_1 _09155_ (.A(_06449_),
    .B(_06457_),
    .X(_02246_));
 sky130_fd_sc_hd__nor2_8 _09156_ (.A(_06407_),
    .B(_06448_),
    .Y(_02247_));
 sky130_fd_sc_hd__or2_1 _09157_ (.A(_06407_),
    .B(_06448_),
    .X(_02248_));
 sky130_fd_sc_hd__nor2_2 _09158_ (.A(_06420_),
    .B(_06457_),
    .Y(_02249_));
 sky130_fd_sc_hd__or2_1 _09159_ (.A(_06420_),
    .B(_06457_),
    .X(_02250_));
 sky130_fd_sc_hd__a21o_1 _09160_ (.A1(net255),
    .A2(net254),
    .B1(_06408_),
    .X(_02251_));
 sky130_fd_sc_hd__a21oi_1 _09161_ (.A1(net208),
    .A2(_02251_),
    .B1(_06409_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_2 _09162_ (.A(_06407_),
    .B(_06428_),
    .Y(_02253_));
 sky130_fd_sc_hd__or2_4 _09163_ (.A(_06407_),
    .B(_06428_),
    .X(_02254_));
 sky130_fd_sc_hd__and4bb_4 _09164_ (.A_N(instruction[4]),
    .B_N(instruction[6]),
    .C(instruction[5]),
    .D(instruction[3]),
    .X(_02255_));
 sky130_fd_sc_hd__or3b_2 _09165_ (.A(_06422_),
    .B(instruction[6]),
    .C_N(instruction[5]),
    .X(_02256_));
 sky130_fd_sc_hd__o21a_1 _09166_ (.A1(_02253_),
    .A2(_02255_),
    .B1(_06408_),
    .X(_02257_));
 sky130_fd_sc_hd__nor2_2 _09167_ (.A(_06420_),
    .B(_06428_),
    .Y(_02258_));
 sky130_fd_sc_hd__or2_1 _09168_ (.A(_06420_),
    .B(_06428_),
    .X(_02259_));
 sky130_fd_sc_hd__nor2_2 _09169_ (.A(_06428_),
    .B(_06449_),
    .Y(_02260_));
 sky130_fd_sc_hd__or2_1 _09170_ (.A(_06428_),
    .B(_06449_),
    .X(_02261_));
 sky130_fd_sc_hd__a221o_1 _09171_ (.A1(\div_shifter[32] ),
    .A2(_02258_),
    .B1(_02260_),
    .B2(\div_res[0] ),
    .C1(_02257_),
    .X(_02262_));
 sky130_fd_sc_hd__and2_2 _09172_ (.A(reg1_val[31]),
    .B(net216),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _09173_ (.A0(_02222_),
    .A1(_02263_),
    .S(net224),
    .X(_02264_));
 sky130_fd_sc_hd__o21a_1 _09174_ (.A1(net232),
    .A2(_02263_),
    .B1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__or2_2 _09175_ (.A(net235),
    .B(_02263_),
    .X(_02266_));
 sky130_fd_sc_hd__and2_1 _09176_ (.A(_02265_),
    .B(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__nor2_1 _09177_ (.A(net238),
    .B(_02263_),
    .Y(_02268_));
 sky130_fd_sc_hd__or2_2 _09178_ (.A(net238),
    .B(_02263_),
    .X(_02269_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(_02267_),
    .B(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _09180_ (.A(net239),
    .B(_02263_),
    .Y(_02271_));
 sky130_fd_sc_hd__or2_4 _09181_ (.A(net239),
    .B(_02263_),
    .X(_02272_));
 sky130_fd_sc_hd__nor2_2 _09182_ (.A(_02270_),
    .B(_02271_),
    .Y(_02273_));
 sky130_fd_sc_hd__a211o_1 _09183_ (.A1(net191),
    .A2(_02273_),
    .B1(_02262_),
    .C1(_02252_),
    .X(_02274_));
 sky130_fd_sc_hd__a211o_1 _09184_ (.A1(_02238_),
    .A2(_02243_),
    .B1(_02274_),
    .C1(_02242_),
    .X(_02275_));
 sky130_fd_sc_hd__a211oi_1 _09185_ (.A1(_06405_),
    .A2(_06458_),
    .B1(_02173_),
    .C1(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__o31a_1 _09186_ (.A1(instruction[5]),
    .A2(_06397_),
    .A3(_06420_),
    .B1(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(net226),
    .A1(_02277_),
    .S(net215),
    .X(_02278_));
 sky130_fd_sc_hd__or2_1 _09188_ (.A(curr_PC[0]),
    .B(net262),
    .X(_02279_));
 sky130_fd_sc_hd__o21ai_4 _09189_ (.A1(net267),
    .A2(_02278_),
    .B1(_02279_),
    .Y(dest_val[0]));
 sky130_fd_sc_hd__a31o_1 _09190_ (.A1(_02069_),
    .A2(_02161_),
    .A3(_02166_),
    .B1(net158),
    .X(_02280_));
 sky130_fd_sc_hd__a21oi_4 _09191_ (.A1(_00494_),
    .A2(_00688_),
    .B1(_00687_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_4 _09192_ (.A(_00683_),
    .B(_00685_),
    .Y(_02282_));
 sky130_fd_sc_hd__a32o_2 _09193_ (.A1(_00581_),
    .A2(_00582_),
    .A3(_00591_),
    .B1(_00592_),
    .B2(_00572_),
    .X(_02283_));
 sky130_fd_sc_hd__o22a_1 _09194_ (.A1(net144),
    .A2(net16),
    .B1(net37),
    .B2(net148),
    .X(_02284_));
 sky130_fd_sc_hd__xnor2_1 _09195_ (.A(net78),
    .B(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__o22a_1 _09196_ (.A1(net23),
    .A2(net140),
    .B1(_00186_),
    .B2(net71),
    .X(_02286_));
 sky130_fd_sc_hd__xor2_1 _09197_ (.A(net110),
    .B(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__or2_1 _09198_ (.A(_02285_),
    .B(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(_02285_),
    .B(_02287_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _09200_ (.A(_02288_),
    .B(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__o22a_1 _09201_ (.A1(net30),
    .A2(net146),
    .B1(net142),
    .B2(net28),
    .X(_02291_));
 sky130_fd_sc_hd__xnor2_1 _09202_ (.A(_06524_),
    .B(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__xnor2_1 _09203_ (.A(_02290_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__a21oi_1 _09204_ (.A1(_00558_),
    .A2(_00560_),
    .B1(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__and3_1 _09205_ (.A(_00558_),
    .B(_00560_),
    .C(_02293_),
    .X(_02295_));
 sky130_fd_sc_hd__or2_2 _09206_ (.A(_02294_),
    .B(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__and2b_1 _09207_ (.A_N(_02296_),
    .B(_02283_),
    .X(_02297_));
 sky130_fd_sc_hd__xnor2_4 _09208_ (.A(_02283_),
    .B(_02296_),
    .Y(_02298_));
 sky130_fd_sc_hd__nand2_2 _09209_ (.A(_00577_),
    .B(_00581_),
    .Y(_02299_));
 sky130_fd_sc_hd__o21ba_1 _09210_ (.A1(_00568_),
    .A2(_00571_),
    .B1_N(_00567_),
    .X(_02300_));
 sky130_fd_sc_hd__o21ba_1 _09211_ (.A1(_00630_),
    .A2(_00635_),
    .B1_N(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__or3b_2 _09212_ (.A(_00630_),
    .B(_00635_),
    .C_N(_02300_),
    .X(_02302_));
 sky130_fd_sc_hd__and2b_1 _09213_ (.A_N(_02301_),
    .B(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__xnor2_2 _09214_ (.A(_02299_),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__o22a_1 _09215_ (.A1(net49),
    .A2(net88),
    .B1(net83),
    .B2(net46),
    .X(_02305_));
 sky130_fd_sc_hd__xnor2_1 _09216_ (.A(_06469_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__o22a_1 _09217_ (.A1(net63),
    .A2(net132),
    .B1(net170),
    .B2(net60),
    .X(_02307_));
 sky130_fd_sc_hd__xnor2_1 _09218_ (.A(net194),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2_1 _09219_ (.A(_02306_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__xor2_1 _09220_ (.A(_02306_),
    .B(_02308_),
    .X(_02310_));
 sky130_fd_sc_hd__o22a_1 _09221_ (.A1(net55),
    .A2(net130),
    .B1(net128),
    .B2(net52),
    .X(_02311_));
 sky130_fd_sc_hd__xnor2_1 _09222_ (.A(net167),
    .B(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__and2b_1 _09223_ (.A_N(_02312_),
    .B(_02310_),
    .X(_02313_));
 sky130_fd_sc_hd__and2b_1 _09224_ (.A_N(_02310_),
    .B(_02312_),
    .X(_02314_));
 sky130_fd_sc_hd__nor2_1 _09225_ (.A(_02313_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__o22a_1 _09226_ (.A1(net125),
    .A2(net43),
    .B1(net40),
    .B2(net121),
    .X(_02316_));
 sky130_fd_sc_hd__xor2_1 _09227_ (.A(net153),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__o22a_1 _09228_ (.A1(_06491_),
    .A2(net69),
    .B1(net95),
    .B2(_06494_),
    .X(_02318_));
 sky130_fd_sc_hd__xnor2_1 _09229_ (.A(net101),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_02317_),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__or2_1 _09231_ (.A(_02317_),
    .B(_02319_),
    .X(_02321_));
 sky130_fd_sc_hd__nand2_2 _09232_ (.A(_02320_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__o22a_1 _09233_ (.A1(net74),
    .A2(net86),
    .B1(net81),
    .B2(net115),
    .X(_02323_));
 sky130_fd_sc_hd__xnor2_2 _09234_ (.A(_06500_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__xor2_2 _09235_ (.A(_02322_),
    .B(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__o22a_1 _09236_ (.A1(net178),
    .A2(net14),
    .B1(net7),
    .B2(net175),
    .X(_02326_));
 sky130_fd_sc_hd__xnor2_1 _09237_ (.A(_00210_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__or2_1 _09238_ (.A(net57),
    .B(net134),
    .X(_02328_));
 sky130_fd_sc_hd__a21o_1 _09239_ (.A1(_00243_),
    .A2(_00244_),
    .B1(net172),
    .X(_02329_));
 sky130_fd_sc_hd__a21o_1 _09240_ (.A1(_02328_),
    .A2(_02329_),
    .B1(net211),
    .X(_02330_));
 sky130_fd_sc_hd__nand3_1 _09241_ (.A(net211),
    .B(_02328_),
    .C(_02329_),
    .Y(_02331_));
 sky130_fd_sc_hd__and3_1 _09242_ (.A(_00213_),
    .B(_02330_),
    .C(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__a21oi_1 _09243_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_00213_),
    .Y(_02333_));
 sky130_fd_sc_hd__a21o_1 _09244_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_00213_),
    .X(_02334_));
 sky130_fd_sc_hd__or3b_1 _09245_ (.A(_02332_),
    .B(_02333_),
    .C_N(_02327_),
    .X(_02335_));
 sky130_fd_sc_hd__o21bai_1 _09246_ (.A1(_02332_),
    .A2(_02333_),
    .B1_N(_02327_),
    .Y(_02336_));
 sky130_fd_sc_hd__nand3_2 _09247_ (.A(_02325_),
    .B(_02335_),
    .C(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__a21o_1 _09248_ (.A1(_02335_),
    .A2(_02336_),
    .B1(_02325_),
    .X(_02338_));
 sky130_fd_sc_hd__nand3_2 _09249_ (.A(_02315_),
    .B(_02337_),
    .C(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__a21o_1 _09250_ (.A1(_02337_),
    .A2(_02338_),
    .B1(_02315_),
    .X(_02340_));
 sky130_fd_sc_hd__nand2_1 _09251_ (.A(_06526_),
    .B(net35),
    .Y(_02341_));
 sky130_fd_sc_hd__a21o_1 _09252_ (.A1(_00585_),
    .A2(_00590_),
    .B1(_00589_),
    .X(_02342_));
 sky130_fd_sc_hd__o22a_1 _09253_ (.A1(net180),
    .A2(net11),
    .B1(net5),
    .B2(net183),
    .X(_02343_));
 sky130_fd_sc_hd__xnor2_1 _09254_ (.A(_00596_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__and2b_1 _09255_ (.A_N(_02344_),
    .B(_02342_),
    .X(_02345_));
 sky130_fd_sc_hd__xnor2_1 _09256_ (.A(_02342_),
    .B(_02344_),
    .Y(_02346_));
 sky130_fd_sc_hd__xnor2_1 _09257_ (.A(_02341_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__and3_1 _09258_ (.A(_02339_),
    .B(_02340_),
    .C(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__a21oi_2 _09259_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_02347_),
    .Y(_02349_));
 sky130_fd_sc_hd__or3_1 _09260_ (.A(_02304_),
    .B(_02348_),
    .C(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__o21ai_1 _09261_ (.A1(_02348_),
    .A2(_02349_),
    .B1(_02304_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(_02350_),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__o21ai_1 _09263_ (.A1(_00537_),
    .A2(_00539_),
    .B1(_00535_),
    .Y(_02353_));
 sky130_fd_sc_hd__or2_1 _09264_ (.A(net117),
    .B(net20),
    .X(_02354_));
 sky130_fd_sc_hd__or2_1 _09265_ (.A(net113),
    .B(net65),
    .X(_02355_));
 sky130_fd_sc_hd__and3_1 _09266_ (.A(net93),
    .B(_02354_),
    .C(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_1 _09267_ (.A1(_02354_),
    .A2(_02355_),
    .B1(net93),
    .Y(_02357_));
 sky130_fd_sc_hd__or2_1 _09268_ (.A(net25),
    .B(net135),
    .X(_02358_));
 sky130_fd_sc_hd__or2_1 _09269_ (.A(_06558_),
    .B(net98),
    .X(_02359_));
 sky130_fd_sc_hd__and3_1 _09270_ (.A(net107),
    .B(_02358_),
    .C(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__a21oi_1 _09271_ (.A1(_02358_),
    .A2(_02359_),
    .B1(net107),
    .Y(_02361_));
 sky130_fd_sc_hd__o22a_1 _09272_ (.A1(_02356_),
    .A2(_02357_),
    .B1(_02360_),
    .B2(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__or4_1 _09273_ (.A(_02356_),
    .B(_02357_),
    .C(_02360_),
    .D(_02361_),
    .X(_02363_));
 sky130_fd_sc_hd__and2b_1 _09274_ (.A_N(_02362_),
    .B(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__o22a_1 _09275_ (.A1(_00166_),
    .A2(net22),
    .B1(net67),
    .B2(net90),
    .X(_02365_));
 sky130_fd_sc_hd__xnor2_2 _09276_ (.A(net103),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__xor2_2 _09277_ (.A(_02364_),
    .B(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__a31o_1 _09278_ (.A1(net224),
    .A2(net35),
    .A3(_00605_),
    .B1(_00604_),
    .X(_02368_));
 sky130_fd_sc_hd__nand2_1 _09279_ (.A(_02367_),
    .B(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__xor2_1 _09280_ (.A(_02367_),
    .B(_02368_),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_1 _09281_ (.A(_02353_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _09282_ (.A(_02352_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(_02352_),
    .B(_02371_),
    .Y(_02373_));
 sky130_fd_sc_hd__and2b_1 _09284_ (.A_N(_02372_),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__xor2_4 _09285_ (.A(_02298_),
    .B(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__a21o_2 _09286_ (.A1(_00550_),
    .A2(_00649_),
    .B1(_00648_),
    .X(_02376_));
 sky130_fd_sc_hd__nand2_4 _09287_ (.A(_00546_),
    .B(_00549_),
    .Y(_02377_));
 sky130_fd_sc_hd__a21bo_1 _09288_ (.A1(_00562_),
    .A2(_00608_),
    .B1_N(_00607_),
    .X(_02378_));
 sky130_fd_sc_hd__a21oi_4 _09289_ (.A1(_00621_),
    .A2(_00646_),
    .B1(_00645_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_1 _09290_ (.A1(_00607_),
    .A2(_00609_),
    .B1(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__xnor2_4 _09291_ (.A(_02378_),
    .B(_02379_),
    .Y(_02381_));
 sky130_fd_sc_hd__xnor2_4 _09292_ (.A(_02377_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__a21oi_4 _09293_ (.A1(_00676_),
    .A2(_00680_),
    .B1(_00679_),
    .Y(_02383_));
 sky130_fd_sc_hd__xnor2_4 _09294_ (.A(_02382_),
    .B(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2b_1 _09295_ (.A_N(_02384_),
    .B(_02376_),
    .Y(_02385_));
 sky130_fd_sc_hd__xnor2_4 _09296_ (.A(_02376_),
    .B(_02384_),
    .Y(_02386_));
 sky130_fd_sc_hd__and2_1 _09297_ (.A(_02375_),
    .B(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__xor2_4 _09298_ (.A(_02375_),
    .B(_02386_),
    .X(_02388_));
 sky130_fd_sc_hd__xnor2_4 _09299_ (.A(_02282_),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__or2_1 _09300_ (.A(_02281_),
    .B(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__and2_1 _09301_ (.A(_02281_),
    .B(_02389_),
    .X(_02391_));
 sky130_fd_sc_hd__xnor2_4 _09302_ (.A(_02281_),
    .B(_02389_),
    .Y(_02392_));
 sky130_fd_sc_hd__o2bb2a_1 _09303_ (.A1_N(_02058_),
    .A2_N(_02059_),
    .B1(_00689_),
    .B2(_00773_),
    .X(_02393_));
 sky130_fd_sc_hd__nor2_1 _09304_ (.A(_00775_),
    .B(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__o32a_1 _09305_ (.A1(_00776_),
    .A2(_02062_),
    .A3(_02162_),
    .B1(_02393_),
    .B2(_00775_),
    .X(_02395_));
 sky130_fd_sc_hd__a2111o_1 _09306_ (.A1(_02155_),
    .A2(_02156_),
    .B1(_02163_),
    .C1(_02062_),
    .D1(_00776_),
    .X(_02396_));
 sky130_fd_sc_hd__and2_1 _09307_ (.A(_02395_),
    .B(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__xnor2_2 _09308_ (.A(_02392_),
    .B(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__a21oi_1 _09309_ (.A1(_02280_),
    .A2(_02398_),
    .B1(net209),
    .Y(_02399_));
 sky130_fd_sc_hd__o21ai_1 _09310_ (.A1(_02280_),
    .A2(_02398_),
    .B1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(_02176_),
    .A1(_02180_),
    .S(_06351_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _09312_ (.A0(_02179_),
    .A1(_02187_),
    .S(net224),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(_02401_),
    .A1(_02402_),
    .S(net230),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(_02183_),
    .A1(_02202_),
    .S(net224),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(_02184_),
    .A1(_02186_),
    .S(net227),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(_02404_),
    .A1(_02405_),
    .S(net231),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(_02403_),
    .A1(_02406_),
    .S(net234),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(_02191_),
    .A1(_02218_),
    .S(net224),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(_02192_),
    .A1(_02194_),
    .S(net227),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(_02408_),
    .A1(_02409_),
    .S(net231),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(_02195_),
    .A1(_02198_),
    .S(net227),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _09322_ (.A0(_02199_),
    .A1(_02201_),
    .S(net228),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(_02411_),
    .A1(_02412_),
    .S(net231),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(_02410_),
    .A1(_02413_),
    .S(_06337_),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(_02407_),
    .A1(_02414_),
    .S(net237),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _09326_ (.A0(_02207_),
    .A1(_02233_),
    .S(net224),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(_02208_),
    .A1(_02210_),
    .S(net227),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _09328_ (.A0(_02416_),
    .A1(_02417_),
    .S(net232),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(_02211_),
    .A1(_02214_),
    .S(net227),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(_02215_),
    .A1(_02217_),
    .S(net227),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(_02419_),
    .A1(_02420_),
    .S(net232),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _09332_ (.A0(_02418_),
    .A1(_02421_),
    .S(net235),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _09333_ (.A0(_02223_),
    .A1(_02225_),
    .S(net228),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _09334_ (.A0(_02264_),
    .A1(_02423_),
    .S(net232),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(_02226_),
    .A1(_02229_),
    .S(net228),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _09336_ (.A0(_02230_),
    .A1(_02232_),
    .S(net228),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(_02425_),
    .A1(_02426_),
    .S(net231),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _09338_ (.A0(_02424_),
    .A1(_02427_),
    .S(net235),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(_02422_),
    .A1(_02428_),
    .S(net236),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _09340_ (.A0(_02415_),
    .A1(_02429_),
    .S(net240),
    .X(_02430_));
 sky130_fd_sc_hd__inv_2 _09341_ (.A(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__nand2_1 _09342_ (.A(net307),
    .B(curr_PC[1]),
    .Y(_02432_));
 sky130_fd_sc_hd__or2_1 _09343_ (.A(net307),
    .B(curr_PC[1]),
    .X(_02433_));
 sky130_fd_sc_hd__nand2_1 _09344_ (.A(_02432_),
    .B(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__xnor2_1 _09345_ (.A(_02239_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__a21o_1 _09346_ (.A1(net268),
    .A2(_02435_),
    .B1(_06447_),
    .X(_02436_));
 sky130_fd_sc_hd__a21oi_1 _09347_ (.A1(net188),
    .A2(_02436_),
    .B1(_02431_),
    .Y(_02437_));
 sky130_fd_sc_hd__a21oi_1 _09348_ (.A1(\div_res[0] ),
    .A2(net165),
    .B1(\div_res[1] ),
    .Y(_02438_));
 sky130_fd_sc_hd__a311o_1 _09349_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .A3(net165),
    .B1(net205),
    .C1(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__xnor2_1 _09350_ (.A(_06348_),
    .B(_06352_),
    .Y(_02440_));
 sky130_fd_sc_hd__nand2_1 _09351_ (.A(net304),
    .B(net224),
    .Y(_02441_));
 sky130_fd_sc_hd__a21oi_1 _09352_ (.A1(_02440_),
    .A2(_02441_),
    .B1(net255),
    .Y(_02442_));
 sky130_fd_sc_hd__o21ai_1 _09353_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__or3b_1 _09354_ (.A(net231),
    .B(net206),
    .C_N(net307),
    .X(_02444_));
 sky130_fd_sc_hd__and2_1 _09355_ (.A(divi1_sign),
    .B(net310),
    .X(_02445_));
 sky130_fd_sc_hd__and3_1 _09356_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .C(net247),
    .X(_02446_));
 sky130_fd_sc_hd__a21oi_1 _09357_ (.A1(\div_shifter[32] ),
    .A2(net247),
    .B1(\div_shifter[33] ),
    .Y(_02447_));
 sky130_fd_sc_hd__o32a_1 _09358_ (.A1(net250),
    .A2(_02446_),
    .A3(_02447_),
    .B1(_06460_),
    .B2(net231),
    .X(_02448_));
 sky130_fd_sc_hd__o2bb2a_1 _09359_ (.A1_N(_06347_),
    .A2_N(_02245_),
    .B1(_02436_),
    .B2(net244),
    .X(_02449_));
 sky130_fd_sc_hd__o2111a_1 _09360_ (.A1(_06348_),
    .A2(net254),
    .B1(_02444_),
    .C1(_02448_),
    .D1(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__and4b_1 _09361_ (.A_N(_02437_),
    .B(_02439_),
    .C(_02443_),
    .D(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__o21ai_1 _09362_ (.A1(net260),
    .A2(net158),
    .B1(_06408_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21oi_1 _09363_ (.A1(net260),
    .A2(net158),
    .B1(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_1 _09364_ (.A(_01770_),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__mux2_1 _09365_ (.A0(_02224_),
    .A1(_02263_),
    .S(net230),
    .X(_02455_));
 sky130_fd_sc_hd__o21ai_2 _09366_ (.A1(net233),
    .A2(_02455_),
    .B1(_02266_),
    .Y(_02456_));
 sky130_fd_sc_hd__inv_2 _09367_ (.A(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__a21oi_2 _09368_ (.A1(net238),
    .A2(_02456_),
    .B1(_02268_),
    .Y(_02458_));
 sky130_fd_sc_hd__o21ai_2 _09369_ (.A1(net240),
    .A2(_02458_),
    .B1(_02272_),
    .Y(_02459_));
 sky130_fd_sc_hd__o22a_1 _09370_ (.A1(_02254_),
    .A2(_02454_),
    .B1(_02459_),
    .B2(net189),
    .X(_02460_));
 sky130_fd_sc_hd__and3_1 _09371_ (.A(_02400_),
    .B(_02451_),
    .C(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(net267),
    .B(_02461_),
    .Y(_02462_));
 sky130_fd_sc_hd__or2_1 _09373_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .X(_02463_));
 sky130_fd_sc_hd__nand2_1 _09374_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .Y(_02464_));
 sky130_fd_sc_hd__a31o_4 _09375_ (.A1(net267),
    .A2(_02463_),
    .A3(_02464_),
    .B1(_02462_),
    .X(dest_val[1]));
 sky130_fd_sc_hd__a31o_1 _09376_ (.A1(_02069_),
    .A2(_02167_),
    .A3(_02398_),
    .B1(net158),
    .X(_02465_));
 sky130_fd_sc_hd__a21oi_4 _09377_ (.A1(_02282_),
    .A2(_02388_),
    .B1(_02387_),
    .Y(_02466_));
 sky130_fd_sc_hd__o21ai_4 _09378_ (.A1(_02382_),
    .A2(_02383_),
    .B1(_02385_),
    .Y(_02467_));
 sky130_fd_sc_hd__nand2_2 _09379_ (.A(_02337_),
    .B(_02339_),
    .Y(_02468_));
 sky130_fd_sc_hd__o22a_1 _09380_ (.A1(net148),
    .A2(net16),
    .B1(net37),
    .B2(net146),
    .X(_02469_));
 sky130_fd_sc_hd__xnor2_1 _09381_ (.A(net78),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__o22a_1 _09382_ (.A1(net23),
    .A2(_00186_),
    .B1(_00191_),
    .B2(net71),
    .X(_02471_));
 sky130_fd_sc_hd__xor2_1 _09383_ (.A(net110),
    .B(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__or2_1 _09384_ (.A(_02470_),
    .B(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(_02470_),
    .B(_02472_),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_2 _09386_ (.A(_02473_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__o22a_2 _09387_ (.A1(net30),
    .A2(net142),
    .B1(_00180_),
    .B2(net28),
    .X(_02476_));
 sky130_fd_sc_hd__xnor2_4 _09388_ (.A(_06524_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__xnor2_4 _09389_ (.A(_02475_),
    .B(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__a21oi_4 _09390_ (.A1(_02299_),
    .A2(_02302_),
    .B1(_02301_),
    .Y(_02479_));
 sky130_fd_sc_hd__xnor2_4 _09391_ (.A(_02478_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__nand2b_1 _09392_ (.A_N(_02480_),
    .B(_02468_),
    .Y(_02481_));
 sky130_fd_sc_hd__xnor2_4 _09393_ (.A(_02468_),
    .B(_02480_),
    .Y(_02482_));
 sky130_fd_sc_hd__o21a_1 _09394_ (.A1(_02290_),
    .A2(_02292_),
    .B1(_02288_),
    .X(_02483_));
 sky130_fd_sc_hd__a21o_1 _09395_ (.A1(_00188_),
    .A2(_00189_),
    .B1(net113),
    .X(_02484_));
 sky130_fd_sc_hd__or2_1 _09396_ (.A(net123),
    .B(net65),
    .X(_02485_));
 sky130_fd_sc_hd__and3_1 _09397_ (.A(net93),
    .B(_02484_),
    .C(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__a21oi_1 _09398_ (.A1(_02484_),
    .A2(_02485_),
    .B1(net93),
    .Y(_02487_));
 sky130_fd_sc_hd__a21o_1 _09399_ (.A1(_06552_),
    .A2(_06553_),
    .B1(net98),
    .X(_02488_));
 sky130_fd_sc_hd__or2_1 _09400_ (.A(_06558_),
    .B(net96),
    .X(_02489_));
 sky130_fd_sc_hd__and3_1 _09401_ (.A(net107),
    .B(_02488_),
    .C(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__a21oi_1 _09402_ (.A1(_02488_),
    .A2(_02489_),
    .B1(net107),
    .Y(_02491_));
 sky130_fd_sc_hd__o22a_1 _09403_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_02490_),
    .B2(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__or4_1 _09404_ (.A(_02486_),
    .B(_02487_),
    .C(_02490_),
    .D(_02491_),
    .X(_02493_));
 sky130_fd_sc_hd__and2b_1 _09405_ (.A_N(_02492_),
    .B(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__o22a_1 _09406_ (.A1(net117),
    .A2(_00181_),
    .B1(net89),
    .B2(net22),
    .X(_02495_));
 sky130_fd_sc_hd__xnor2_2 _09407_ (.A(net103),
    .B(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__xor2_2 _09408_ (.A(_02494_),
    .B(_02496_),
    .X(_02497_));
 sky130_fd_sc_hd__a31o_1 _09409_ (.A1(_06526_),
    .A2(net35),
    .A3(_02346_),
    .B1(_02345_),
    .X(_02498_));
 sky130_fd_sc_hd__nand2_1 _09410_ (.A(_02497_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__xor2_1 _09411_ (.A(_02497_),
    .B(_02498_),
    .X(_02500_));
 sky130_fd_sc_hd__nand2b_1 _09412_ (.A_N(_02483_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__xnor2_1 _09413_ (.A(_02483_),
    .B(_02500_),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ai_2 _09414_ (.A1(_02322_),
    .A2(_02324_),
    .B1(_02320_),
    .Y(_02503_));
 sky130_fd_sc_hd__or2_1 _09415_ (.A(_02309_),
    .B(_02313_),
    .X(_02504_));
 sky130_fd_sc_hd__a21oi_2 _09416_ (.A1(_02363_),
    .A2(_02366_),
    .B1(_02362_),
    .Y(_02505_));
 sky130_fd_sc_hd__o21bai_1 _09417_ (.A1(_02309_),
    .A2(_02313_),
    .B1_N(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__xnor2_1 _09418_ (.A(_02504_),
    .B(_02505_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _09419_ (.A(_02503_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__xnor2_1 _09420_ (.A(_02503_),
    .B(_02507_),
    .Y(_02509_));
 sky130_fd_sc_hd__or2_1 _09421_ (.A(net183),
    .B(net32),
    .X(_02510_));
 sky130_fd_sc_hd__a21o_1 _09422_ (.A1(_02327_),
    .A2(_02334_),
    .B1(_02332_),
    .X(_02511_));
 sky130_fd_sc_hd__o22a_1 _09423_ (.A1(net144),
    .A2(net11),
    .B1(net5),
    .B2(net180),
    .X(_02512_));
 sky130_fd_sc_hd__xnor2_1 _09424_ (.A(net35),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__nand2_1 _09425_ (.A(_02511_),
    .B(_02513_),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _09426_ (.A(_02511_),
    .B(_02513_),
    .Y(_02515_));
 sky130_fd_sc_hd__or2_1 _09427_ (.A(_02511_),
    .B(_02513_),
    .X(_02516_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(_02514_),
    .B(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__xor2_1 _09429_ (.A(_02510_),
    .B(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__o22a_1 _09430_ (.A1(net46),
    .A2(net88),
    .B1(net83),
    .B2(net55),
    .X(_02519_));
 sky130_fd_sc_hd__xnor2_1 _09431_ (.A(_06469_),
    .B(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__o22a_1 _09432_ (.A1(net60),
    .A2(net132),
    .B1(net170),
    .B2(net57),
    .X(_02521_));
 sky130_fd_sc_hd__xnor2_1 _09433_ (.A(net195),
    .B(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__nor2_1 _09434_ (.A(_02520_),
    .B(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__xor2_1 _09435_ (.A(_02520_),
    .B(_02522_),
    .X(_02524_));
 sky130_fd_sc_hd__o22a_1 _09436_ (.A1(net52),
    .A2(net130),
    .B1(net128),
    .B2(net63),
    .X(_02525_));
 sky130_fd_sc_hd__xnor2_1 _09437_ (.A(net167),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__inv_2 _09438_ (.A(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__xnor2_1 _09439_ (.A(_02524_),
    .B(_02526_),
    .Y(_02528_));
 sky130_fd_sc_hd__o22a_1 _09440_ (.A1(net19),
    .A2(net134),
    .B1(net172),
    .B2(net14),
    .X(_02529_));
 sky130_fd_sc_hd__xnor2_2 _09441_ (.A(net211),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _09442_ (.A(net260),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__xnor2_2 _09443_ (.A(_00213_),
    .B(_02530_),
    .Y(_02532_));
 sky130_fd_sc_hd__nor2_1 _09444_ (.A(net178),
    .B(net7),
    .Y(_02533_));
 sky130_fd_sc_hd__xnor2_2 _09445_ (.A(net213),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__xnor2_2 _09446_ (.A(_02532_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__o22a_1 _09447_ (.A1(net121),
    .A2(net48),
    .B1(net39),
    .B2(net125),
    .X(_02536_));
 sky130_fd_sc_hd__xnor2_1 _09448_ (.A(net153),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__o22a_1 _09449_ (.A1(net119),
    .A2(net69),
    .B1(net95),
    .B2(net85),
    .X(_02538_));
 sky130_fd_sc_hd__xnor2_1 _09450_ (.A(_00153_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__or2_1 _09451_ (.A(_02537_),
    .B(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_02537_),
    .B(_02539_),
    .Y(_02541_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(_02540_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__o22a_1 _09454_ (.A1(net75),
    .A2(net80),
    .B1(net42),
    .B2(_06507_),
    .X(_02543_));
 sky130_fd_sc_hd__xnor2_2 _09455_ (.A(_06500_),
    .B(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__xnor2_2 _09456_ (.A(_02542_),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _09457_ (.A(_02535_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand2_1 _09458_ (.A(_02535_),
    .B(_02545_),
    .Y(_02547_));
 sky130_fd_sc_hd__xnor2_1 _09459_ (.A(_02535_),
    .B(_02545_),
    .Y(_02548_));
 sky130_fd_sc_hd__xnor2_1 _09460_ (.A(_02528_),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_1 _09461_ (.A(_02518_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__xnor2_1 _09462_ (.A(_02518_),
    .B(_02549_),
    .Y(_02551_));
 sky130_fd_sc_hd__xor2_1 _09463_ (.A(_02509_),
    .B(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__and2_1 _09464_ (.A(_02502_),
    .B(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__nor2_1 _09465_ (.A(_02502_),
    .B(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_2 _09466_ (.A(_02553_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__xor2_4 _09467_ (.A(_02482_),
    .B(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__a21o_2 _09468_ (.A1(_02298_),
    .A2(_02373_),
    .B1(_02372_),
    .X(_02557_));
 sky130_fd_sc_hd__or2_4 _09469_ (.A(_02294_),
    .B(_02297_),
    .X(_02558_));
 sky130_fd_sc_hd__o21bai_4 _09470_ (.A1(_02304_),
    .A2(_02349_),
    .B1_N(_02348_),
    .Y(_02559_));
 sky130_fd_sc_hd__a21bo_2 _09471_ (.A1(_02353_),
    .A2(_02370_),
    .B1_N(_02369_),
    .X(_02560_));
 sky130_fd_sc_hd__nand2_1 _09472_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__xor2_4 _09473_ (.A(_02559_),
    .B(_02560_),
    .X(_02562_));
 sky130_fd_sc_hd__xnor2_4 _09474_ (.A(_02558_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__a21oi_4 _09475_ (.A1(_02377_),
    .A2(_02381_),
    .B1(_02380_),
    .Y(_02564_));
 sky130_fd_sc_hd__xnor2_2 _09476_ (.A(_02563_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand2b_1 _09477_ (.A_N(_02565_),
    .B(_02557_),
    .Y(_02566_));
 sky130_fd_sc_hd__xnor2_4 _09478_ (.A(_02557_),
    .B(_02565_),
    .Y(_02567_));
 sky130_fd_sc_hd__and2_1 _09479_ (.A(_02556_),
    .B(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__xor2_4 _09480_ (.A(_02556_),
    .B(_02567_),
    .X(_02569_));
 sky130_fd_sc_hd__xnor2_4 _09481_ (.A(_02467_),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__or2_2 _09482_ (.A(_02466_),
    .B(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__and2_1 _09483_ (.A(_02466_),
    .B(_02570_),
    .X(_02572_));
 sky130_fd_sc_hd__xnor2_4 _09484_ (.A(_02466_),
    .B(_02570_),
    .Y(_02573_));
 sky130_fd_sc_hd__or4_1 _09485_ (.A(_00776_),
    .B(_02057_),
    .C(_02062_),
    .D(_02392_),
    .X(_02574_));
 sky130_fd_sc_hd__a21o_1 _09486_ (.A1(_00774_),
    .A2(_02390_),
    .B1(_02391_),
    .X(_02575_));
 sky130_fd_sc_hd__or4_1 _09487_ (.A(_00776_),
    .B(_02060_),
    .C(_02064_),
    .D(_02392_),
    .X(_02576_));
 sky130_fd_sc_hd__o211a_2 _09488_ (.A1(_02159_),
    .A2(_02574_),
    .B1(_02575_),
    .C1(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__xnor2_1 _09489_ (.A(_02573_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__o21ai_1 _09490_ (.A1(_02465_),
    .A2(_02578_),
    .B1(_02171_),
    .Y(_02579_));
 sky130_fd_sc_hd__a21o_1 _09491_ (.A1(_02465_),
    .A2(_02578_),
    .B1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__a21oi_1 _09492_ (.A1(_01771_),
    .A2(net161),
    .B1(_02075_),
    .Y(_02581_));
 sky130_fd_sc_hd__a311o_1 _09493_ (.A1(_01769_),
    .A2(_01771_),
    .A3(net161),
    .B1(_02254_),
    .C1(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__o21ai_1 _09494_ (.A1(net233),
    .A2(_02424_),
    .B1(_02266_),
    .Y(_02583_));
 sky130_fd_sc_hd__a21oi_2 _09495_ (.A1(net238),
    .A2(_02583_),
    .B1(_02268_),
    .Y(_02584_));
 sky130_fd_sc_hd__inv_2 _09496_ (.A(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__o21ai_2 _09497_ (.A1(net240),
    .A2(_02584_),
    .B1(_02272_),
    .Y(_02586_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(_02181_),
    .A1(_02188_),
    .S(net230),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _09499_ (.A0(_02185_),
    .A1(_02203_),
    .S(net230),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(_02587_),
    .A1(_02588_),
    .S(net233),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _09501_ (.A0(_02193_),
    .A1(_02219_),
    .S(net230),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _09502_ (.A0(_02196_),
    .A1(_02200_),
    .S(net231),
    .X(_02591_));
 sky130_fd_sc_hd__mux2_1 _09503_ (.A0(_02590_),
    .A1(_02591_),
    .S(_06337_),
    .X(_02592_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(_02589_),
    .A1(_02592_),
    .S(net237),
    .X(_02593_));
 sky130_fd_sc_hd__mux2_1 _09505_ (.A0(_02209_),
    .A1(_02234_),
    .S(_06345_),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(_02212_),
    .A1(_02216_),
    .S(net232),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _09507_ (.A0(_02594_),
    .A1(_02595_),
    .S(net235),
    .X(_02596_));
 sky130_fd_sc_hd__mux2_1 _09508_ (.A0(_02227_),
    .A1(_02231_),
    .S(net231),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_1 _09509_ (.A0(_02455_),
    .A1(_02597_),
    .S(net235),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _09510_ (.A0(_02596_),
    .A1(_02598_),
    .S(net236),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _09511_ (.A0(_02593_),
    .A1(_02599_),
    .S(net240),
    .X(_02600_));
 sky130_fd_sc_hd__inv_2 _09512_ (.A(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__o21a_1 _09513_ (.A1(_02239_),
    .A2(_02434_),
    .B1(_02432_),
    .X(_02602_));
 sky130_fd_sc_hd__nor2_1 _09514_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02603_));
 sky130_fd_sc_hd__nand2_1 _09515_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02604_));
 sky130_fd_sc_hd__nand2b_1 _09516_ (.A_N(_02603_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__xor2_1 _09517_ (.A(_02602_),
    .B(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__nor2_1 _09518_ (.A(net243),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__or2_1 _09519_ (.A(\div_res[1] ),
    .B(\div_res[0] ),
    .X(_02608_));
 sky130_fd_sc_hd__a21oi_1 _09520_ (.A1(net165),
    .A2(_02608_),
    .B1(\div_res[2] ),
    .Y(_02609_));
 sky130_fd_sc_hd__a31o_1 _09521_ (.A1(\div_res[2] ),
    .A2(net165),
    .A3(_02608_),
    .B1(net205),
    .X(_02610_));
 sky130_fd_sc_hd__a22o_1 _09522_ (.A1(net307),
    .A2(_06345_),
    .B1(net224),
    .B2(net308),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _09523_ (.A(_06347_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__mux2_1 _09524_ (.A0(_06353_),
    .A1(_02612_),
    .S(net304),
    .X(_02613_));
 sky130_fd_sc_hd__nor2_1 _09525_ (.A(_06342_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__a21o_1 _09526_ (.A1(_06342_),
    .A2(_02613_),
    .B1(net255),
    .X(_02615_));
 sky130_fd_sc_hd__or2_1 _09527_ (.A(_06342_),
    .B(net253),
    .X(_02616_));
 sky130_fd_sc_hd__or2_1 _09528_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .X(_02617_));
 sky130_fd_sc_hd__a21oi_1 _09529_ (.A1(net247),
    .A2(_02617_),
    .B1(\div_shifter[34] ),
    .Y(_02618_));
 sky130_fd_sc_hd__a31o_1 _09530_ (.A1(\div_shifter[34] ),
    .A2(net247),
    .A3(_02617_),
    .B1(net250),
    .X(_02619_));
 sky130_fd_sc_hd__o22a_1 _09531_ (.A1(net235),
    .A2(net215),
    .B1(_02618_),
    .B2(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__nor2_1 _09532_ (.A(net309),
    .B(_02600_),
    .Y(_02621_));
 sky130_fd_sc_hd__a211o_1 _09533_ (.A1(net309),
    .A2(_02586_),
    .B1(_02621_),
    .C1(_06451_),
    .X(_02622_));
 sky130_fd_sc_hd__a211o_1 _09534_ (.A1(net244),
    .A2(_02601_),
    .B1(_02607_),
    .C1(_06447_),
    .X(_02623_));
 sky130_fd_sc_hd__o221a_1 _09535_ (.A1(_06340_),
    .A2(net208),
    .B1(net206),
    .B2(_06341_),
    .C1(_02620_),
    .X(_02624_));
 sky130_fd_sc_hd__o211a_1 _09536_ (.A1(_02609_),
    .A2(_02610_),
    .B1(_02616_),
    .C1(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__o211a_1 _09537_ (.A1(_02614_),
    .A2(_02615_),
    .B1(_02623_),
    .C1(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__a41o_2 _09538_ (.A1(_02580_),
    .A2(_02582_),
    .A3(_02622_),
    .A4(_02626_),
    .B1(_06424_),
    .X(_02627_));
 sky130_fd_sc_hd__and3_1 _09539_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .X(_02628_));
 sky130_fd_sc_hd__a21oi_2 _09540_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .B1(curr_PC[2]),
    .Y(_02629_));
 sky130_fd_sc_hd__o31ai_4 _09541_ (.A1(net262),
    .A2(_02628_),
    .A3(_02629_),
    .B1(_02627_),
    .Y(dest_val[2]));
 sky130_fd_sc_hd__and3_1 _09542_ (.A(_02069_),
    .B(_02398_),
    .C(_02578_),
    .X(_02630_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_02167_),
    .B(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__a21oi_4 _09544_ (.A1(_02467_),
    .A2(_02569_),
    .B1(_02568_),
    .Y(_02632_));
 sky130_fd_sc_hd__o21ai_4 _09545_ (.A1(_02563_),
    .A2(_02564_),
    .B1(_02566_),
    .Y(_02633_));
 sky130_fd_sc_hd__a21o_2 _09546_ (.A1(_02528_),
    .A2(_02547_),
    .B1(_02546_),
    .X(_02634_));
 sky130_fd_sc_hd__o22a_1 _09547_ (.A1(net146),
    .A2(net16),
    .B1(_00354_),
    .B2(net142),
    .X(_02635_));
 sky130_fd_sc_hd__xnor2_1 _09548_ (.A(net78),
    .B(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__o22a_1 _09549_ (.A1(_00143_),
    .A2(net99),
    .B1(net135),
    .B2(net23),
    .X(_02637_));
 sky130_fd_sc_hd__xor2_1 _09550_ (.A(net110),
    .B(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__or2_1 _09551_ (.A(_02636_),
    .B(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__nand2_1 _09552_ (.A(_02636_),
    .B(_02638_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _09553_ (.A(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__o22a_1 _09554_ (.A1(net30),
    .A2(_00180_),
    .B1(net137),
    .B2(net28),
    .X(_02642_));
 sky130_fd_sc_hd__xnor2_2 _09555_ (.A(_06524_),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__xnor2_1 _09556_ (.A(_02641_),
    .B(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__a21oi_1 _09557_ (.A1(_02506_),
    .A2(_02508_),
    .B1(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__and3_1 _09558_ (.A(_02506_),
    .B(_02508_),
    .C(_02644_),
    .X(_02646_));
 sky130_fd_sc_hd__nor2_2 _09559_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__xor2_4 _09560_ (.A(_02634_),
    .B(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__o21a_1 _09561_ (.A1(_02542_),
    .A2(_02544_),
    .B1(_02540_),
    .X(_02649_));
 sky130_fd_sc_hd__a21o_1 _09562_ (.A1(_02524_),
    .A2(_02527_),
    .B1(_02523_),
    .X(_02650_));
 sky130_fd_sc_hd__a21o_1 _09563_ (.A1(_02493_),
    .A2(_02496_),
    .B1(_02492_),
    .X(_02651_));
 sky130_fd_sc_hd__xor2_2 _09564_ (.A(_02650_),
    .B(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__and2b_1 _09565_ (.A_N(_02649_),
    .B(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__xnor2_2 _09566_ (.A(_02649_),
    .B(_02652_),
    .Y(_02654_));
 sky130_fd_sc_hd__or2_1 _09567_ (.A(net57),
    .B(net132),
    .X(_02655_));
 sky130_fd_sc_hd__or2_1 _09568_ (.A(net18),
    .B(net170),
    .X(_02656_));
 sky130_fd_sc_hd__a21o_1 _09569_ (.A1(_02655_),
    .A2(_02656_),
    .B1(net194),
    .X(_02657_));
 sky130_fd_sc_hd__nand3_1 _09570_ (.A(net194),
    .B(_02655_),
    .C(_02656_),
    .Y(_02658_));
 sky130_fd_sc_hd__o22a_1 _09571_ (.A1(net54),
    .A2(net88),
    .B1(net83),
    .B2(net51),
    .X(_02659_));
 sky130_fd_sc_hd__xnor2_1 _09572_ (.A(_06470_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__and3_1 _09573_ (.A(_02657_),
    .B(_02658_),
    .C(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__a21oi_1 _09574_ (.A1(_02657_),
    .A2(_02658_),
    .B1(_02660_),
    .Y(_02662_));
 sky130_fd_sc_hd__nor2_1 _09575_ (.A(_02661_),
    .B(_02662_),
    .Y(_02663_));
 sky130_fd_sc_hd__o22a_1 _09576_ (.A1(net63),
    .A2(net130),
    .B1(net128),
    .B2(net60),
    .X(_02664_));
 sky130_fd_sc_hd__xnor2_2 _09577_ (.A(net167),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__xnor2_2 _09578_ (.A(_02663_),
    .B(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__o22a_1 _09579_ (.A1(net125),
    .A2(net47),
    .B1(net45),
    .B2(net121),
    .X(_02667_));
 sky130_fd_sc_hd__xnor2_1 _09580_ (.A(net152),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__o22a_1 _09581_ (.A1(net68),
    .A2(net85),
    .B1(net79),
    .B2(net94),
    .X(_02669_));
 sky130_fd_sc_hd__xnor2_1 _09582_ (.A(_00153_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nor2_1 _09583_ (.A(_02668_),
    .B(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__xnor2_1 _09584_ (.A(_02668_),
    .B(_02670_),
    .Y(_02672_));
 sky130_fd_sc_hd__o22a_1 _09585_ (.A1(net75),
    .A2(net41),
    .B1(net38),
    .B2(net116),
    .X(_02673_));
 sky130_fd_sc_hd__xnor2_1 _09586_ (.A(_06500_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__nor2_1 _09587_ (.A(_02672_),
    .B(_02674_),
    .Y(_02675_));
 sky130_fd_sc_hd__and2_1 _09588_ (.A(_02672_),
    .B(_02674_),
    .X(_02676_));
 sky130_fd_sc_hd__or2_1 _09589_ (.A(_02675_),
    .B(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__o22a_1 _09590_ (.A1(net134),
    .A2(net14),
    .B1(net7),
    .B2(_00258_),
    .X(_02678_));
 sky130_fd_sc_hd__xnor2_1 _09591_ (.A(_00250_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__or2_1 _09592_ (.A(_00213_),
    .B(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__xnor2_2 _09593_ (.A(_00213_),
    .B(_02679_),
    .Y(_02681_));
 sky130_fd_sc_hd__xnor2_2 _09594_ (.A(_00210_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__nor2_1 _09595_ (.A(_02677_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__xor2_2 _09596_ (.A(_02677_),
    .B(_02682_),
    .X(_02684_));
 sky130_fd_sc_hd__xor2_2 _09597_ (.A(_02666_),
    .B(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_1 _09598_ (.A(_06565_),
    .B(net35),
    .Y(_02686_));
 sky130_fd_sc_hd__a21oi_2 _09599_ (.A1(_02532_),
    .A2(_02534_),
    .B1(_02531_),
    .Y(_02687_));
 sky130_fd_sc_hd__o22a_1 _09600_ (.A1(_06547_),
    .A2(net11),
    .B1(net5),
    .B2(net144),
    .X(_02688_));
 sky130_fd_sc_hd__xnor2_2 _09601_ (.A(net35),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__and2b_1 _09602_ (.A_N(_02687_),
    .B(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__xnor2_2 _09603_ (.A(_02687_),
    .B(_02689_),
    .Y(_02691_));
 sky130_fd_sc_hd__xnor2_2 _09604_ (.A(_02686_),
    .B(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__and2_1 _09605_ (.A(_02685_),
    .B(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__xor2_2 _09606_ (.A(_02685_),
    .B(_02692_),
    .X(_02694_));
 sky130_fd_sc_hd__xor2_1 _09607_ (.A(_02654_),
    .B(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__o21a_1 _09608_ (.A1(_02475_),
    .A2(_02477_),
    .B1(_02473_),
    .X(_02696_));
 sky130_fd_sc_hd__or2_1 _09609_ (.A(net123),
    .B(net21),
    .X(_02697_));
 sky130_fd_sc_hd__or2_1 _09610_ (.A(net119),
    .B(_00192_),
    .X(_02698_));
 sky130_fd_sc_hd__and3_1 _09611_ (.A(net93),
    .B(_02697_),
    .C(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__a21oi_1 _09612_ (.A1(_02697_),
    .A2(_02698_),
    .B1(net93),
    .Y(_02700_));
 sky130_fd_sc_hd__or2_1 _09613_ (.A(net26),
    .B(net96),
    .X(_02701_));
 sky130_fd_sc_hd__or2_1 _09614_ (.A(net73),
    .B(net89),
    .X(_02702_));
 sky130_fd_sc_hd__and3_1 _09615_ (.A(net107),
    .B(_02701_),
    .C(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__a21oi_1 _09616_ (.A1(_02701_),
    .A2(_02702_),
    .B1(net107),
    .Y(_02704_));
 sky130_fd_sc_hd__o22a_1 _09617_ (.A1(_02699_),
    .A2(_02700_),
    .B1(_02703_),
    .B2(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__or4_1 _09618_ (.A(_02699_),
    .B(_02700_),
    .C(_02703_),
    .D(_02704_),
    .X(_02706_));
 sky130_fd_sc_hd__nand2b_1 _09619_ (.A_N(_02705_),
    .B(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__o22a_1 _09620_ (.A1(net117),
    .A2(net22),
    .B1(net67),
    .B2(net113),
    .X(_02708_));
 sky130_fd_sc_hd__xnor2_2 _09621_ (.A(net103),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__xnor2_2 _09622_ (.A(_02707_),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__o21ai_1 _09623_ (.A1(_02510_),
    .A2(_02515_),
    .B1(_02514_),
    .Y(_02711_));
 sky130_fd_sc_hd__xor2_1 _09624_ (.A(_02710_),
    .B(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__and2b_1 _09625_ (.A_N(_02696_),
    .B(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__xnor2_1 _09626_ (.A(_02696_),
    .B(_02712_),
    .Y(_02714_));
 sky130_fd_sc_hd__and2_1 _09627_ (.A(_02695_),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__nor2_1 _09628_ (.A(_02695_),
    .B(_02714_),
    .Y(_02716_));
 sky130_fd_sc_hd__nor2_2 _09629_ (.A(_02715_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__xor2_4 _09630_ (.A(_02648_),
    .B(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__a21o_2 _09631_ (.A1(_02482_),
    .A2(_02555_),
    .B1(_02553_),
    .X(_02719_));
 sky130_fd_sc_hd__o21ai_4 _09632_ (.A1(_02478_),
    .A2(_02479_),
    .B1(_02481_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand2_2 _09633_ (.A(_02499_),
    .B(_02501_),
    .Y(_02721_));
 sky130_fd_sc_hd__o21a_2 _09634_ (.A1(_02509_),
    .A2(_02551_),
    .B1(_02550_),
    .X(_02722_));
 sky130_fd_sc_hd__a21o_1 _09635_ (.A1(_02499_),
    .A2(_02501_),
    .B1(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__xnor2_4 _09636_ (.A(_02721_),
    .B(_02722_),
    .Y(_02724_));
 sky130_fd_sc_hd__xnor2_4 _09637_ (.A(_02720_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__a21boi_4 _09638_ (.A1(_02558_),
    .A2(_02562_),
    .B1_N(_02561_),
    .Y(_02726_));
 sky130_fd_sc_hd__xnor2_4 _09639_ (.A(_02725_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__nand2b_1 _09640_ (.A_N(_02727_),
    .B(_02719_),
    .Y(_02728_));
 sky130_fd_sc_hd__xnor2_4 _09641_ (.A(_02719_),
    .B(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__and2_1 _09642_ (.A(_02718_),
    .B(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__xor2_4 _09643_ (.A(_02718_),
    .B(_02729_),
    .X(_02731_));
 sky130_fd_sc_hd__xnor2_4 _09644_ (.A(_02633_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__or2_2 _09645_ (.A(_02632_),
    .B(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__and2_1 _09646_ (.A(_02632_),
    .B(_02732_),
    .X(_02734_));
 sky130_fd_sc_hd__xnor2_4 _09647_ (.A(_02632_),
    .B(_02732_),
    .Y(_02735_));
 sky130_fd_sc_hd__nor2_1 _09648_ (.A(_02392_),
    .B(_02573_),
    .Y(_02736_));
 sky130_fd_sc_hd__nor4_1 _09649_ (.A(_00776_),
    .B(_02062_),
    .C(_02392_),
    .D(_02573_),
    .Y(_02737_));
 sky130_fd_sc_hd__a21oi_2 _09650_ (.A1(_02390_),
    .A2(_02571_),
    .B1(_02572_),
    .Y(_02738_));
 sky130_fd_sc_hd__a221oi_4 _09651_ (.A1(_02394_),
    .A2(_02736_),
    .B1(net3),
    .B2(_02165_),
    .C1(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__xor2_4 _09652_ (.A(_02735_),
    .B(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__nand3_1 _09653_ (.A(net161),
    .B(_02631_),
    .C(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__a21o_1 _09654_ (.A1(net161),
    .A2(_02631_),
    .B1(_02740_),
    .X(_02742_));
 sky130_fd_sc_hd__and3_1 _09655_ (.A(_02171_),
    .B(_02741_),
    .C(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__or3_1 _09656_ (.A(net158),
    .B(_02073_),
    .C(_02076_),
    .X(_02744_));
 sky130_fd_sc_hd__o21ai_1 _09657_ (.A1(net158),
    .A2(_02076_),
    .B1(_02073_),
    .Y(_02745_));
 sky130_fd_sc_hd__and3_1 _09658_ (.A(_02253_),
    .B(_02744_),
    .C(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _09659_ (.A0(_02402_),
    .A1(_02405_),
    .S(net230),
    .X(_02747_));
 sky130_fd_sc_hd__mux2_1 _09660_ (.A0(_02404_),
    .A1(_02412_),
    .S(net230),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _09661_ (.A0(_02747_),
    .A1(_02748_),
    .S(net233),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _09662_ (.A0(_02408_),
    .A1(_02420_),
    .S(net230),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _09663_ (.A0(_02409_),
    .A1(_02411_),
    .S(net231),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(_02750_),
    .A1(_02751_),
    .S(net235),
    .X(_02752_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(_02749_),
    .A1(_02752_),
    .S(net237),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _09666_ (.A0(_02416_),
    .A1(_02426_),
    .S(net230),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(_02417_),
    .A1(_02419_),
    .S(net232),
    .X(_02755_));
 sky130_fd_sc_hd__mux2_1 _09668_ (.A0(_02754_),
    .A1(_02755_),
    .S(net235),
    .X(_02756_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(_02423_),
    .A1(_02425_),
    .S(net232),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(_02265_),
    .A1(_02757_),
    .S(net235),
    .X(_02758_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(_02756_),
    .A1(_02758_),
    .S(net236),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_2 _09672_ (.A0(_02753_),
    .A1(_02759_),
    .S(net240),
    .X(_02760_));
 sky130_fd_sc_hd__o21a_1 _09673_ (.A1(_02602_),
    .A2(_02603_),
    .B1(_02604_),
    .X(_02761_));
 sky130_fd_sc_hd__nor2_1 _09674_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02762_));
 sky130_fd_sc_hd__or2_1 _09675_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .X(_02763_));
 sky130_fd_sc_hd__nand2_1 _09676_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02764_));
 sky130_fd_sc_hd__a21oi_1 _09677_ (.A1(_02763_),
    .A2(_02764_),
    .B1(_02761_),
    .Y(_02765_));
 sky130_fd_sc_hd__a31o_1 _09678_ (.A1(_02761_),
    .A2(_02763_),
    .A3(_02764_),
    .B1(net243),
    .X(_02766_));
 sky130_fd_sc_hd__o221a_1 _09679_ (.A1(net268),
    .A2(_02760_),
    .B1(_02765_),
    .B2(_02766_),
    .C1(net216),
    .X(_02767_));
 sky130_fd_sc_hd__o21a_1 _09680_ (.A1(net233),
    .A2(_02228_),
    .B1(_02266_),
    .X(_02768_));
 sky130_fd_sc_hd__o21a_1 _09681_ (.A1(net236),
    .A2(_02768_),
    .B1(_02269_),
    .X(_02769_));
 sky130_fd_sc_hd__o21a_1 _09682_ (.A1(net240),
    .A2(_02769_),
    .B1(_02272_),
    .X(_02770_));
 sky130_fd_sc_hd__a21boi_1 _09683_ (.A1(_06347_),
    .A2(_02611_),
    .B1_N(_06341_),
    .Y(_02771_));
 sky130_fd_sc_hd__or3_1 _09684_ (.A(net310),
    .B(_06340_),
    .C(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__o21ai_1 _09685_ (.A1(net304),
    .A2(_06354_),
    .B1(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2b_1 _09686_ (.A_N(_02773_),
    .B(_06335_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2b_1 _09687_ (.A_N(_06335_),
    .B(_02773_),
    .Y(_02775_));
 sky130_fd_sc_hd__or3_1 _09688_ (.A(\div_res[2] ),
    .B(\div_res[1] ),
    .C(\div_res[0] ),
    .X(_02776_));
 sky130_fd_sc_hd__a21oi_1 _09689_ (.A1(net165),
    .A2(_02776_),
    .B1(\div_res[3] ),
    .Y(_02777_));
 sky130_fd_sc_hd__a31o_1 _09690_ (.A1(\div_res[3] ),
    .A2(net165),
    .A3(_02776_),
    .B1(net205),
    .X(_02778_));
 sky130_fd_sc_hd__o31a_1 _09691_ (.A1(\div_shifter[34] ),
    .A2(\div_shifter[33] ),
    .A3(\div_shifter[32] ),
    .B1(net247),
    .X(_02779_));
 sky130_fd_sc_hd__o21ai_1 _09692_ (.A1(\div_shifter[35] ),
    .A2(_02779_),
    .B1(_02258_),
    .Y(_02780_));
 sky130_fd_sc_hd__a21o_1 _09693_ (.A1(\div_shifter[35] ),
    .A2(_02779_),
    .B1(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__o221a_1 _09694_ (.A1(net238),
    .A2(_06460_),
    .B1(net206),
    .B2(_06334_),
    .C1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__o221a_1 _09695_ (.A1(_06333_),
    .A2(net208),
    .B1(net254),
    .B2(_06335_),
    .C1(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__o21ai_1 _09696_ (.A1(_02777_),
    .A2(_02778_),
    .B1(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__a31o_1 _09697_ (.A1(_02247_),
    .A2(_02774_),
    .A3(_02775_),
    .B1(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__a221o_1 _09698_ (.A1(_02243_),
    .A2(_02760_),
    .B1(_02770_),
    .B2(net192),
    .C1(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__or4_2 _09699_ (.A(_02743_),
    .B(_02746_),
    .C(_02767_),
    .D(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__or2_1 _09700_ (.A(curr_PC[3]),
    .B(_02628_),
    .X(_02788_));
 sky130_fd_sc_hd__and2_1 _09701_ (.A(curr_PC[3]),
    .B(_02628_),
    .X(_02789_));
 sky130_fd_sc_hd__nor2_1 _09702_ (.A(net262),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__a22o_4 _09703_ (.A1(net262),
    .A2(_02787_),
    .B1(_02788_),
    .B2(_02790_),
    .X(dest_val[3]));
 sky130_fd_sc_hd__o21a_1 _09704_ (.A1(_02631_),
    .A2(_02740_),
    .B1(net161),
    .X(_02791_));
 sky130_fd_sc_hd__or2_1 _09705_ (.A(_02573_),
    .B(_02735_),
    .X(_02792_));
 sky130_fd_sc_hd__or4_1 _09706_ (.A(_00776_),
    .B(_02392_),
    .C(_02573_),
    .D(_02735_),
    .X(_02793_));
 sky130_fd_sc_hd__a21o_1 _09707_ (.A1(_02063_),
    .A2(_02067_),
    .B1(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__a21o_1 _09708_ (.A1(_02571_),
    .A2(_02733_),
    .B1(_02734_),
    .X(_02795_));
 sky130_fd_sc_hd__o21a_2 _09709_ (.A1(_02575_),
    .A2(_02792_),
    .B1(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__a21oi_4 _09710_ (.A1(_02633_),
    .A2(_02731_),
    .B1(_02730_),
    .Y(_02797_));
 sky130_fd_sc_hd__o21ai_4 _09711_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02728_),
    .Y(_02798_));
 sky130_fd_sc_hd__a21o_2 _09712_ (.A1(_02666_),
    .A2(_02684_),
    .B1(_02683_),
    .X(_02799_));
 sky130_fd_sc_hd__o22a_1 _09713_ (.A1(net142),
    .A2(net16),
    .B1(net37),
    .B2(net140),
    .X(_02800_));
 sky130_fd_sc_hd__xnor2_1 _09714_ (.A(net77),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__o22a_1 _09715_ (.A1(net23),
    .A2(net98),
    .B1(net96),
    .B2(net71),
    .X(_02802_));
 sky130_fd_sc_hd__xor2_1 _09716_ (.A(net110),
    .B(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__or2_2 _09717_ (.A(_02801_),
    .B(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(_02801_),
    .B(_02803_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2_4 _09719_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__o22a_2 _09720_ (.A1(net30),
    .A2(net137),
    .B1(net135),
    .B2(net28),
    .X(_02807_));
 sky130_fd_sc_hd__xnor2_4 _09721_ (.A(_06524_),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__xnor2_4 _09722_ (.A(_02806_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__a21oi_2 _09723_ (.A1(_02650_),
    .A2(_02651_),
    .B1(_02653_),
    .Y(_02810_));
 sky130_fd_sc_hd__xnor2_2 _09724_ (.A(_02809_),
    .B(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2b_1 _09725_ (.A_N(_02811_),
    .B(_02799_),
    .Y(_02812_));
 sky130_fd_sc_hd__xnor2_4 _09726_ (.A(_02799_),
    .B(_02811_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21oi_1 _09727_ (.A1(_02706_),
    .A2(_02709_),
    .B1(_02705_),
    .Y(_02814_));
 sky130_fd_sc_hd__o21ba_1 _09728_ (.A1(_02662_),
    .A2(_02665_),
    .B1_N(_02661_),
    .X(_02815_));
 sky130_fd_sc_hd__nor2_1 _09729_ (.A(_02814_),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__xor2_1 _09730_ (.A(_02814_),
    .B(_02815_),
    .X(_02817_));
 sky130_fd_sc_hd__o21a_1 _09731_ (.A1(_02671_),
    .A2(_02675_),
    .B1(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__nor3_1 _09732_ (.A(_02671_),
    .B(_02675_),
    .C(_02817_),
    .Y(_02819_));
 sky130_fd_sc_hd__or2_1 _09733_ (.A(_02818_),
    .B(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__o22a_1 _09734_ (.A1(net51),
    .A2(net88),
    .B1(net83),
    .B2(net62),
    .X(_02821_));
 sky130_fd_sc_hd__xnor2_2 _09735_ (.A(net186),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__o22a_1 _09736_ (.A1(net121),
    .A2(net54),
    .B1(net44),
    .B2(net125),
    .X(_02823_));
 sky130_fd_sc_hd__xnor2_1 _09737_ (.A(net152),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__o22a_1 _09738_ (.A1(net59),
    .A2(net130),
    .B1(net128),
    .B2(net57),
    .X(_02825_));
 sky130_fd_sc_hd__xnor2_1 _09739_ (.A(net167),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__or2_1 _09740_ (.A(_02824_),
    .B(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_02824_),
    .B(_02826_),
    .Y(_02828_));
 sky130_fd_sc_hd__nand2_1 _09742_ (.A(_02827_),
    .B(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__xor2_2 _09743_ (.A(_02822_),
    .B(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__a21o_1 _09744_ (.A1(_00188_),
    .A2(_00189_),
    .B1(net119),
    .X(_02831_));
 sky130_fd_sc_hd__or2_1 _09745_ (.A(_00192_),
    .B(net85),
    .X(_02832_));
 sky130_fd_sc_hd__nand3_1 _09746_ (.A(net93),
    .B(_02831_),
    .C(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__a21o_1 _09747_ (.A1(_02831_),
    .A2(_02832_),
    .B1(net93),
    .X(_02834_));
 sky130_fd_sc_hd__o22a_1 _09748_ (.A1(net115),
    .A2(net47),
    .B1(net38),
    .B2(net74),
    .X(_02835_));
 sky130_fd_sc_hd__xnor2_1 _09749_ (.A(net149),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__a21oi_1 _09750_ (.A1(_02833_),
    .A2(_02834_),
    .B1(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__and3_1 _09751_ (.A(_02833_),
    .B(_02834_),
    .C(_02836_),
    .X(_02838_));
 sky130_fd_sc_hd__nor2_1 _09752_ (.A(_02837_),
    .B(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__o22a_1 _09753_ (.A1(net68),
    .A2(net79),
    .B1(net41),
    .B2(net94),
    .X(_02840_));
 sky130_fd_sc_hd__xnor2_2 _09754_ (.A(net100),
    .B(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__xor2_2 _09755_ (.A(_02839_),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__o22a_1 _09756_ (.A1(net18),
    .A2(net132),
    .B1(net170),
    .B2(net13),
    .X(_02843_));
 sky130_fd_sc_hd__xor2_1 _09757_ (.A(net194),
    .B(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__or2_1 _09758_ (.A(_00255_),
    .B(net7),
    .X(_02845_));
 sky130_fd_sc_hd__a2bb2o_1 _09759_ (.A1_N(_00254_),
    .A2_N(net7),
    .B1(_02845_),
    .B2(_00249_),
    .X(_02846_));
 sky130_fd_sc_hd__nor2_1 _09760_ (.A(_02844_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__and2_1 _09761_ (.A(_02844_),
    .B(_02846_),
    .X(_02848_));
 sky130_fd_sc_hd__or2_1 _09762_ (.A(_02847_),
    .B(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__and2_1 _09763_ (.A(_02842_),
    .B(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__xor2_2 _09764_ (.A(_02842_),
    .B(_02849_),
    .X(_02851_));
 sky130_fd_sc_hd__xor2_1 _09765_ (.A(_02830_),
    .B(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__or2_1 _09766_ (.A(_00142_),
    .B(net32),
    .X(_02853_));
 sky130_fd_sc_hd__o21a_1 _09767_ (.A1(_00210_),
    .A2(_02681_),
    .B1(_02680_),
    .X(_02854_));
 sky130_fd_sc_hd__o22a_1 _09768_ (.A1(net146),
    .A2(net11),
    .B1(net5),
    .B2(_06547_),
    .X(_02855_));
 sky130_fd_sc_hd__xnor2_1 _09769_ (.A(net35),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__and2b_1 _09770_ (.A_N(_02854_),
    .B(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__xnor2_2 _09771_ (.A(_02854_),
    .B(_02856_),
    .Y(_02858_));
 sky130_fd_sc_hd__xnor2_2 _09772_ (.A(_02853_),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(_02852_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__xnor2_1 _09774_ (.A(_02852_),
    .B(_02859_),
    .Y(_02861_));
 sky130_fd_sc_hd__xnor2_1 _09775_ (.A(_02820_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__o21ai_2 _09776_ (.A1(_02641_),
    .A2(_02643_),
    .B1(_02639_),
    .Y(_02863_));
 sky130_fd_sc_hd__o22a_1 _09777_ (.A1(net117),
    .A2(net72),
    .B1(net89),
    .B2(net26),
    .X(_02864_));
 sky130_fd_sc_hd__xnor2_2 _09778_ (.A(net105),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__o22a_1 _09779_ (.A1(net113),
    .A2(net22),
    .B1(net67),
    .B2(net123),
    .X(_02866_));
 sky130_fd_sc_hd__xnor2_2 _09780_ (.A(net102),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__nand2_1 _09781_ (.A(_02865_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__or2_1 _09782_ (.A(_02865_),
    .B(_02867_),
    .X(_02869_));
 sky130_fd_sc_hd__and2_1 _09783_ (.A(_02868_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__a31o_1 _09784_ (.A1(_06565_),
    .A2(net35),
    .A3(_02691_),
    .B1(_02690_),
    .X(_02871_));
 sky130_fd_sc_hd__nand2_1 _09785_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__xor2_2 _09786_ (.A(_02870_),
    .B(_02871_),
    .X(_02873_));
 sky130_fd_sc_hd__xnor2_1 _09787_ (.A(_02863_),
    .B(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__nor2_1 _09788_ (.A(_02862_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _09789_ (.A(_02862_),
    .B(_02874_),
    .Y(_02876_));
 sky130_fd_sc_hd__and2b_1 _09790_ (.A_N(_02875_),
    .B(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__xor2_4 _09791_ (.A(_02813_),
    .B(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__a21o_2 _09792_ (.A1(_02648_),
    .A2(_02717_),
    .B1(_02715_),
    .X(_02879_));
 sky130_fd_sc_hd__a21bo_1 _09793_ (.A1(_02720_),
    .A2(_02724_),
    .B1_N(_02723_),
    .X(_02880_));
 sky130_fd_sc_hd__a21o_1 _09794_ (.A1(_02634_),
    .A2(_02647_),
    .B1(_02645_),
    .X(_02881_));
 sky130_fd_sc_hd__a21oi_2 _09795_ (.A1(_02654_),
    .A2(_02694_),
    .B1(_02693_),
    .Y(_02882_));
 sky130_fd_sc_hd__a21o_1 _09796_ (.A1(_02710_),
    .A2(_02711_),
    .B1(_02713_),
    .X(_02883_));
 sky130_fd_sc_hd__and2b_1 _09797_ (.A_N(_02882_),
    .B(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__xnor2_2 _09798_ (.A(_02882_),
    .B(_02883_),
    .Y(_02885_));
 sky130_fd_sc_hd__xor2_2 _09799_ (.A(_02881_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__xnor2_2 _09800_ (.A(_02880_),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__nand2b_1 _09801_ (.A_N(_02887_),
    .B(_02879_),
    .Y(_02888_));
 sky130_fd_sc_hd__xnor2_4 _09802_ (.A(_02879_),
    .B(_02887_),
    .Y(_02889_));
 sky130_fd_sc_hd__and2_1 _09803_ (.A(_02878_),
    .B(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__xor2_4 _09804_ (.A(_02878_),
    .B(_02889_),
    .X(_02891_));
 sky130_fd_sc_hd__xnor2_4 _09805_ (.A(_02798_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__or2_1 _09806_ (.A(_02797_),
    .B(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__and2_1 _09807_ (.A(_02797_),
    .B(_02892_),
    .X(_02894_));
 sky130_fd_sc_hd__xnor2_4 _09808_ (.A(_02797_),
    .B(_02892_),
    .Y(_02895_));
 sky130_fd_sc_hd__a21o_1 _09809_ (.A1(_02794_),
    .A2(_02796_),
    .B1(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__nand3_1 _09810_ (.A(_02794_),
    .B(_02796_),
    .C(_02895_),
    .Y(_02897_));
 sky130_fd_sc_hd__and2_1 _09811_ (.A(_02896_),
    .B(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__a21oi_1 _09812_ (.A1(_02791_),
    .A2(_02898_),
    .B1(_02172_),
    .Y(_02899_));
 sky130_fd_sc_hd__o21ai_1 _09813_ (.A1(_02791_),
    .A2(_02898_),
    .B1(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__a21oi_1 _09814_ (.A1(net161),
    .A2(_02077_),
    .B1(_02078_),
    .Y(_02901_));
 sky130_fd_sc_hd__a31o_1 _09815_ (.A1(net161),
    .A2(_02077_),
    .A3(_02078_),
    .B1(_02254_),
    .X(_02902_));
 sky130_fd_sc_hd__o31a_1 _09816_ (.A1(_06333_),
    .A2(_06340_),
    .A3(_02771_),
    .B1(_06334_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(_06355_),
    .A1(_02903_),
    .S(net304),
    .X(_02904_));
 sky130_fd_sc_hd__a21oi_1 _09818_ (.A1(_06328_),
    .A2(_02904_),
    .B1(net255),
    .Y(_02905_));
 sky130_fd_sc_hd__o21ai_1 _09819_ (.A1(_06328_),
    .A2(_02904_),
    .B1(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__o21ai_1 _09820_ (.A1(net236),
    .A2(_02758_),
    .B1(_02269_),
    .Y(_02907_));
 sky130_fd_sc_hd__a21o_1 _09821_ (.A1(net239),
    .A2(_02907_),
    .B1(_02271_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _09822_ (.A0(_02189_),
    .A1(_02204_),
    .S(net233),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(_02197_),
    .A1(_02220_),
    .S(net234),
    .X(_02910_));
 sky130_fd_sc_hd__or2_1 _09824_ (.A(net237),
    .B(_02909_),
    .X(_02911_));
 sky130_fd_sc_hd__o211a_1 _09825_ (.A1(net238),
    .A2(_02910_),
    .B1(_02911_),
    .C1(net239),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _09826_ (.A0(_02213_),
    .A1(_02235_),
    .S(net233),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(_02768_),
    .A1(_02913_),
    .S(net238),
    .X(_02914_));
 sky130_fd_sc_hd__a21oi_1 _09828_ (.A1(net242),
    .A2(_02914_),
    .B1(_02912_),
    .Y(_02915_));
 sky130_fd_sc_hd__a21o_1 _09829_ (.A1(net244),
    .A2(net216),
    .B1(_02243_),
    .X(_02916_));
 sky130_fd_sc_hd__inv_2 _09830_ (.A(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__or4_2 _09831_ (.A(\div_res[3] ),
    .B(\div_res[2] ),
    .C(\div_res[1] ),
    .D(\div_res[0] ),
    .X(_02918_));
 sky130_fd_sc_hd__a21oi_1 _09832_ (.A1(net165),
    .A2(_02918_),
    .B1(\div_res[4] ),
    .Y(_02919_));
 sky130_fd_sc_hd__a31o_1 _09833_ (.A1(\div_res[4] ),
    .A2(net165),
    .A3(_02918_),
    .B1(net204),
    .X(_02920_));
 sky130_fd_sc_hd__or4_2 _09834_ (.A(\div_shifter[35] ),
    .B(\div_shifter[34] ),
    .C(\div_shifter[33] ),
    .D(\div_shifter[32] ),
    .X(_02921_));
 sky130_fd_sc_hd__and3_1 _09835_ (.A(\div_shifter[36] ),
    .B(net247),
    .C(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__a21oi_1 _09836_ (.A1(net247),
    .A2(_02921_),
    .B1(\div_shifter[36] ),
    .Y(_02923_));
 sky130_fd_sc_hd__or3_2 _09837_ (.A(net250),
    .B(_02922_),
    .C(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__o221a_1 _09838_ (.A1(net239),
    .A2(net215),
    .B1(net206),
    .B2(_06327_),
    .C1(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__o21a_1 _09839_ (.A1(_02761_),
    .A2(_02762_),
    .B1(_02764_),
    .X(_02926_));
 sky130_fd_sc_hd__nor2_1 _09840_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02927_));
 sky130_fd_sc_hd__nand2_1 _09841_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2b_1 _09842_ (.A_N(_02927_),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__xnor2_2 _09843_ (.A(_02926_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__o32a_1 _09844_ (.A1(net244),
    .A2(_06447_),
    .A3(_02930_),
    .B1(net208),
    .B2(_06326_),
    .X(_02931_));
 sky130_fd_sc_hd__o211a_1 _09845_ (.A1(_06328_),
    .A2(net253),
    .B1(_02925_),
    .C1(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__o221a_1 _09846_ (.A1(_02915_),
    .A2(_02917_),
    .B1(_02919_),
    .B2(_02920_),
    .C1(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__o211a_1 _09847_ (.A1(net190),
    .A2(_02908_),
    .B1(_02933_),
    .C1(_02906_),
    .X(_02934_));
 sky130_fd_sc_hd__o21a_1 _09848_ (.A1(_02901_),
    .A2(_02902_),
    .B1(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__a21oi_2 _09849_ (.A1(_02900_),
    .A2(_02935_),
    .B1(_06424_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(curr_PC[4]),
    .B(_02789_),
    .Y(_02937_));
 sky130_fd_sc_hd__or2_1 _09851_ (.A(curr_PC[4]),
    .B(_02789_),
    .X(_02938_));
 sky130_fd_sc_hd__a31o_4 _09852_ (.A1(net267),
    .A2(_02937_),
    .A3(_02938_),
    .B1(_02936_),
    .X(dest_val[4]));
 sky130_fd_sc_hd__nor3_1 _09853_ (.A(_02631_),
    .B(_02740_),
    .C(_02898_),
    .Y(_02939_));
 sky130_fd_sc_hd__or2_1 _09854_ (.A(net157),
    .B(_02939_),
    .X(_02940_));
 sky130_fd_sc_hd__a21oi_4 _09855_ (.A1(_02798_),
    .A2(_02891_),
    .B1(_02890_),
    .Y(_02941_));
 sky130_fd_sc_hd__a21bo_2 _09856_ (.A1(_02880_),
    .A2(_02886_),
    .B1_N(_02888_),
    .X(_02942_));
 sky130_fd_sc_hd__a21oi_4 _09857_ (.A1(_02830_),
    .A2(_02851_),
    .B1(_02850_),
    .Y(_02943_));
 sky130_fd_sc_hd__o22a_1 _09858_ (.A1(net117),
    .A2(net25),
    .B1(net72),
    .B2(net113),
    .X(_02944_));
 sky130_fd_sc_hd__xnor2_1 _09859_ (.A(net105),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__o22a_1 _09860_ (.A1(_06538_),
    .A2(net98),
    .B1(net135),
    .B2(net30),
    .X(_02946_));
 sky130_fd_sc_hd__xnor2_1 _09861_ (.A(net112),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__and2_1 _09862_ (.A(_02945_),
    .B(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__nor2_1 _09863_ (.A(_02945_),
    .B(_02947_),
    .Y(_02949_));
 sky130_fd_sc_hd__nor2_1 _09864_ (.A(_02948_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__o22a_1 _09865_ (.A1(net23),
    .A2(net96),
    .B1(net89),
    .B2(net70),
    .X(_02951_));
 sky130_fd_sc_hd__xor2_1 _09866_ (.A(net108),
    .B(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__xnor2_1 _09867_ (.A(_02950_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_2 _09868_ (.A1(_02816_),
    .A2(_02818_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__or3_1 _09869_ (.A(_02816_),
    .B(_02818_),
    .C(_02953_),
    .X(_02955_));
 sky130_fd_sc_hd__nand2_2 _09870_ (.A(_02954_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__xor2_4 _09871_ (.A(_02943_),
    .B(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__o21ai_4 _09872_ (.A1(_02806_),
    .A2(_02808_),
    .B1(_02804_),
    .Y(_02958_));
 sky130_fd_sc_hd__o22a_2 _09873_ (.A1(net68),
    .A2(net41),
    .B1(net38),
    .B2(net94),
    .X(_02959_));
 sky130_fd_sc_hd__xnor2_4 _09874_ (.A(net100),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__o32a_1 _09875_ (.A1(net123),
    .A2(_00176_),
    .A3(_00177_),
    .B1(net66),
    .B2(net119),
    .X(_02961_));
 sky130_fd_sc_hd__xnor2_2 _09876_ (.A(net102),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__and2_1 _09877_ (.A(_02960_),
    .B(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__xor2_4 _09878_ (.A(_02960_),
    .B(_02962_),
    .X(_02964_));
 sky130_fd_sc_hd__o22a_1 _09879_ (.A1(net21),
    .A2(net85),
    .B1(net80),
    .B2(net65),
    .X(_02965_));
 sky130_fd_sc_hd__xnor2_2 _09880_ (.A(net91),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__xor2_4 _09881_ (.A(_02964_),
    .B(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__a41o_2 _09882_ (.A1(_00140_),
    .A2(_00141_),
    .A3(net35),
    .A4(_02858_),
    .B1(_02857_),
    .X(_02968_));
 sky130_fd_sc_hd__nand2_1 _09883_ (.A(_02967_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__xor2_4 _09884_ (.A(_02967_),
    .B(_02968_),
    .X(_02970_));
 sky130_fd_sc_hd__xor2_4 _09885_ (.A(_02958_),
    .B(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__o21ai_1 _09886_ (.A1(_02822_),
    .A2(_02829_),
    .B1(_02827_),
    .Y(_02972_));
 sky130_fd_sc_hd__a21oi_2 _09887_ (.A1(_02839_),
    .A2(_02841_),
    .B1(_02837_),
    .Y(_02973_));
 sky130_fd_sc_hd__nor2_1 _09888_ (.A(_02847_),
    .B(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__xnor2_1 _09889_ (.A(_02847_),
    .B(_02973_),
    .Y(_02975_));
 sky130_fd_sc_hd__and2b_1 _09890_ (.A_N(_02975_),
    .B(_02972_),
    .X(_02976_));
 sky130_fd_sc_hd__and2b_1 _09891_ (.A_N(_02972_),
    .B(_02975_),
    .X(_02977_));
 sky130_fd_sc_hd__or2_2 _09892_ (.A(_02976_),
    .B(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__o22a_1 _09893_ (.A1(net132),
    .A2(net13),
    .B1(net6),
    .B2(_00283_),
    .X(_02979_));
 sky130_fd_sc_hd__xnor2_2 _09894_ (.A(net194),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__o22a_1 _09895_ (.A1(net57),
    .A2(net130),
    .B1(net128),
    .B2(net18),
    .X(_02981_));
 sky130_fd_sc_hd__xnor2_2 _09896_ (.A(net167),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__or2_1 _09897_ (.A(_00249_),
    .B(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__xnor2_2 _09898_ (.A(_00250_),
    .B(_02982_),
    .Y(_02984_));
 sky130_fd_sc_hd__nand2b_1 _09899_ (.A_N(_02980_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__xnor2_2 _09900_ (.A(_02980_),
    .B(_02984_),
    .Y(_02986_));
 sky130_fd_sc_hd__o22a_1 _09901_ (.A1(net125),
    .A2(net54),
    .B1(net51),
    .B2(net121),
    .X(_02987_));
 sky130_fd_sc_hd__xnor2_1 _09902_ (.A(net152),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__o22a_1 _09903_ (.A1(net62),
    .A2(net88),
    .B1(net83),
    .B2(net59),
    .X(_02989_));
 sky130_fd_sc_hd__xnor2_1 _09904_ (.A(net186),
    .B(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__o22a_1 _09905_ (.A1(net75),
    .A2(net47),
    .B1(net44),
    .B2(net116),
    .X(_02991_));
 sky130_fd_sc_hd__xnor2_1 _09906_ (.A(_06500_),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__nor2_1 _09907_ (.A(_02990_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__xnor2_1 _09908_ (.A(_02990_),
    .B(_02992_),
    .Y(_02994_));
 sky130_fd_sc_hd__nor2_1 _09909_ (.A(_02988_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__and2_1 _09910_ (.A(_02988_),
    .B(_02994_),
    .X(_02996_));
 sky130_fd_sc_hd__nor2_2 _09911_ (.A(_02995_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__xnor2_2 _09912_ (.A(_02868_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__xnor2_1 _09913_ (.A(_02986_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21oi_1 _09914_ (.A1(_00599_),
    .A2(_00600_),
    .B1(_06557_),
    .Y(_03000_));
 sky130_fd_sc_hd__nor2_1 _09915_ (.A(net142),
    .B(net10),
    .Y(_03001_));
 sky130_fd_sc_hd__o21ai_1 _09916_ (.A1(_03000_),
    .A2(_03001_),
    .B1(net33),
    .Y(_03002_));
 sky130_fd_sc_hd__or3_1 _09917_ (.A(net33),
    .B(_03000_),
    .C(_03001_),
    .X(_03003_));
 sky130_fd_sc_hd__or2_1 _09918_ (.A(net148),
    .B(net32),
    .X(_03004_));
 sky130_fd_sc_hd__o32a_1 _09919_ (.A1(net140),
    .A2(_00351_),
    .A3(_00352_),
    .B1(net36),
    .B2(net137),
    .X(_03005_));
 sky130_fd_sc_hd__xnor2_2 _09920_ (.A(_00348_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__and2b_1 _09921_ (.A_N(_03004_),
    .B(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__xnor2_1 _09922_ (.A(_03004_),
    .B(_03006_),
    .Y(_03008_));
 sky130_fd_sc_hd__and3_1 _09923_ (.A(_03002_),
    .B(_03003_),
    .C(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__a21oi_1 _09924_ (.A1(_03002_),
    .A2(_03003_),
    .B1(_03008_),
    .Y(_03010_));
 sky130_fd_sc_hd__or2_1 _09925_ (.A(_03009_),
    .B(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__nor2_1 _09926_ (.A(_02999_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__and2_1 _09927_ (.A(_02999_),
    .B(_03011_),
    .X(_03013_));
 sky130_fd_sc_hd__nor2_2 _09928_ (.A(_03012_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__xnor2_4 _09929_ (.A(_02978_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__and2_1 _09930_ (.A(_02971_),
    .B(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__xor2_4 _09931_ (.A(_02971_),
    .B(_03015_),
    .X(_03017_));
 sky130_fd_sc_hd__xor2_4 _09932_ (.A(_02957_),
    .B(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__a21o_1 _09933_ (.A1(_02813_),
    .A2(_02876_),
    .B1(_02875_),
    .X(_03019_));
 sky130_fd_sc_hd__a21o_1 _09934_ (.A1(_02881_),
    .A2(_02885_),
    .B1(_02884_),
    .X(_03020_));
 sky130_fd_sc_hd__o21ai_4 _09935_ (.A1(_02809_),
    .A2(_02810_),
    .B1(_02812_),
    .Y(_03021_));
 sky130_fd_sc_hd__o21a_2 _09936_ (.A1(_02820_),
    .A2(_02861_),
    .B1(_02860_),
    .X(_03022_));
 sky130_fd_sc_hd__a21boi_4 _09937_ (.A1(_02863_),
    .A2(_02873_),
    .B1_N(_02872_),
    .Y(_03023_));
 sky130_fd_sc_hd__nor2_1 _09938_ (.A(_03022_),
    .B(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__xor2_4 _09939_ (.A(_03022_),
    .B(_03023_),
    .X(_03025_));
 sky130_fd_sc_hd__xor2_2 _09940_ (.A(_03021_),
    .B(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__xnor2_2 _09941_ (.A(_03020_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__nand2b_1 _09942_ (.A_N(_03027_),
    .B(_03019_),
    .Y(_03028_));
 sky130_fd_sc_hd__xnor2_2 _09943_ (.A(_03019_),
    .B(_03027_),
    .Y(_03029_));
 sky130_fd_sc_hd__and2_1 _09944_ (.A(_03018_),
    .B(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__xor2_4 _09945_ (.A(_03018_),
    .B(_03029_),
    .X(_03031_));
 sky130_fd_sc_hd__xnor2_4 _09946_ (.A(_02942_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__or2_1 _09947_ (.A(_02941_),
    .B(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__and2_1 _09948_ (.A(_02941_),
    .B(_03032_),
    .X(_03034_));
 sky130_fd_sc_hd__xnor2_4 _09949_ (.A(_02941_),
    .B(_03032_),
    .Y(_03035_));
 sky130_fd_sc_hd__a21oi_1 _09950_ (.A1(_02733_),
    .A2(_02893_),
    .B1(_02894_),
    .Y(_03036_));
 sky130_fd_sc_hd__a2111oi_2 _09951_ (.A1(_02390_),
    .A2(_02571_),
    .B1(_02572_),
    .C1(_02735_),
    .D1(_02895_),
    .Y(_03037_));
 sky130_fd_sc_hd__nor2_1 _09952_ (.A(_03036_),
    .B(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__or4_1 _09953_ (.A(_02392_),
    .B(_02573_),
    .C(_02735_),
    .D(_02895_),
    .X(_03039_));
 sky130_fd_sc_hd__a21o_1 _09954_ (.A1(_02395_),
    .A2(_02396_),
    .B1(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__a21o_1 _09955_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03035_),
    .X(_03041_));
 sky130_fd_sc_hd__nand3_1 _09956_ (.A(_03035_),
    .B(_03038_),
    .C(_03040_),
    .Y(_03042_));
 sky130_fd_sc_hd__nand2_2 _09957_ (.A(_03041_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__or2_1 _09958_ (.A(_02940_),
    .B(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__a21oi_1 _09959_ (.A1(_02940_),
    .A2(_03043_),
    .B1(net209),
    .Y(_03045_));
 sky130_fd_sc_hd__nor2_1 _09960_ (.A(net157),
    .B(_02079_),
    .Y(_03046_));
 sky130_fd_sc_hd__xnor2_1 _09961_ (.A(_02080_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__o21a_1 _09962_ (.A1(_06326_),
    .A2(_02903_),
    .B1(_06327_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(_06356_),
    .A1(_03048_),
    .S(net304),
    .X(_03049_));
 sky130_fd_sc_hd__xor2_1 _09964_ (.A(_06321_),
    .B(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__o21ai_1 _09965_ (.A1(net236),
    .A2(_02598_),
    .B1(_02269_),
    .Y(_03051_));
 sky130_fd_sc_hd__inv_2 _09966_ (.A(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__a21o_1 _09967_ (.A1(net239),
    .A2(_03051_),
    .B1(_02271_),
    .X(_03053_));
 sky130_fd_sc_hd__inv_2 _09968_ (.A(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(_02406_),
    .A1(_02413_),
    .S(net233),
    .X(_03055_));
 sky130_fd_sc_hd__or2_1 _09970_ (.A(net235),
    .B(_02421_),
    .X(_03056_));
 sky130_fd_sc_hd__o21ai_1 _09971_ (.A1(net234),
    .A2(_02410_),
    .B1(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2_1 _09972_ (.A(net237),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__o211a_1 _09973_ (.A1(net237),
    .A2(_03055_),
    .B1(_03058_),
    .C1(net239),
    .X(_03059_));
 sky130_fd_sc_hd__or2_1 _09974_ (.A(net235),
    .B(_02427_),
    .X(_03060_));
 sky130_fd_sc_hd__o21ai_1 _09975_ (.A1(net233),
    .A2(_02418_),
    .B1(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__or2_1 _09976_ (.A(net238),
    .B(_02583_),
    .X(_03062_));
 sky130_fd_sc_hd__o21ai_1 _09977_ (.A1(net236),
    .A2(_03061_),
    .B1(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__a21o_1 _09978_ (.A1(net240),
    .A2(_03063_),
    .B1(_03059_),
    .X(_03064_));
 sky130_fd_sc_hd__o21ai_1 _09979_ (.A1(\div_res[4] ),
    .A2(_02918_),
    .B1(net165),
    .Y(_03065_));
 sky130_fd_sc_hd__xnor2_1 _09980_ (.A(\div_res[5] ),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__o21a_1 _09981_ (.A1(\div_shifter[36] ),
    .A2(_02921_),
    .B1(net247),
    .X(_03067_));
 sky130_fd_sc_hd__and2_1 _09982_ (.A(\div_shifter[37] ),
    .B(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__nor2_1 _09983_ (.A(\div_shifter[37] ),
    .B(_03067_),
    .Y(_03069_));
 sky130_fd_sc_hd__o32a_1 _09984_ (.A1(net250),
    .A2(_03068_),
    .A3(_03069_),
    .B1(_06460_),
    .B2(_06316_),
    .X(_03070_));
 sky130_fd_sc_hd__o221a_1 _09985_ (.A1(_06319_),
    .A2(net208),
    .B1(_02256_),
    .B2(_06320_),
    .C1(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__o21ai_1 _09986_ (.A1(_06321_),
    .A2(net254),
    .B1(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__o21a_1 _09987_ (.A1(_02926_),
    .A2(_02927_),
    .B1(_02928_),
    .X(_03073_));
 sky130_fd_sc_hd__nor2_1 _09988_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03075_));
 sky130_fd_sc_hd__and2b_1 _09990_ (.A_N(_03074_),
    .B(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__xnor2_1 _09991_ (.A(_03073_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__a31o_1 _09992_ (.A1(net269),
    .A2(net216),
    .A3(_03077_),
    .B1(_03072_),
    .X(_03078_));
 sky130_fd_sc_hd__a221o_1 _09993_ (.A1(_02916_),
    .A2(_03064_),
    .B1(_03066_),
    .B2(_02260_),
    .C1(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__a221o_1 _09994_ (.A1(_02247_),
    .A2(_03050_),
    .B1(_03054_),
    .B2(net192),
    .C1(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__a221o_1 _09995_ (.A1(_03044_),
    .A2(_03045_),
    .B1(_03047_),
    .B2(net252),
    .C1(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__a31o_1 _09996_ (.A1(curr_PC[3]),
    .A2(curr_PC[4]),
    .A3(_02628_),
    .B1(curr_PC[5]),
    .X(_03082_));
 sky130_fd_sc_hd__and3_1 _09997_ (.A(curr_PC[4]),
    .B(curr_PC[5]),
    .C(_02789_),
    .X(_03083_));
 sky130_fd_sc_hd__nor2_1 _09998_ (.A(net262),
    .B(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__a22o_4 _09999_ (.A1(net262),
    .A2(_03081_),
    .B1(_03082_),
    .B2(_03084_),
    .X(dest_val[5]));
 sky130_fd_sc_hd__a21o_1 _10000_ (.A1(_02939_),
    .A2(_03043_),
    .B1(net157),
    .X(_03085_));
 sky130_fd_sc_hd__a21oi_4 _10001_ (.A1(_02942_),
    .A2(_03031_),
    .B1(_03030_),
    .Y(_03086_));
 sky130_fd_sc_hd__a21bo_2 _10002_ (.A1(_03020_),
    .A2(_03026_),
    .B1_N(_03028_),
    .X(_03087_));
 sky130_fd_sc_hd__o211a_1 _10003_ (.A1(_02993_),
    .A2(_02995_),
    .B1(_06556_),
    .C1(net33),
    .X(_03088_));
 sky130_fd_sc_hd__a211oi_1 _10004_ (.A1(_06556_),
    .A2(net35),
    .B1(_02993_),
    .C1(_02995_),
    .Y(_03089_));
 sky130_fd_sc_hd__a211oi_2 _10005_ (.A1(_02983_),
    .A2(_02985_),
    .B1(_03088_),
    .C1(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__o211a_1 _10006_ (.A1(_03088_),
    .A2(_03089_),
    .B1(_02983_),
    .C1(_02985_),
    .X(_03091_));
 sky130_fd_sc_hd__or2_2 _10007_ (.A(_03090_),
    .B(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__o22a_1 _10008_ (.A1(_06492_),
    .A2(net62),
    .B1(net51),
    .B2(net125),
    .X(_03093_));
 sky130_fd_sc_hd__xor2_1 _10009_ (.A(net152),
    .B(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__inv_2 _10010_ (.A(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__o22a_1 _10011_ (.A1(net59),
    .A2(net88),
    .B1(net83),
    .B2(net57),
    .X(_03096_));
 sky130_fd_sc_hd__xnor2_2 _10012_ (.A(net186),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__o22a_1 _10013_ (.A1(net115),
    .A2(net54),
    .B1(net45),
    .B2(net74),
    .X(_03098_));
 sky130_fd_sc_hd__xnor2_2 _10014_ (.A(net149),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__or2_1 _10015_ (.A(_03097_),
    .B(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__xnor2_2 _10016_ (.A(_03097_),
    .B(_03099_),
    .Y(_03101_));
 sky130_fd_sc_hd__or2_1 _10017_ (.A(_03095_),
    .B(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(_03095_),
    .B(_03101_),
    .Y(_03103_));
 sky130_fd_sc_hd__xnor2_1 _10019_ (.A(_03095_),
    .B(_03101_),
    .Y(_03104_));
 sky130_fd_sc_hd__a21o_1 _10020_ (.A1(_02964_),
    .A2(_02966_),
    .B1(_02963_),
    .X(_03105_));
 sky130_fd_sc_hd__xnor2_2 _10021_ (.A(_03104_),
    .B(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__o22a_1 _10022_ (.A1(net18),
    .A2(net130),
    .B1(net128),
    .B2(net13),
    .X(_03107_));
 sky130_fd_sc_hd__xnor2_1 _10023_ (.A(net167),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__nor2_1 _10024_ (.A(_00279_),
    .B(net7),
    .Y(_03109_));
 sky130_fd_sc_hd__o22a_1 _10025_ (.A1(_00278_),
    .A2(net7),
    .B1(_03109_),
    .B2(net195),
    .X(_03110_));
 sky130_fd_sc_hd__and2_1 _10026_ (.A(_03108_),
    .B(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__nor2_1 _10027_ (.A(_03108_),
    .B(_03110_),
    .Y(_03112_));
 sky130_fd_sc_hd__or2_1 _10028_ (.A(_03111_),
    .B(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__xor2_2 _10029_ (.A(_03106_),
    .B(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__o22a_1 _10030_ (.A1(net137),
    .A2(net16),
    .B1(net37),
    .B2(net135),
    .X(_03115_));
 sky130_fd_sc_hd__xnor2_1 _10031_ (.A(_00348_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__inv_2 _10032_ (.A(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__a21oi_1 _10033_ (.A1(_00599_),
    .A2(_00600_),
    .B1(_00171_),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_1 _10034_ (.A(net140),
    .B(net10),
    .Y(_03119_));
 sky130_fd_sc_hd__o21ai_1 _10035_ (.A1(_03118_),
    .A2(_03119_),
    .B1(net33),
    .Y(_03120_));
 sky130_fd_sc_hd__or3_1 _10036_ (.A(net33),
    .B(_03118_),
    .C(_03119_),
    .X(_03121_));
 sky130_fd_sc_hd__o22a_1 _10037_ (.A1(net29),
    .A2(net98),
    .B1(net96),
    .B2(net27),
    .X(_03122_));
 sky130_fd_sc_hd__xnor2_1 _10038_ (.A(net112),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__and3_1 _10039_ (.A(_03120_),
    .B(_03121_),
    .C(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__nand3_1 _10040_ (.A(_03120_),
    .B(_03121_),
    .C(_03123_),
    .Y(_03125_));
 sky130_fd_sc_hd__a21oi_1 _10041_ (.A1(_03120_),
    .A2(_03121_),
    .B1(_03123_),
    .Y(_03126_));
 sky130_fd_sc_hd__or3_1 _10042_ (.A(_03117_),
    .B(_03124_),
    .C(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__o21ai_1 _10043_ (.A1(_03124_),
    .A2(_03126_),
    .B1(_03117_),
    .Y(_03128_));
 sky130_fd_sc_hd__and2_1 _10044_ (.A(_03127_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__nand2_1 _10045_ (.A(_03114_),
    .B(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__xnor2_2 _10046_ (.A(_03114_),
    .B(_03129_),
    .Y(_03131_));
 sky130_fd_sc_hd__xor2_1 _10047_ (.A(_03092_),
    .B(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__o21ba_1 _10048_ (.A1(_02949_),
    .A2(_02952_),
    .B1_N(_02948_),
    .X(_03133_));
 sky130_fd_sc_hd__o22a_1 _10049_ (.A1(net94),
    .A2(net48),
    .B1(net39),
    .B2(net68),
    .X(_03134_));
 sky130_fd_sc_hd__xnor2_1 _10050_ (.A(net100),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__o22a_1 _10051_ (.A1(net20),
    .A2(net80),
    .B1(net41),
    .B2(net64),
    .X(_03136_));
 sky130_fd_sc_hd__xnor2_1 _10052_ (.A(net92),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__and2_1 _10053_ (.A(_03135_),
    .B(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__xor2_1 _10054_ (.A(_03135_),
    .B(_03137_),
    .X(_03139_));
 sky130_fd_sc_hd__o21ai_1 _10055_ (.A1(_03007_),
    .A2(_03009_),
    .B1(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__or3_1 _10056_ (.A(_03007_),
    .B(_03009_),
    .C(_03139_),
    .X(_03141_));
 sky130_fd_sc_hd__and2_1 _10057_ (.A(_03140_),
    .B(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__nand2b_1 _10058_ (.A_N(_03133_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__xnor2_1 _10059_ (.A(_03133_),
    .B(_03142_),
    .Y(_03144_));
 sky130_fd_sc_hd__and2_1 _10060_ (.A(_03132_),
    .B(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(_03132_),
    .B(_03144_),
    .Y(_03146_));
 sky130_fd_sc_hd__nor2_2 _10062_ (.A(_03145_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__a32oi_4 _10063_ (.A1(_02865_),
    .A2(_02867_),
    .A3(_02997_),
    .B1(_02998_),
    .B2(_02986_),
    .Y(_03148_));
 sky130_fd_sc_hd__o22a_1 _10064_ (.A1(net117),
    .A2(net70),
    .B1(net89),
    .B2(net24),
    .X(_03149_));
 sky130_fd_sc_hd__xnor2_1 _10065_ (.A(net108),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__o22a_1 _10066_ (.A1(net119),
    .A2(_00178_),
    .B1(net66),
    .B2(net85),
    .X(_03151_));
 sky130_fd_sc_hd__xnor2_1 _10067_ (.A(net102),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__and2_1 _10068_ (.A(_03150_),
    .B(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__nor2_1 _10069_ (.A(_03150_),
    .B(_03152_),
    .Y(_03154_));
 sky130_fd_sc_hd__nor2_1 _10070_ (.A(_03153_),
    .B(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__o22a_1 _10071_ (.A1(net113),
    .A2(net25),
    .B1(net72),
    .B2(net123),
    .X(_03156_));
 sky130_fd_sc_hd__xor2_2 _10072_ (.A(net105),
    .B(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__xnor2_2 _10073_ (.A(_03155_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__o21a_1 _10074_ (.A1(_02974_),
    .A2(_02976_),
    .B1(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__o21ai_1 _10075_ (.A1(_02974_),
    .A2(_02976_),
    .B1(_03158_),
    .Y(_03160_));
 sky130_fd_sc_hd__nor3_2 _10076_ (.A(_02974_),
    .B(_02976_),
    .C(_03158_),
    .Y(_03161_));
 sky130_fd_sc_hd__nor2_2 _10077_ (.A(_03159_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__xnor2_4 _10078_ (.A(_03148_),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__xor2_4 _10079_ (.A(_03147_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__a21o_1 _10080_ (.A1(_02957_),
    .A2(_03017_),
    .B1(_03016_),
    .X(_03165_));
 sky130_fd_sc_hd__o21ai_2 _10081_ (.A1(_02943_),
    .A2(_02956_),
    .B1(_02954_),
    .Y(_03166_));
 sky130_fd_sc_hd__a21boi_2 _10082_ (.A1(_02958_),
    .A2(_02970_),
    .B1_N(_02969_),
    .Y(_03167_));
 sky130_fd_sc_hd__o21ba_1 _10083_ (.A1(_02978_),
    .A2(_03013_),
    .B1_N(_03012_),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_1 _10084_ (.A(_03167_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__xor2_2 _10085_ (.A(_03167_),
    .B(_03168_),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_2 _10086_ (.A(_03166_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__a21oi_4 _10087_ (.A1(_03021_),
    .A2(_03025_),
    .B1(_03024_),
    .Y(_03172_));
 sky130_fd_sc_hd__xnor2_2 _10088_ (.A(_03171_),
    .B(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__and2b_1 _10089_ (.A_N(_03173_),
    .B(_03165_),
    .X(_03174_));
 sky130_fd_sc_hd__xnor2_2 _10090_ (.A(_03165_),
    .B(_03173_),
    .Y(_03175_));
 sky130_fd_sc_hd__and2_1 _10091_ (.A(_03164_),
    .B(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__xor2_4 _10092_ (.A(_03164_),
    .B(_03175_),
    .X(_03177_));
 sky130_fd_sc_hd__xnor2_4 _10093_ (.A(_03087_),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__or2_1 _10094_ (.A(_03086_),
    .B(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__and2_1 _10095_ (.A(_03086_),
    .B(_03178_),
    .X(_03180_));
 sky130_fd_sc_hd__xnor2_4 _10096_ (.A(_03086_),
    .B(_03178_),
    .Y(_03181_));
 sky130_fd_sc_hd__or3_2 _10097_ (.A(_02792_),
    .B(_02895_),
    .C(_03035_),
    .X(_03182_));
 sky130_fd_sc_hd__a21oi_2 _10098_ (.A1(_02893_),
    .A2(_03033_),
    .B1(_03034_),
    .Y(_03183_));
 sky130_fd_sc_hd__a2111oi_2 _10099_ (.A1(_02571_),
    .A2(_02733_),
    .B1(_02734_),
    .C1(_02895_),
    .D1(_03035_),
    .Y(_03184_));
 sky130_fd_sc_hd__nor2_1 _10100_ (.A(_03183_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__o21a_1 _10101_ (.A1(_02577_),
    .A2(_03182_),
    .B1(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__xnor2_4 _10102_ (.A(_03181_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__o21ai_1 _10103_ (.A1(_03085_),
    .A2(_03187_),
    .B1(_02171_),
    .Y(_03188_));
 sky130_fd_sc_hd__a21oi_1 _10104_ (.A1(_03085_),
    .A2(_03187_),
    .B1(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__nor2_1 _10105_ (.A(net157),
    .B(_02081_),
    .Y(_03190_));
 sky130_fd_sc_hd__xnor2_1 _10106_ (.A(_02082_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__o21ai_1 _10107_ (.A1(_06319_),
    .A2(_03048_),
    .B1(_06320_),
    .Y(_03192_));
 sky130_fd_sc_hd__mux2_1 _10108_ (.A0(_06357_),
    .A1(_03192_),
    .S(net304),
    .X(_03193_));
 sky130_fd_sc_hd__nand2_1 _10109_ (.A(_06313_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__o21a_1 _10110_ (.A1(_06313_),
    .A2(_03193_),
    .B1(_02247_),
    .X(_03195_));
 sky130_fd_sc_hd__o21a_1 _10111_ (.A1(net236),
    .A2(_02428_),
    .B1(_02269_),
    .X(_03196_));
 sky130_fd_sc_hd__o21ai_2 _10112_ (.A1(net240),
    .A2(_03196_),
    .B1(_02272_),
    .Y(_03197_));
 sky130_fd_sc_hd__nor2_1 _10113_ (.A(net190),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(_02588_),
    .A1(_02591_),
    .S(net233),
    .X(_03199_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(_02590_),
    .A1(_02595_),
    .S(net233),
    .X(_03200_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(_03199_),
    .A1(_03200_),
    .S(net236),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(_02594_),
    .A1(_02597_),
    .S(net233),
    .X(_03202_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(_02457_),
    .A1(_03202_),
    .S(net238),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _10119_ (.A0(_03201_),
    .A1(_03203_),
    .S(net240),
    .X(_03204_));
 sky130_fd_sc_hd__or3_1 _10120_ (.A(\div_res[5] ),
    .B(\div_res[4] ),
    .C(_02918_),
    .X(_03205_));
 sky130_fd_sc_hd__a21oi_1 _10121_ (.A1(net165),
    .A2(_03205_),
    .B1(\div_res[6] ),
    .Y(_03206_));
 sky130_fd_sc_hd__a31o_1 _10122_ (.A1(\div_res[6] ),
    .A2(net165),
    .A3(_03205_),
    .B1(net205),
    .X(_03207_));
 sky130_fd_sc_hd__nor2_1 _10123_ (.A(_03206_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__or3_2 _10124_ (.A(\div_shifter[37] ),
    .B(\div_shifter[36] ),
    .C(_02921_),
    .X(_03209_));
 sky130_fd_sc_hd__a21oi_1 _10125_ (.A1(net249),
    .A2(_03209_),
    .B1(\div_shifter[38] ),
    .Y(_03210_));
 sky130_fd_sc_hd__a311oi_4 _10126_ (.A1(\div_shifter[38] ),
    .A2(net249),
    .A3(_03209_),
    .B1(_03210_),
    .C1(net250),
    .Y(_03211_));
 sky130_fd_sc_hd__a221o_1 _10127_ (.A1(_06307_),
    .A2(_06459_),
    .B1(_02255_),
    .B2(_06312_),
    .C1(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__a221o_1 _10128_ (.A1(_06311_),
    .A2(_02245_),
    .B1(_02249_),
    .B2(_06313_),
    .C1(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__o21a_1 _10129_ (.A1(_03073_),
    .A2(_03074_),
    .B1(_03075_),
    .X(_03214_));
 sky130_fd_sc_hd__nor2_1 _10130_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03215_));
 sky130_fd_sc_hd__nand2_1 _10131_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03216_));
 sky130_fd_sc_hd__and2b_1 _10132_ (.A_N(_03215_),
    .B(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__xnor2_1 _10133_ (.A(_03214_),
    .B(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__a311o_1 _10134_ (.A1(net268),
    .A2(net216),
    .A3(_03218_),
    .B1(_03213_),
    .C1(_03208_),
    .X(_03219_));
 sky130_fd_sc_hd__a211o_1 _10135_ (.A1(_02916_),
    .A2(_03204_),
    .B1(_03219_),
    .C1(_03198_),
    .X(_03220_));
 sky130_fd_sc_hd__a21o_1 _10136_ (.A1(_03194_),
    .A2(_03195_),
    .B1(_03220_),
    .X(_03221_));
 sky130_fd_sc_hd__a211o_1 _10137_ (.A1(net252),
    .A2(_03191_),
    .B1(_03221_),
    .C1(_03189_),
    .X(_03222_));
 sky130_fd_sc_hd__and2_1 _10138_ (.A(curr_PC[6]),
    .B(_03083_),
    .X(_03223_));
 sky130_fd_sc_hd__o21ai_1 _10139_ (.A1(curr_PC[6]),
    .A2(_03083_),
    .B1(net267),
    .Y(_03224_));
 sky130_fd_sc_hd__a2bb2o_4 _10140_ (.A1_N(_03223_),
    .A2_N(_03224_),
    .B1(net262),
    .B2(_03222_),
    .X(dest_val[6]));
 sky130_fd_sc_hd__a31o_1 _10141_ (.A1(_02939_),
    .A2(_03043_),
    .A3(_03187_),
    .B1(net158),
    .X(_03225_));
 sky130_fd_sc_hd__a21oi_4 _10142_ (.A1(_03087_),
    .A2(_03177_),
    .B1(_03176_),
    .Y(_03226_));
 sky130_fd_sc_hd__o21bai_4 _10143_ (.A1(_03171_),
    .A2(_03172_),
    .B1_N(_03174_),
    .Y(_03227_));
 sky130_fd_sc_hd__o22a_1 _10144_ (.A1(net137),
    .A2(net10),
    .B1(net5),
    .B2(net140),
    .X(_03228_));
 sky130_fd_sc_hd__xnor2_1 _10145_ (.A(net33),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2b_1 _10146_ (.A_N(_03111_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__xor2_1 _10147_ (.A(_03111_),
    .B(_03229_),
    .X(_03231_));
 sky130_fd_sc_hd__or2_1 _10148_ (.A(_00171_),
    .B(net32),
    .X(_03232_));
 sky130_fd_sc_hd__xnor2_1 _10149_ (.A(_03231_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__o22a_1 _10150_ (.A1(net135),
    .A2(net15),
    .B1(net37),
    .B2(net98),
    .X(_03234_));
 sky130_fd_sc_hd__xnor2_1 _10151_ (.A(net77),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__o22a_1 _10152_ (.A1(net117),
    .A2(net23),
    .B1(net70),
    .B2(net113),
    .X(_03236_));
 sky130_fd_sc_hd__xnor2_1 _10153_ (.A(net108),
    .B(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__nand2b_1 _10154_ (.A_N(_03235_),
    .B(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__xor2_1 _10155_ (.A(_03235_),
    .B(_03237_),
    .X(_03239_));
 sky130_fd_sc_hd__o22a_1 _10156_ (.A1(net29),
    .A2(net96),
    .B1(net89),
    .B2(net28),
    .X(_03240_));
 sky130_fd_sc_hd__xnor2_1 _10157_ (.A(net112),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__inv_2 _10158_ (.A(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__xnor2_1 _10159_ (.A(_03239_),
    .B(_03241_),
    .Y(_03243_));
 sky130_fd_sc_hd__o21ai_1 _10160_ (.A1(_03095_),
    .A2(_03101_),
    .B1(_03100_),
    .Y(_03244_));
 sky130_fd_sc_hd__or2_1 _10161_ (.A(net57),
    .B(net88),
    .X(_03245_));
 sky130_fd_sc_hd__a21o_1 _10162_ (.A1(_00243_),
    .A2(_00244_),
    .B1(net83),
    .X(_03246_));
 sky130_fd_sc_hd__a21o_1 _10163_ (.A1(_03245_),
    .A2(_03246_),
    .B1(net186),
    .X(_03247_));
 sky130_fd_sc_hd__nand3_1 _10164_ (.A(net186),
    .B(_03245_),
    .C(_03246_),
    .Y(_03248_));
 sky130_fd_sc_hd__nand3_1 _10165_ (.A(net194),
    .B(_03247_),
    .C(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__a21o_1 _10166_ (.A1(_03247_),
    .A2(_03248_),
    .B1(net194),
    .X(_03250_));
 sky130_fd_sc_hd__o22a_1 _10167_ (.A1(net130),
    .A2(net13),
    .B1(net6),
    .B2(_00313_),
    .X(_03251_));
 sky130_fd_sc_hd__xor2_1 _10168_ (.A(net167),
    .B(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__nand3_1 _10169_ (.A(_03249_),
    .B(_03250_),
    .C(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__a21o_1 _10170_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_03252_),
    .X(_03254_));
 sky130_fd_sc_hd__and3_1 _10171_ (.A(_03244_),
    .B(_03253_),
    .C(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__nand3_1 _10172_ (.A(_03244_),
    .B(_03253_),
    .C(_03254_),
    .Y(_03256_));
 sky130_fd_sc_hd__a21o_1 _10173_ (.A1(_03253_),
    .A2(_03254_),
    .B1(_03244_),
    .X(_03257_));
 sky130_fd_sc_hd__and3_1 _10174_ (.A(_03138_),
    .B(_03256_),
    .C(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__a21oi_1 _10175_ (.A1(_03256_),
    .A2(_03257_),
    .B1(_03138_),
    .Y(_03259_));
 sky130_fd_sc_hd__nor3b_1 _10176_ (.A(_03258_),
    .B(_03259_),
    .C_N(_03243_),
    .Y(_03260_));
 sky130_fd_sc_hd__o21ba_1 _10177_ (.A1(_03258_),
    .A2(_03259_),
    .B1_N(_03243_),
    .X(_03261_));
 sky130_fd_sc_hd__or3_1 _10178_ (.A(_03233_),
    .B(_03260_),
    .C(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__o21ai_1 _10179_ (.A1(_03260_),
    .A2(_03261_),
    .B1(_03233_),
    .Y(_03263_));
 sky130_fd_sc_hd__o21ba_1 _10180_ (.A1(_03154_),
    .A2(_03157_),
    .B1_N(_03153_),
    .X(_03264_));
 sky130_fd_sc_hd__o22a_1 _10181_ (.A1(net125),
    .A2(net62),
    .B1(net59),
    .B2(net121),
    .X(_03265_));
 sky130_fd_sc_hd__xnor2_1 _10182_ (.A(net152),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__o22a_1 _10183_ (.A1(net68),
    .A2(net48),
    .B1(net45),
    .B2(net94),
    .X(_03267_));
 sky130_fd_sc_hd__xnor2_1 _10184_ (.A(_00153_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__nor2_1 _10185_ (.A(_03266_),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__and2_1 _10186_ (.A(_03266_),
    .B(_03268_),
    .X(_03270_));
 sky130_fd_sc_hd__or2_1 _10187_ (.A(_03269_),
    .B(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__o22a_1 _10188_ (.A1(net74),
    .A2(net54),
    .B1(net51),
    .B2(net115),
    .X(_03272_));
 sky130_fd_sc_hd__xnor2_1 _10189_ (.A(net149),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__xnor2_1 _10190_ (.A(_03271_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21oi_1 _10191_ (.A1(_03125_),
    .A2(_03127_),
    .B1(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__and3_1 _10192_ (.A(_03125_),
    .B(_03127_),
    .C(_03274_),
    .X(_03276_));
 sky130_fd_sc_hd__or2_1 _10193_ (.A(_03275_),
    .B(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__xor2_1 _10194_ (.A(_03264_),
    .B(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__and3_1 _10195_ (.A(_03262_),
    .B(_03263_),
    .C(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__a21oi_1 _10196_ (.A1(_03262_),
    .A2(_03263_),
    .B1(_03278_),
    .Y(_03280_));
 sky130_fd_sc_hd__nor2_2 _10197_ (.A(_03279_),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__a32o_2 _10198_ (.A1(_03102_),
    .A2(_03103_),
    .A3(_03105_),
    .B1(_03106_),
    .B2(_03113_),
    .X(_03282_));
 sky130_fd_sc_hd__o22a_1 _10199_ (.A1(net123),
    .A2(net25),
    .B1(net72),
    .B2(net119),
    .X(_03283_));
 sky130_fd_sc_hd__xnor2_1 _10200_ (.A(net105),
    .B(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__o22a_1 _10201_ (.A1(net20),
    .A2(net42),
    .B1(net39),
    .B2(net64),
    .X(_03285_));
 sky130_fd_sc_hd__xnor2_1 _10202_ (.A(net91),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__and2_1 _10203_ (.A(_03284_),
    .B(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(_03284_),
    .B(_03286_),
    .Y(_03288_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(_03284_),
    .B(_03286_),
    .Y(_03289_));
 sky130_fd_sc_hd__nor2_1 _10206_ (.A(_03287_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__o22a_1 _10207_ (.A1(_00178_),
    .A2(net84),
    .B1(net80),
    .B2(net66),
    .X(_03291_));
 sky130_fd_sc_hd__xor2_1 _10208_ (.A(net103),
    .B(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__xnor2_1 _10209_ (.A(_03290_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__o21a_1 _10210_ (.A1(_03088_),
    .A2(_03090_),
    .B1(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__or3_1 _10211_ (.A(_03088_),
    .B(_03090_),
    .C(_03293_),
    .X(_03295_));
 sky130_fd_sc_hd__and2b_1 _10212_ (.A_N(_03294_),
    .B(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__xnor2_4 _10213_ (.A(_03282_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__xnor2_4 _10214_ (.A(_03281_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__a21o_2 _10215_ (.A1(_03147_),
    .A2(_03163_),
    .B1(_03145_),
    .X(_03299_));
 sky130_fd_sc_hd__o21ai_4 _10216_ (.A1(_03148_),
    .A2(_03161_),
    .B1(_03160_),
    .Y(_03300_));
 sky130_fd_sc_hd__o21ai_4 _10217_ (.A1(_03092_),
    .A2(_03131_),
    .B1(_03130_),
    .Y(_03301_));
 sky130_fd_sc_hd__and2_1 _10218_ (.A(_03140_),
    .B(_03143_),
    .X(_03302_));
 sky130_fd_sc_hd__a21bo_1 _10219_ (.A1(_03140_),
    .A2(_03143_),
    .B1_N(_03301_),
    .X(_03303_));
 sky130_fd_sc_hd__xnor2_4 _10220_ (.A(_03301_),
    .B(_03302_),
    .Y(_03304_));
 sky130_fd_sc_hd__xnor2_4 _10221_ (.A(_03300_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__a21oi_2 _10222_ (.A1(_03166_),
    .A2(_03170_),
    .B1(_03169_),
    .Y(_03306_));
 sky130_fd_sc_hd__nor2_1 _10223_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__xor2_4 _10224_ (.A(_03305_),
    .B(_03306_),
    .X(_03308_));
 sky130_fd_sc_hd__xor2_4 _10225_ (.A(_03299_),
    .B(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__and2_1 _10226_ (.A(_03298_),
    .B(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__xor2_4 _10227_ (.A(_03298_),
    .B(_03309_),
    .X(_03311_));
 sky130_fd_sc_hd__xnor2_4 _10228_ (.A(_03227_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__or2_1 _10229_ (.A(_03226_),
    .B(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__and2_1 _10230_ (.A(_03226_),
    .B(_03312_),
    .X(_03314_));
 sky130_fd_sc_hd__xnor2_4 _10231_ (.A(_03226_),
    .B(_03312_),
    .Y(_03315_));
 sky130_fd_sc_hd__or4_1 _10232_ (.A(_02735_),
    .B(_02895_),
    .C(_03035_),
    .D(_03181_),
    .X(_03316_));
 sky130_fd_sc_hd__a21o_1 _10233_ (.A1(_03033_),
    .A2(_03179_),
    .B1(_03180_),
    .X(_03317_));
 sky130_fd_sc_hd__a2111o_1 _10234_ (.A1(_02733_),
    .A2(_02893_),
    .B1(_02894_),
    .C1(_03035_),
    .D1(_03181_),
    .X(_03318_));
 sky130_fd_sc_hd__o211a_1 _10235_ (.A1(_02739_),
    .A2(_03316_),
    .B1(_03317_),
    .C1(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__xnor2_4 _10236_ (.A(_03315_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__a21oi_1 _10237_ (.A1(_03225_),
    .A2(_03320_),
    .B1(net209),
    .Y(_03321_));
 sky130_fd_sc_hd__o21a_1 _10238_ (.A1(_03225_),
    .A2(_03320_),
    .B1(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__a21oi_1 _10239_ (.A1(net161),
    .A2(_02083_),
    .B1(_02084_),
    .Y(_03323_));
 sky130_fd_sc_hd__a311oi_1 _10240_ (.A1(net161),
    .A2(_02083_),
    .A3(_02084_),
    .B1(_02254_),
    .C1(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__a21oi_1 _10241_ (.A1(_06311_),
    .A2(_03192_),
    .B1(_06312_),
    .Y(_03325_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(_06358_),
    .A1(_03325_),
    .S(net304),
    .X(_03326_));
 sky130_fd_sc_hd__a21oi_1 _10243_ (.A1(_06291_),
    .A2(_03326_),
    .B1(net255),
    .Y(_03327_));
 sky130_fd_sc_hd__o21a_1 _10244_ (.A1(_06291_),
    .A2(_03326_),
    .B1(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__o21a_1 _10245_ (.A1(net236),
    .A2(_02236_),
    .B1(_02269_),
    .X(_03329_));
 sky130_fd_sc_hd__o21a_1 _10246_ (.A1(net241),
    .A2(_03329_),
    .B1(_02272_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _10247_ (.A0(_02748_),
    .A1(_02751_),
    .S(net233),
    .X(_03331_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(_02750_),
    .A1(_02755_),
    .S(net234),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(_03331_),
    .A1(_03332_),
    .S(net237),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(_02754_),
    .A1(_02757_),
    .S(net233),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(_02267_),
    .A1(_03334_),
    .S(net238),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _10252_ (.A0(_03333_),
    .A1(_03335_),
    .S(net241),
    .X(_03336_));
 sky130_fd_sc_hd__or2_1 _10253_ (.A(\div_res[6] ),
    .B(_03205_),
    .X(_03337_));
 sky130_fd_sc_hd__a21oi_1 _10254_ (.A1(net165),
    .A2(_03337_),
    .B1(\div_res[7] ),
    .Y(_03338_));
 sky130_fd_sc_hd__a31o_1 _10255_ (.A1(\div_res[7] ),
    .A2(net165),
    .A3(_03337_),
    .B1(net205),
    .X(_03339_));
 sky130_fd_sc_hd__or2_1 _10256_ (.A(\div_shifter[38] ),
    .B(_03209_),
    .X(_03340_));
 sky130_fd_sc_hd__a21oi_2 _10257_ (.A1(net247),
    .A2(_03340_),
    .B1(\div_shifter[39] ),
    .Y(_03341_));
 sky130_fd_sc_hd__a31o_1 _10258_ (.A1(\div_shifter[39] ),
    .A2(net247),
    .A3(_03340_),
    .B1(net250),
    .X(_03342_));
 sky130_fd_sc_hd__o2bb2a_1 _10259_ (.A1_N(_06256_),
    .A2_N(_06459_),
    .B1(net208),
    .B2(_06274_),
    .X(_03343_));
 sky130_fd_sc_hd__o22a_1 _10260_ (.A1(_06282_),
    .A2(_02256_),
    .B1(_03341_),
    .B2(_03342_),
    .X(_03344_));
 sky130_fd_sc_hd__o211a_1 _10261_ (.A1(_06291_),
    .A2(net254),
    .B1(_03343_),
    .C1(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__o21ai_1 _10262_ (.A1(_03338_),
    .A2(_03339_),
    .B1(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__o21a_1 _10263_ (.A1(_03214_),
    .A2(_03215_),
    .B1(_03216_),
    .X(_03347_));
 sky130_fd_sc_hd__nor2_1 _10264_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03348_));
 sky130_fd_sc_hd__nand2_1 _10265_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03349_));
 sky130_fd_sc_hd__and2b_1 _10266_ (.A_N(_03348_),
    .B(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__xnor2_1 _10267_ (.A(_03347_),
    .B(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__a31o_1 _10268_ (.A1(net268),
    .A2(net216),
    .A3(_03351_),
    .B1(_03346_),
    .X(_03352_));
 sky130_fd_sc_hd__a221o_1 _10269_ (.A1(net192),
    .A2(_03330_),
    .B1(_03336_),
    .B2(_02916_),
    .C1(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__or4_2 _10270_ (.A(_03322_),
    .B(_03324_),
    .C(_03328_),
    .D(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__or2_1 _10271_ (.A(curr_PC[7]),
    .B(_03223_),
    .X(_03355_));
 sky130_fd_sc_hd__a21oi_1 _10272_ (.A1(curr_PC[7]),
    .A2(_03223_),
    .B1(net262),
    .Y(_03356_));
 sky130_fd_sc_hd__a22o_4 _10273_ (.A1(net262),
    .A2(_03354_),
    .B1(_03355_),
    .B2(_03356_),
    .X(dest_val[7]));
 sky130_fd_sc_hd__a221oi_2 _10274_ (.A1(_02896_),
    .A2(_02897_),
    .B1(_03041_),
    .B2(_03042_),
    .C1(_02740_),
    .Y(_03357_));
 sky130_fd_sc_hd__nand4_2 _10275_ (.A(_02630_),
    .B(_03187_),
    .C(_03320_),
    .D(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__or2_1 _10276_ (.A(_02168_),
    .B(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__a21o_2 _10277_ (.A1(_03227_),
    .A2(_03311_),
    .B1(_03310_),
    .X(_03360_));
 sky130_fd_sc_hd__a21o_2 _10278_ (.A1(_03299_),
    .A2(_03308_),
    .B1(_03307_),
    .X(_03361_));
 sky130_fd_sc_hd__o22a_1 _10279_ (.A1(net94),
    .A2(net54),
    .B1(net45),
    .B2(net68),
    .X(_03362_));
 sky130_fd_sc_hd__xnor2_1 _10280_ (.A(net100),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__o22a_1 _10281_ (.A1(_00178_),
    .A2(net80),
    .B1(net42),
    .B2(net66),
    .X(_03364_));
 sky130_fd_sc_hd__xnor2_1 _10282_ (.A(net102),
    .B(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__and2_1 _10283_ (.A(_03363_),
    .B(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__nor2_1 _10284_ (.A(_03363_),
    .B(_03365_),
    .Y(_03367_));
 sky130_fd_sc_hd__nor2_1 _10285_ (.A(_03366_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__o22a_1 _10286_ (.A1(net64),
    .A2(net48),
    .B1(net39),
    .B2(net20),
    .X(_03369_));
 sky130_fd_sc_hd__xnor2_2 _10287_ (.A(net91),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__xnor2_2 _10288_ (.A(_03368_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__o21a_1 _10289_ (.A1(_03231_),
    .A2(_03232_),
    .B1(_03230_),
    .X(_03372_));
 sky130_fd_sc_hd__xor2_1 _10290_ (.A(_03371_),
    .B(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__o21ai_1 _10291_ (.A1(_03255_),
    .A2(_03258_),
    .B1(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__or3_1 _10292_ (.A(_03255_),
    .B(_03258_),
    .C(_03373_),
    .X(_03375_));
 sky130_fd_sc_hd__and2_2 _10293_ (.A(_03374_),
    .B(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__o21ai_1 _10294_ (.A1(_03289_),
    .A2(_03292_),
    .B1(_03288_),
    .Y(_03377_));
 sky130_fd_sc_hd__o22a_1 _10295_ (.A1(net125),
    .A2(net59),
    .B1(net57),
    .B2(net121),
    .X(_03378_));
 sky130_fd_sc_hd__xnor2_1 _10296_ (.A(net152),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__o22a_1 _10297_ (.A1(net115),
    .A2(net62),
    .B1(net51),
    .B2(net74),
    .X(_03380_));
 sky130_fd_sc_hd__xnor2_1 _10298_ (.A(net149),
    .B(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__xnor2_1 _10299_ (.A(_03379_),
    .B(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__o21a_1 _10300_ (.A1(_03239_),
    .A2(_03242_),
    .B1(_03238_),
    .X(_03383_));
 sky130_fd_sc_hd__nor2_1 _10301_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_1 _10302_ (.A(_03382_),
    .B(_03383_),
    .Y(_03385_));
 sky130_fd_sc_hd__and2b_1 _10303_ (.A_N(_03385_),
    .B(_03377_),
    .X(_03386_));
 sky130_fd_sc_hd__and2b_1 _10304_ (.A_N(_03377_),
    .B(_03385_),
    .X(_03387_));
 sky130_fd_sc_hd__nor2_1 _10305_ (.A(_03386_),
    .B(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__o22a_1 _10306_ (.A1(net135),
    .A2(net9),
    .B1(net5),
    .B2(net137),
    .X(_03389_));
 sky130_fd_sc_hd__xnor2_1 _10307_ (.A(net33),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__o22a_1 _10308_ (.A1(net98),
    .A2(net16),
    .B1(net37),
    .B2(net96),
    .X(_03391_));
 sky130_fd_sc_hd__xnor2_1 _10309_ (.A(net77),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__or2_1 _10310_ (.A(net140),
    .B(net32),
    .X(_03393_));
 sky130_fd_sc_hd__nor2_1 _10311_ (.A(_03392_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__xor2_1 _10312_ (.A(_03392_),
    .B(_03393_),
    .X(_03395_));
 sky130_fd_sc_hd__and2_1 _10313_ (.A(_03390_),
    .B(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__nor2_1 _10314_ (.A(_03390_),
    .B(_03395_),
    .Y(_03397_));
 sky130_fd_sc_hd__or2_1 _10315_ (.A(_03396_),
    .B(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__o21ba_1 _10316_ (.A1(_03271_),
    .A2(_03273_),
    .B1_N(_03269_),
    .X(_03399_));
 sky130_fd_sc_hd__a21boi_1 _10317_ (.A1(_03250_),
    .A2(_03252_),
    .B1_N(_03249_),
    .Y(_03400_));
 sky130_fd_sc_hd__o22a_1 _10318_ (.A1(net18),
    .A2(net88),
    .B1(net83),
    .B2(net13),
    .X(_03401_));
 sky130_fd_sc_hd__xnor2_1 _10319_ (.A(_06470_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__or2_1 _10320_ (.A(_00308_),
    .B(net7),
    .X(_03403_));
 sky130_fd_sc_hd__nor2_1 _10321_ (.A(_00307_),
    .B(net7),
    .Y(_03404_));
 sky130_fd_sc_hd__mux2_2 _10322_ (.A0(_03403_),
    .A1(_03404_),
    .S(net167),
    .X(_03405_));
 sky130_fd_sc_hd__or2_1 _10323_ (.A(_03402_),
    .B(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__xnor2_1 _10324_ (.A(_03402_),
    .B(_03405_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2b_1 _10325_ (.A_N(_03400_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__xnor2_1 _10326_ (.A(_03400_),
    .B(_03407_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2b_1 _10327_ (.A_N(_03399_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__xnor2_1 _10328_ (.A(_03399_),
    .B(_03409_),
    .Y(_03411_));
 sky130_fd_sc_hd__o22a_1 _10329_ (.A1(net119),
    .A2(net25),
    .B1(net72),
    .B2(net84),
    .X(_03412_));
 sky130_fd_sc_hd__xor2_1 _10330_ (.A(net105),
    .B(_03412_),
    .X(_03413_));
 sky130_fd_sc_hd__o22a_1 _10331_ (.A1(net117),
    .A2(net28),
    .B1(net89),
    .B2(net29),
    .X(_03414_));
 sky130_fd_sc_hd__xnor2_1 _10332_ (.A(_06524_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nor2_1 _10333_ (.A(_03413_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__xor2_1 _10334_ (.A(_03413_),
    .B(_03415_),
    .X(_03417_));
 sky130_fd_sc_hd__o22a_1 _10335_ (.A1(net113),
    .A2(net23),
    .B1(net70),
    .B2(net123),
    .X(_03418_));
 sky130_fd_sc_hd__xnor2_1 _10336_ (.A(net108),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__and2_1 _10337_ (.A(_03417_),
    .B(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__nor2_1 _10338_ (.A(_03417_),
    .B(_03419_),
    .Y(_03421_));
 sky130_fd_sc_hd__nor2_1 _10339_ (.A(_03420_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand2_1 _10340_ (.A(_03411_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__xnor2_1 _10341_ (.A(_03411_),
    .B(_03422_),
    .Y(_03424_));
 sky130_fd_sc_hd__xor2_1 _10342_ (.A(_03398_),
    .B(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__and2_1 _10343_ (.A(_03388_),
    .B(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__nor2_1 _10344_ (.A(_03388_),
    .B(_03425_),
    .Y(_03427_));
 sky130_fd_sc_hd__nor2_2 _10345_ (.A(_03426_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__xor2_4 _10346_ (.A(_03376_),
    .B(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__o21ba_1 _10347_ (.A1(_03280_),
    .A2(_03297_),
    .B1_N(_03279_),
    .X(_03430_));
 sky130_fd_sc_hd__a21o_1 _10348_ (.A1(_03282_),
    .A2(_03295_),
    .B1(_03294_),
    .X(_03431_));
 sky130_fd_sc_hd__o21ba_1 _10349_ (.A1(_03233_),
    .A2(_03261_),
    .B1_N(_03260_),
    .X(_03432_));
 sky130_fd_sc_hd__o21ba_1 _10350_ (.A1(_03264_),
    .A2(_03276_),
    .B1_N(_03275_),
    .X(_03433_));
 sky130_fd_sc_hd__nor2_1 _10351_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__xor2_2 _10352_ (.A(_03432_),
    .B(_03433_),
    .X(_03435_));
 sky130_fd_sc_hd__xnor2_2 _10353_ (.A(_03431_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21bo_1 _10354_ (.A1(_03300_),
    .A2(_03304_),
    .B1_N(_03303_),
    .X(_03437_));
 sky130_fd_sc_hd__nand2b_1 _10355_ (.A_N(_03436_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_2 _10356_ (.A(_03436_),
    .B(_03437_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2b_1 _10357_ (.A_N(_03430_),
    .B(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__xnor2_2 _10358_ (.A(_03430_),
    .B(_03439_),
    .Y(_03441_));
 sky130_fd_sc_hd__and2_1 _10359_ (.A(_03429_),
    .B(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__xor2_4 _10360_ (.A(_03429_),
    .B(_03441_),
    .X(_03443_));
 sky130_fd_sc_hd__xor2_4 _10361_ (.A(_03361_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(_03360_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__or2_1 _10363_ (.A(_03360_),
    .B(_03444_),
    .X(_03446_));
 sky130_fd_sc_hd__xnor2_4 _10364_ (.A(_03360_),
    .B(_03444_),
    .Y(_03447_));
 sky130_fd_sc_hd__a21oi_1 _10365_ (.A1(_03179_),
    .A2(_03313_),
    .B1(_03314_),
    .Y(_03448_));
 sky130_fd_sc_hd__nor2_1 _10366_ (.A(_03181_),
    .B(_03315_),
    .Y(_03449_));
 sky130_fd_sc_hd__a21oi_2 _10367_ (.A1(_03183_),
    .A2(_03449_),
    .B1(_03448_),
    .Y(_03450_));
 sky130_fd_sc_hd__or4_2 _10368_ (.A(_02895_),
    .B(_03035_),
    .C(_03181_),
    .D(_03315_),
    .X(_03451_));
 sky130_fd_sc_hd__a211o_1 _10369_ (.A1(_02063_),
    .A2(_02067_),
    .B1(_02793_),
    .C1(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__o211ai_4 _10370_ (.A1(_02796_),
    .A2(_03451_),
    .B1(_03452_),
    .C1(_03450_),
    .Y(_03453_));
 sky130_fd_sc_hd__xnor2_2 _10371_ (.A(_03447_),
    .B(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21oi_1 _10372_ (.A1(net159),
    .A2(_03359_),
    .B1(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__and3_1 _10373_ (.A(net159),
    .B(_03359_),
    .C(_03454_),
    .X(_03456_));
 sky130_fd_sc_hd__a21oi_1 _10374_ (.A1(net161),
    .A2(_02085_),
    .B1(_02086_),
    .Y(_03457_));
 sky130_fd_sc_hd__a31o_1 _10375_ (.A1(net161),
    .A2(_02085_),
    .A3(_02086_),
    .B1(_02254_),
    .X(_03458_));
 sky130_fd_sc_hd__o21a_1 _10376_ (.A1(_06274_),
    .A2(_03325_),
    .B1(_06282_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _10377_ (.A0(_06359_),
    .A1(_03459_),
    .S(net304),
    .X(_03460_));
 sky130_fd_sc_hd__nor2_1 _10378_ (.A(_06238_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a211o_1 _10379_ (.A1(_06238_),
    .A2(_03460_),
    .B1(_03461_),
    .C1(net255),
    .X(_03462_));
 sky130_fd_sc_hd__o21a_1 _10380_ (.A1(_03347_),
    .A2(_03348_),
    .B1(_03349_),
    .X(_03463_));
 sky130_fd_sc_hd__nor2_1 _10381_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03465_));
 sky130_fd_sc_hd__nand2b_1 _10383_ (.A_N(_03464_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__xnor2_1 _10384_ (.A(_03463_),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__or2_1 _10385_ (.A(net238),
    .B(_02221_),
    .X(_03468_));
 sky130_fd_sc_hd__o211a_1 _10386_ (.A1(net237),
    .A2(_02205_),
    .B1(_03468_),
    .C1(net239),
    .X(_03469_));
 sky130_fd_sc_hd__a21oi_2 _10387_ (.A1(net241),
    .A2(_03329_),
    .B1(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(_03467_),
    .A1(_03470_),
    .S(net243),
    .X(_03471_));
 sky130_fd_sc_hd__or2_1 _10389_ (.A(\div_res[7] ),
    .B(_03337_),
    .X(_03472_));
 sky130_fd_sc_hd__a21oi_1 _10390_ (.A1(net165),
    .A2(_03472_),
    .B1(\div_res[8] ),
    .Y(_03473_));
 sky130_fd_sc_hd__a31o_1 _10391_ (.A1(\div_res[8] ),
    .A2(net165),
    .A3(_03472_),
    .B1(net204),
    .X(_03474_));
 sky130_fd_sc_hd__a21oi_1 _10392_ (.A1(_06229_),
    .A2(_02249_),
    .B1(_02245_),
    .Y(_03475_));
 sky130_fd_sc_hd__or2_1 _10393_ (.A(\div_shifter[39] ),
    .B(_03340_),
    .X(_03476_));
 sky130_fd_sc_hd__a21oi_1 _10394_ (.A1(net247),
    .A2(_03476_),
    .B1(\div_shifter[40] ),
    .Y(_03477_));
 sky130_fd_sc_hd__a31o_1 _10395_ (.A1(\div_shifter[40] ),
    .A2(net247),
    .A3(_03476_),
    .B1(net250),
    .X(_03478_));
 sky130_fd_sc_hd__o2bb2a_1 _10396_ (.A1_N(_06202_),
    .A2_N(_06459_),
    .B1(_03477_),
    .B2(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__o221a_1 _10397_ (.A1(_06229_),
    .A2(net206),
    .B1(_03475_),
    .B2(_06220_),
    .C1(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__o21ai_2 _10398_ (.A1(net241),
    .A2(_03335_),
    .B1(_02272_),
    .Y(_03481_));
 sky130_fd_sc_hd__o221a_1 _10399_ (.A1(_03473_),
    .A2(_03474_),
    .B1(_03481_),
    .B2(net190),
    .C1(_03480_),
    .X(_03482_));
 sky130_fd_sc_hd__o221a_1 _10400_ (.A1(net188),
    .A2(_03470_),
    .B1(_03471_),
    .B2(_06447_),
    .C1(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__o211a_1 _10401_ (.A1(_03457_),
    .A2(_03458_),
    .B1(_03462_),
    .C1(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__o31a_1 _10402_ (.A1(net209),
    .A2(_03455_),
    .A3(_03456_),
    .B1(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__and3_1 _10403_ (.A(curr_PC[7]),
    .B(curr_PC[8]),
    .C(_03223_),
    .X(_03486_));
 sky130_fd_sc_hd__a21oi_1 _10404_ (.A1(curr_PC[7]),
    .A2(_03223_),
    .B1(curr_PC[8]),
    .Y(_03487_));
 sky130_fd_sc_hd__or3_1 _10405_ (.A(net262),
    .B(_03486_),
    .C(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__o21ai_4 _10406_ (.A1(net267),
    .A2(_03485_),
    .B1(_03488_),
    .Y(dest_val[8]));
 sky130_fd_sc_hd__nand2_1 _10407_ (.A(curr_PC[9]),
    .B(_03486_),
    .Y(_03489_));
 sky130_fd_sc_hd__or2_1 _10408_ (.A(curr_PC[9]),
    .B(_03486_),
    .X(_03490_));
 sky130_fd_sc_hd__and2_1 _10409_ (.A(_03489_),
    .B(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__nor2_1 _10410_ (.A(_03359_),
    .B(_03454_),
    .Y(_03492_));
 sky130_fd_sc_hd__a21o_2 _10411_ (.A1(_03361_),
    .A2(_03443_),
    .B1(_03442_),
    .X(_03493_));
 sky130_fd_sc_hd__and2_2 _10412_ (.A(_03438_),
    .B(_03440_),
    .X(_03494_));
 sky130_fd_sc_hd__or4_1 _10413_ (.A(net137),
    .B(net32),
    .C(_03379_),
    .D(_03381_),
    .X(_03495_));
 sky130_fd_sc_hd__o22ai_1 _10414_ (.A1(net137),
    .A2(net32),
    .B1(_03379_),
    .B2(_03381_),
    .Y(_03496_));
 sky130_fd_sc_hd__and2_1 _10415_ (.A(_03495_),
    .B(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__xor2_1 _10416_ (.A(_03406_),
    .B(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_1 _10417_ (.A1(_00137_),
    .A2(_00138_),
    .B1(net123),
    .X(_03499_));
 sky130_fd_sc_hd__or2_1 _10418_ (.A(net119),
    .B(net70),
    .X(_03500_));
 sky130_fd_sc_hd__nand3_1 _10419_ (.A(net108),
    .B(_03499_),
    .C(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__a21o_1 _10420_ (.A1(_03499_),
    .A2(_03500_),
    .B1(net108),
    .X(_03502_));
 sky130_fd_sc_hd__o32a_1 _10421_ (.A1(_00176_),
    .A2(_00177_),
    .A3(net42),
    .B1(net39),
    .B2(net66),
    .X(_03503_));
 sky130_fd_sc_hd__xor2_1 _10422_ (.A(net103),
    .B(_03503_),
    .X(_03504_));
 sky130_fd_sc_hd__a21oi_1 _10423_ (.A1(_03501_),
    .A2(_03502_),
    .B1(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand3_1 _10424_ (.A(_03501_),
    .B(_03502_),
    .C(_03504_),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2b_1 _10425_ (.A_N(_03505_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__o22a_1 _10426_ (.A1(net25),
    .A2(net84),
    .B1(net80),
    .B2(net72),
    .X(_03508_));
 sky130_fd_sc_hd__xnor2_1 _10427_ (.A(net105),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__xnor2_1 _10428_ (.A(_03507_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__and2_1 _10429_ (.A(_03498_),
    .B(_03510_),
    .X(_03511_));
 sky130_fd_sc_hd__xor2_1 _10430_ (.A(_03498_),
    .B(_03510_),
    .X(_03512_));
 sky130_fd_sc_hd__o22a_1 _10431_ (.A1(net96),
    .A2(net16),
    .B1(net37),
    .B2(net89),
    .X(_03513_));
 sky130_fd_sc_hd__xnor2_1 _10432_ (.A(net77),
    .B(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__inv_2 _10433_ (.A(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__o22a_1 _10434_ (.A1(net98),
    .A2(net10),
    .B1(net5),
    .B2(net135),
    .X(_03516_));
 sky130_fd_sc_hd__xnor2_1 _10435_ (.A(net33),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__o22a_1 _10436_ (.A1(net117),
    .A2(net30),
    .B1(net28),
    .B2(net113),
    .X(_03518_));
 sky130_fd_sc_hd__xnor2_1 _10437_ (.A(net112),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__nand2_1 _10438_ (.A(_03517_),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__xor2_1 _10439_ (.A(_03517_),
    .B(_03519_),
    .X(_03521_));
 sky130_fd_sc_hd__xnor2_1 _10440_ (.A(_03514_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__xnor2_1 _10441_ (.A(_03512_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__a21o_1 _10442_ (.A1(_03368_),
    .A2(_03370_),
    .B1(_03366_),
    .X(_03524_));
 sky130_fd_sc_hd__o22a_1 _10443_ (.A1(net88),
    .A2(net13),
    .B1(net6),
    .B2(_00299_),
    .X(_03525_));
 sky130_fd_sc_hd__xnor2_1 _10444_ (.A(_06470_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__or2_1 _10445_ (.A(net125),
    .B(net57),
    .X(_03527_));
 sky130_fd_sc_hd__a21o_1 _10446_ (.A1(_00243_),
    .A2(_00244_),
    .B1(net121),
    .X(_03528_));
 sky130_fd_sc_hd__a21o_1 _10447_ (.A1(_03527_),
    .A2(_03528_),
    .B1(net152),
    .X(_03529_));
 sky130_fd_sc_hd__nand3_1 _10448_ (.A(net152),
    .B(_03527_),
    .C(_03528_),
    .Y(_03530_));
 sky130_fd_sc_hd__and3_1 _10449_ (.A(net167),
    .B(_03529_),
    .C(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__a21o_1 _10450_ (.A1(_03529_),
    .A2(_03530_),
    .B1(net167),
    .X(_03532_));
 sky130_fd_sc_hd__nand2b_1 _10451_ (.A_N(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__xnor2_1 _10452_ (.A(_03526_),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__o21ai_1 _10453_ (.A1(_03416_),
    .A2(_03420_),
    .B1(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__or3_1 _10454_ (.A(_03416_),
    .B(_03420_),
    .C(_03534_),
    .X(_03536_));
 sky130_fd_sc_hd__and3_1 _10455_ (.A(_03524_),
    .B(_03535_),
    .C(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__a21oi_1 _10456_ (.A1(_03535_),
    .A2(_03536_),
    .B1(_03524_),
    .Y(_03538_));
 sky130_fd_sc_hd__or2_1 _10457_ (.A(_03537_),
    .B(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__nor2_1 _10458_ (.A(_03523_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__nand2_1 _10459_ (.A(_03523_),
    .B(_03539_),
    .Y(_03541_));
 sky130_fd_sc_hd__nand2b_2 _10460_ (.A_N(_03540_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__o22a_1 _10461_ (.A1(net74),
    .A2(net62),
    .B1(net59),
    .B2(net115),
    .X(_03543_));
 sky130_fd_sc_hd__xnor2_1 _10462_ (.A(net149),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__o22a_1 _10463_ (.A1(net20),
    .A2(net48),
    .B1(net45),
    .B2(net64),
    .X(_03545_));
 sky130_fd_sc_hd__xor2_1 _10464_ (.A(net91),
    .B(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__xnor2_1 _10465_ (.A(_03544_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__o22a_1 _10466_ (.A1(net68),
    .A2(net54),
    .B1(net51),
    .B2(net94),
    .X(_03548_));
 sky130_fd_sc_hd__xnor2_1 _10467_ (.A(net100),
    .B(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__and2b_1 _10468_ (.A_N(_03547_),
    .B(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__xnor2_1 _10469_ (.A(_03547_),
    .B(_03549_),
    .Y(_03551_));
 sky130_fd_sc_hd__o21a_1 _10470_ (.A1(_03394_),
    .A2(_03396_),
    .B1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__nor3_1 _10471_ (.A(_03394_),
    .B(_03396_),
    .C(_03551_),
    .Y(_03553_));
 sky130_fd_sc_hd__or2_1 _10472_ (.A(_03552_),
    .B(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__a21oi_2 _10473_ (.A1(_03408_),
    .A2(_03410_),
    .B1(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__and3_1 _10474_ (.A(_03408_),
    .B(_03410_),
    .C(_03554_),
    .X(_03556_));
 sky130_fd_sc_hd__nor2_2 _10475_ (.A(_03555_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__xnor2_4 _10476_ (.A(_03542_),
    .B(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__a21o_1 _10477_ (.A1(_03376_),
    .A2(_03428_),
    .B1(_03426_),
    .X(_03559_));
 sky130_fd_sc_hd__a21o_1 _10478_ (.A1(_03431_),
    .A2(_03435_),
    .B1(_03434_),
    .X(_03560_));
 sky130_fd_sc_hd__o21ai_2 _10479_ (.A1(_03371_),
    .A2(_03372_),
    .B1(_03374_),
    .Y(_03561_));
 sky130_fd_sc_hd__or2_1 _10480_ (.A(_03384_),
    .B(_03386_),
    .X(_03562_));
 sky130_fd_sc_hd__o21a_1 _10481_ (.A1(_03398_),
    .A2(_03424_),
    .B1(_03423_),
    .X(_03563_));
 sky130_fd_sc_hd__o21ba_1 _10482_ (.A1(_03384_),
    .A2(_03386_),
    .B1_N(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__xnor2_2 _10483_ (.A(_03562_),
    .B(_03563_),
    .Y(_03565_));
 sky130_fd_sc_hd__xor2_2 _10484_ (.A(_03561_),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__xnor2_2 _10485_ (.A(_03560_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__and2b_1 _10486_ (.A_N(_03567_),
    .B(_03559_),
    .X(_03568_));
 sky130_fd_sc_hd__xnor2_4 _10487_ (.A(_03559_),
    .B(_03567_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _10488_ (.A(_03558_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__xnor2_4 _10489_ (.A(_03558_),
    .B(_03569_),
    .Y(_03571_));
 sky130_fd_sc_hd__xnor2_4 _10490_ (.A(_03494_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2b_1 _10491_ (.A_N(_03572_),
    .B(_03493_),
    .Y(_03573_));
 sky130_fd_sc_hd__and2b_1 _10492_ (.A_N(_03493_),
    .B(_03572_),
    .X(_03574_));
 sky130_fd_sc_hd__xor2_4 _10493_ (.A(_03493_),
    .B(_03572_),
    .X(_03575_));
 sky130_fd_sc_hd__a21bo_1 _10494_ (.A1(_03313_),
    .A2(_03445_),
    .B1_N(_03446_),
    .X(_03576_));
 sky130_fd_sc_hd__o31a_1 _10495_ (.A1(_03315_),
    .A2(_03317_),
    .A3(_03447_),
    .B1(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__or4_1 _10496_ (.A(_03035_),
    .B(_03181_),
    .C(_03315_),
    .D(_03447_),
    .X(_03578_));
 sky130_fd_sc_hd__o21bai_2 _10497_ (.A1(_03036_),
    .A2(_03037_),
    .B1_N(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__a211o_1 _10498_ (.A1(_02395_),
    .A2(_02396_),
    .B1(_03039_),
    .C1(_03578_),
    .X(_03580_));
 sky130_fd_sc_hd__and3_1 _10499_ (.A(_03577_),
    .B(_03579_),
    .C(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__xnor2_2 _10500_ (.A(_03575_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__o21ai_1 _10501_ (.A1(net155),
    .A2(_03492_),
    .B1(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__o311a_1 _10502_ (.A1(net155),
    .A2(_03492_),
    .A3(_03582_),
    .B1(_03583_),
    .C1(_02171_),
    .X(_03584_));
 sky130_fd_sc_hd__or3_1 _10503_ (.A(net157),
    .B(_02087_),
    .C(_02091_),
    .X(_03585_));
 sky130_fd_sc_hd__o21ai_1 _10504_ (.A1(net157),
    .A2(_02087_),
    .B1(_02091_),
    .Y(_03586_));
 sky130_fd_sc_hd__o21a_1 _10505_ (.A1(_06220_),
    .A2(_03459_),
    .B1(_06229_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(_06360_),
    .A1(_03587_),
    .S(net304),
    .X(_03588_));
 sky130_fd_sc_hd__nor2_1 _10507_ (.A(_06185_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__a211o_1 _10508_ (.A1(_06185_),
    .A2(_03588_),
    .B1(_03589_),
    .C1(net255),
    .X(_03590_));
 sky130_fd_sc_hd__o21a_1 _10509_ (.A1(_03463_),
    .A2(_03464_),
    .B1(_03465_),
    .X(_03591_));
 sky130_fd_sc_hd__nor2_1 _10510_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_1 _10511_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2b_1 _10512_ (.A_N(_03592_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__xnor2_1 _10513_ (.A(_03591_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(_02414_),
    .A1(_02422_),
    .S(net236),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(_03196_),
    .A1(_03596_),
    .S(net239),
    .X(_03597_));
 sky130_fd_sc_hd__inv_2 _10516_ (.A(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(_03595_),
    .A1(_03598_),
    .S(net243),
    .X(_03599_));
 sky130_fd_sc_hd__or2_1 _10518_ (.A(\div_res[8] ),
    .B(_03472_),
    .X(_03600_));
 sky130_fd_sc_hd__a21oi_1 _10519_ (.A1(net163),
    .A2(_03600_),
    .B1(\div_res[9] ),
    .Y(_03601_));
 sky130_fd_sc_hd__a31o_1 _10520_ (.A1(\div_res[9] ),
    .A2(net163),
    .A3(_03600_),
    .B1(net204),
    .X(_03602_));
 sky130_fd_sc_hd__a21oi_1 _10521_ (.A1(_06176_),
    .A2(_02249_),
    .B1(_02245_),
    .Y(_03603_));
 sky130_fd_sc_hd__or3_2 _10522_ (.A(\div_shifter[40] ),
    .B(\div_shifter[39] ),
    .C(_03340_),
    .X(_03604_));
 sky130_fd_sc_hd__a21oi_2 _10523_ (.A1(net247),
    .A2(_03604_),
    .B1(\div_shifter[41] ),
    .Y(_03605_));
 sky130_fd_sc_hd__a31o_1 _10524_ (.A1(\div_shifter[41] ),
    .A2(net249),
    .A3(_03604_),
    .B1(net250),
    .X(_03606_));
 sky130_fd_sc_hd__a221oi_1 _10525_ (.A1(_06150_),
    .A2(_06459_),
    .B1(_02255_),
    .B2(_06168_),
    .C1(_06424_),
    .Y(_03607_));
 sky130_fd_sc_hd__o221a_1 _10526_ (.A1(_06162_),
    .A2(_03603_),
    .B1(_03605_),
    .B2(_03606_),
    .C1(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__o21a_1 _10527_ (.A1(_03601_),
    .A2(_03602_),
    .B1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__o21ai_2 _10528_ (.A1(net240),
    .A2(_03203_),
    .B1(_02272_),
    .Y(_03610_));
 sky130_fd_sc_hd__o221a_1 _10529_ (.A1(net188),
    .A2(_03598_),
    .B1(_03610_),
    .B2(net190),
    .C1(_03609_),
    .X(_03611_));
 sky130_fd_sc_hd__o211ai_2 _10530_ (.A1(_06447_),
    .A2(_03599_),
    .B1(_03611_),
    .C1(_03590_),
    .Y(_03612_));
 sky130_fd_sc_hd__a31o_1 _10531_ (.A1(net252),
    .A2(_03585_),
    .A3(_03586_),
    .B1(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__o22a_4 _10532_ (.A1(net262),
    .A2(_03491_),
    .B1(_03584_),
    .B2(_03613_),
    .X(dest_val[9]));
 sky130_fd_sc_hd__a21o_1 _10533_ (.A1(_03492_),
    .A2(_03582_),
    .B1(net155),
    .X(_03614_));
 sky130_fd_sc_hd__o21a_2 _10534_ (.A1(_03494_),
    .A2(_03571_),
    .B1(_03570_),
    .X(_03615_));
 sky130_fd_sc_hd__a21o_2 _10535_ (.A1(_03560_),
    .A2(_03566_),
    .B1(_03568_),
    .X(_03616_));
 sky130_fd_sc_hd__a21bo_1 _10536_ (.A1(_03406_),
    .A2(_03496_),
    .B1_N(_03495_),
    .X(_03617_));
 sky130_fd_sc_hd__o22a_1 _10537_ (.A1(net126),
    .A2(net18),
    .B1(net13),
    .B2(net121),
    .X(_03618_));
 sky130_fd_sc_hd__xnor2_1 _10538_ (.A(net153),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__o22a_1 _10539_ (.A1(net94),
    .A2(net62),
    .B1(net51),
    .B2(net68),
    .X(_03620_));
 sky130_fd_sc_hd__xnor2_1 _10540_ (.A(_00153_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__nor2_1 _10541_ (.A(_03619_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__and2_1 _10542_ (.A(_03619_),
    .B(_03621_),
    .X(_03623_));
 sky130_fd_sc_hd__or2_2 _10543_ (.A(_03622_),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__o22a_1 _10544_ (.A1(net74),
    .A2(net59),
    .B1(net56),
    .B2(net115),
    .X(_03625_));
 sky130_fd_sc_hd__xnor2_2 _10545_ (.A(net149),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__xnor2_2 _10546_ (.A(_03624_),
    .B(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__a21bo_1 _10547_ (.A1(_03515_),
    .A2(_03521_),
    .B1_N(_03520_),
    .X(_03628_));
 sky130_fd_sc_hd__nand2b_1 _10548_ (.A_N(_03627_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__xor2_2 _10549_ (.A(_03627_),
    .B(_03628_),
    .X(_03630_));
 sky130_fd_sc_hd__nand2b_1 _10550_ (.A_N(_03630_),
    .B(_03617_),
    .Y(_03631_));
 sky130_fd_sc_hd__xor2_2 _10551_ (.A(_03617_),
    .B(_03630_),
    .X(_03632_));
 sky130_fd_sc_hd__o22a_1 _10552_ (.A1(net89),
    .A2(net16),
    .B1(net37),
    .B2(net117),
    .X(_03633_));
 sky130_fd_sc_hd__xnor2_1 _10553_ (.A(net77),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__inv_2 _10554_ (.A(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__o22a_1 _10555_ (.A1(net119),
    .A2(net23),
    .B1(net70),
    .B2(net85),
    .X(_03636_));
 sky130_fd_sc_hd__xnor2_1 _10556_ (.A(net108),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__xor2_1 _10557_ (.A(_03634_),
    .B(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__o22a_1 _10558_ (.A1(net113),
    .A2(net30),
    .B1(net28),
    .B2(net123),
    .X(_03639_));
 sky130_fd_sc_hd__xnor2_1 _10559_ (.A(net112),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__and2b_1 _10560_ (.A_N(_03638_),
    .B(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__and2b_1 _10561_ (.A_N(_03640_),
    .B(_03638_),
    .X(_03642_));
 sky130_fd_sc_hd__or2_2 _10562_ (.A(_03641_),
    .B(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__a21o_1 _10563_ (.A1(_03526_),
    .A2(_03532_),
    .B1(_03531_),
    .X(_03644_));
 sky130_fd_sc_hd__o22a_1 _10564_ (.A1(net96),
    .A2(net10),
    .B1(net5),
    .B2(net98),
    .X(_03645_));
 sky130_fd_sc_hd__xnor2_2 _10565_ (.A(net33),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__xor2_2 _10566_ (.A(_03644_),
    .B(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__or2_1 _10567_ (.A(net135),
    .B(net32),
    .X(_03648_));
 sky130_fd_sc_hd__and3b_1 _10568_ (.A_N(net135),
    .B(net33),
    .C(_03647_),
    .X(_03649_));
 sky130_fd_sc_hd__xnor2_2 _10569_ (.A(_03647_),
    .B(_03648_),
    .Y(_03650_));
 sky130_fd_sc_hd__or2_1 _10570_ (.A(net20),
    .B(net45),
    .X(_03651_));
 sky130_fd_sc_hd__or2_1 _10571_ (.A(net64),
    .B(net54),
    .X(_03652_));
 sky130_fd_sc_hd__and3_1 _10572_ (.A(net91),
    .B(_03651_),
    .C(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__a21oi_1 _10573_ (.A1(_03651_),
    .A2(_03652_),
    .B1(net91),
    .Y(_03654_));
 sky130_fd_sc_hd__or2_1 _10574_ (.A(net25),
    .B(net80),
    .X(_03655_));
 sky130_fd_sc_hd__or2_1 _10575_ (.A(net72),
    .B(net42),
    .X(_03656_));
 sky130_fd_sc_hd__and3_1 _10576_ (.A(net105),
    .B(_03655_),
    .C(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__a21oi_1 _10577_ (.A1(_03655_),
    .A2(_03656_),
    .B1(net105),
    .Y(_03658_));
 sky130_fd_sc_hd__o22a_1 _10578_ (.A1(_03653_),
    .A2(_03654_),
    .B1(_03657_),
    .B2(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__or4_1 _10579_ (.A(_03653_),
    .B(_03654_),
    .C(_03657_),
    .D(_03658_),
    .X(_03660_));
 sky130_fd_sc_hd__and2b_1 _10580_ (.A_N(_03659_),
    .B(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__o22a_1 _10581_ (.A1(net66),
    .A2(net48),
    .B1(net39),
    .B2(_00178_),
    .X(_03662_));
 sky130_fd_sc_hd__xnor2_2 _10582_ (.A(net102),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__xor2_2 _10583_ (.A(_03661_),
    .B(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__nand2_1 _10584_ (.A(_03650_),
    .B(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__xnor2_2 _10585_ (.A(_03650_),
    .B(_03664_),
    .Y(_03666_));
 sky130_fd_sc_hd__xor2_2 _10586_ (.A(_03643_),
    .B(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__o21ba_1 _10587_ (.A1(_03544_),
    .A2(_03546_),
    .B1_N(_03550_),
    .X(_03668_));
 sky130_fd_sc_hd__a21o_1 _10588_ (.A1(_03506_),
    .A2(_03509_),
    .B1(_03505_),
    .X(_03669_));
 sky130_fd_sc_hd__nor2_1 _10589_ (.A(net88),
    .B(net6),
    .Y(_03670_));
 sky130_fd_sc_hd__xnor2_2 _10590_ (.A(net186),
    .B(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__and2b_1 _10591_ (.A_N(_03671_),
    .B(_03669_),
    .X(_03672_));
 sky130_fd_sc_hd__xnor2_2 _10592_ (.A(_03669_),
    .B(_03671_),
    .Y(_03673_));
 sky130_fd_sc_hd__and2b_1 _10593_ (.A_N(_03668_),
    .B(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__xnor2_2 _10594_ (.A(_03668_),
    .B(_03673_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _10595_ (.A(_03667_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__xnor2_2 _10596_ (.A(_03667_),
    .B(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__xor2_2 _10597_ (.A(_03632_),
    .B(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__a21oi_2 _10598_ (.A1(_03541_),
    .A2(_03557_),
    .B1(_03540_),
    .Y(_03679_));
 sky130_fd_sc_hd__a21o_1 _10599_ (.A1(_03512_),
    .A2(_03522_),
    .B1(_03511_),
    .X(_03680_));
 sky130_fd_sc_hd__a21bo_1 _10600_ (.A1(_03524_),
    .A2(_03536_),
    .B1_N(_03535_),
    .X(_03681_));
 sky130_fd_sc_hd__xor2_1 _10601_ (.A(_03680_),
    .B(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__o21a_1 _10602_ (.A1(_03552_),
    .A2(_03555_),
    .B1(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__nor3_1 _10603_ (.A(_03552_),
    .B(_03555_),
    .C(_03682_),
    .Y(_03684_));
 sky130_fd_sc_hd__or2_2 _10604_ (.A(_03683_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__a21oi_2 _10605_ (.A1(_03561_),
    .A2(_03565_),
    .B1(_03564_),
    .Y(_03686_));
 sky130_fd_sc_hd__xor2_2 _10606_ (.A(_03685_),
    .B(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__nand2b_1 _10607_ (.A_N(_03679_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__xnor2_2 _10608_ (.A(_03679_),
    .B(_03687_),
    .Y(_03689_));
 sky130_fd_sc_hd__and2_1 _10609_ (.A(_03678_),
    .B(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__or2_1 _10610_ (.A(_03678_),
    .B(_03689_),
    .X(_03691_));
 sky130_fd_sc_hd__xor2_2 _10611_ (.A(_03678_),
    .B(_03689_),
    .X(_03692_));
 sky130_fd_sc_hd__xnor2_4 _10612_ (.A(_03616_),
    .B(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__or2_1 _10613_ (.A(_03615_),
    .B(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__and2_1 _10614_ (.A(_03615_),
    .B(_03693_),
    .X(_03695_));
 sky130_fd_sc_hd__xnor2_4 _10615_ (.A(_03615_),
    .B(_03693_),
    .Y(_03696_));
 sky130_fd_sc_hd__nor2_1 _10616_ (.A(_03447_),
    .B(_03575_),
    .Y(_03697_));
 sky130_fd_sc_hd__or4_2 _10617_ (.A(_03181_),
    .B(_03315_),
    .C(_03447_),
    .D(_03575_),
    .X(_03698_));
 sky130_fd_sc_hd__o21bai_2 _10618_ (.A1(_03183_),
    .A2(_03184_),
    .B1_N(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21oi_1 _10619_ (.A1(_03445_),
    .A2(_03573_),
    .B1(_03574_),
    .Y(_03700_));
 sky130_fd_sc_hd__a21oi_1 _10620_ (.A1(_03448_),
    .A2(_03697_),
    .B1(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__o311ai_4 _10621_ (.A1(_02577_),
    .A2(_03182_),
    .A3(_03698_),
    .B1(_03699_),
    .C1(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__xor2_2 _10622_ (.A(_03696_),
    .B(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__nand2_1 _10623_ (.A(_03614_),
    .B(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__or2_1 _10624_ (.A(_03614_),
    .B(_03703_),
    .X(_03705_));
 sky130_fd_sc_hd__or3_1 _10625_ (.A(net157),
    .B(_02092_),
    .C(_02093_),
    .X(_03706_));
 sky130_fd_sc_hd__o21ai_1 _10626_ (.A1(net157),
    .A2(_02092_),
    .B1(_02093_),
    .Y(_03707_));
 sky130_fd_sc_hd__o21ai_1 _10627_ (.A1(_06162_),
    .A2(_03587_),
    .B1(_06176_),
    .Y(_03708_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(_06361_),
    .A1(_03708_),
    .S(net303),
    .X(_03709_));
 sky130_fd_sc_hd__nand2_1 _10629_ (.A(_06138_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__o211a_1 _10630_ (.A1(_06138_),
    .A2(_03709_),
    .B1(_03710_),
    .C1(_02247_),
    .X(_03711_));
 sky130_fd_sc_hd__or2_1 _10631_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03712_));
 sky130_fd_sc_hd__and2_1 _10632_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03713_));
 sky130_fd_sc_hd__nand2_1 _10633_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03714_));
 sky130_fd_sc_hd__o21ai_1 _10634_ (.A1(_03591_),
    .A2(_03592_),
    .B1(_03593_),
    .Y(_03715_));
 sky130_fd_sc_hd__a21oi_1 _10635_ (.A1(_03712_),
    .A2(_03714_),
    .B1(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__and3_1 _10636_ (.A(_03712_),
    .B(_03714_),
    .C(_03715_),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(_02592_),
    .A1(_02596_),
    .S(net236),
    .X(_03718_));
 sky130_fd_sc_hd__mux2_2 _10638_ (.A0(_03052_),
    .A1(_03718_),
    .S(net239),
    .X(_03719_));
 sky130_fd_sc_hd__o21ai_1 _10639_ (.A1(_03716_),
    .A2(_03717_),
    .B1(net268),
    .Y(_03720_));
 sky130_fd_sc_hd__o211a_1 _10640_ (.A1(net268),
    .A2(_03719_),
    .B1(_03720_),
    .C1(net216),
    .X(_03721_));
 sky130_fd_sc_hd__or2_1 _10641_ (.A(\div_res[9] ),
    .B(_03600_),
    .X(_03722_));
 sky130_fd_sc_hd__a21oi_1 _10642_ (.A1(net163),
    .A2(_03722_),
    .B1(\div_res[10] ),
    .Y(_03723_));
 sky130_fd_sc_hd__a31o_1 _10643_ (.A1(\div_res[10] ),
    .A2(net163),
    .A3(_03722_),
    .B1(net204),
    .X(_03724_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(net253),
    .A1(net206),
    .S(_06126_),
    .X(_03725_));
 sky130_fd_sc_hd__a21oi_1 _10645_ (.A1(net207),
    .A2(_03725_),
    .B1(_06132_),
    .Y(_03726_));
 sky130_fd_sc_hd__or2_1 _10646_ (.A(\div_shifter[41] ),
    .B(_03604_),
    .X(_03727_));
 sky130_fd_sc_hd__a21oi_1 _10647_ (.A1(net247),
    .A2(_03727_),
    .B1(\div_shifter[42] ),
    .Y(_03728_));
 sky130_fd_sc_hd__a311o_2 _10648_ (.A1(\div_shifter[42] ),
    .A2(net247),
    .A3(_03727_),
    .B1(_03728_),
    .C1(net250),
    .X(_03729_));
 sky130_fd_sc_hd__a21oi_1 _10649_ (.A1(_06114_),
    .A2(_06459_),
    .B1(_03726_),
    .Y(_03730_));
 sky130_fd_sc_hd__o211a_1 _10650_ (.A1(_03723_),
    .A2(_03724_),
    .B1(_03729_),
    .C1(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__o21ai_2 _10651_ (.A1(net240),
    .A2(_03063_),
    .B1(_02272_),
    .Y(_03732_));
 sky130_fd_sc_hd__o21ai_1 _10652_ (.A1(net190),
    .A2(_03732_),
    .B1(_03731_),
    .Y(_03733_));
 sky130_fd_sc_hd__a2111o_1 _10653_ (.A1(_02243_),
    .A2(_03719_),
    .B1(_03721_),
    .C1(_03733_),
    .D1(_03711_),
    .X(_03734_));
 sky130_fd_sc_hd__a31o_1 _10654_ (.A1(net252),
    .A2(_03706_),
    .A3(_03707_),
    .B1(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__a31o_1 _10655_ (.A1(_02171_),
    .A2(_03704_),
    .A3(_03705_),
    .B1(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__xnor2_1 _10656_ (.A(curr_PC[10]),
    .B(_03489_),
    .Y(_03737_));
 sky130_fd_sc_hd__mux2_8 _10657_ (.A0(_03736_),
    .A1(_03737_),
    .S(net267),
    .X(dest_val[10]));
 sky130_fd_sc_hd__or4bb_1 _10658_ (.A(_02168_),
    .B(_03454_),
    .C_N(_03582_),
    .D_N(_03703_),
    .X(_03738_));
 sky130_fd_sc_hd__nor2_1 _10659_ (.A(_03358_),
    .B(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__or2_1 _10660_ (.A(net156),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__o21ai_4 _10661_ (.A1(_03685_),
    .A2(_03686_),
    .B1(_03688_),
    .Y(_03741_));
 sky130_fd_sc_hd__o22a_1 _10662_ (.A1(net117),
    .A2(net15),
    .B1(net36),
    .B2(net113),
    .X(_03742_));
 sky130_fd_sc_hd__xnor2_1 _10663_ (.A(net77),
    .B(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__or2_1 _10664_ (.A(net98),
    .B(net32),
    .X(_03744_));
 sky130_fd_sc_hd__xor2_1 _10665_ (.A(_03743_),
    .B(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__o22ai_1 _10666_ (.A1(net89),
    .A2(net10),
    .B1(net4),
    .B2(net96),
    .Y(_03746_));
 sky130_fd_sc_hd__nand2_1 _10667_ (.A(net33),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__or2_1 _10668_ (.A(net33),
    .B(_03746_),
    .X(_03748_));
 sky130_fd_sc_hd__and3_1 _10669_ (.A(_03745_),
    .B(_03747_),
    .C(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__a21oi_1 _10670_ (.A1(_03747_),
    .A2(_03748_),
    .B1(_03745_),
    .Y(_03750_));
 sky130_fd_sc_hd__o22a_1 _10671_ (.A1(net68),
    .A2(net61),
    .B1(net58),
    .B2(net94),
    .X(_03751_));
 sky130_fd_sc_hd__xnor2_1 _10672_ (.A(net100),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__o32a_1 _10673_ (.A1(_00176_),
    .A2(_00177_),
    .A3(net48),
    .B1(net45),
    .B2(net66),
    .X(_03753_));
 sky130_fd_sc_hd__xnor2_1 _10674_ (.A(net102),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__and2_1 _10675_ (.A(_03752_),
    .B(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__nor2_1 _10676_ (.A(_03752_),
    .B(_03754_),
    .Y(_03756_));
 sky130_fd_sc_hd__nor2_1 _10677_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__o22a_1 _10678_ (.A1(net20),
    .A2(net54),
    .B1(net50),
    .B2(net64),
    .X(_03758_));
 sky130_fd_sc_hd__xnor2_1 _10679_ (.A(net91),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__xor2_1 _10680_ (.A(_03757_),
    .B(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__nor3b_1 _10681_ (.A(_03749_),
    .B(_03750_),
    .C_N(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__o21bai_1 _10682_ (.A1(_03749_),
    .A2(_03750_),
    .B1_N(_03760_),
    .Y(_03762_));
 sky130_fd_sc_hd__inv_2 _10683_ (.A(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__o22a_1 _10684_ (.A1(net123),
    .A2(net30),
    .B1(net27),
    .B2(net119),
    .X(_03764_));
 sky130_fd_sc_hd__xnor2_1 _10685_ (.A(net112),
    .B(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__o22a_1 _10686_ (.A1(net25),
    .A2(net42),
    .B1(net39),
    .B2(net72),
    .X(_03766_));
 sky130_fd_sc_hd__xnor2_1 _10687_ (.A(net105),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__and2_1 _10688_ (.A(_03765_),
    .B(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__xor2_1 _10689_ (.A(_03765_),
    .B(_03767_),
    .X(_03769_));
 sky130_fd_sc_hd__o22a_1 _10690_ (.A1(net23),
    .A2(net85),
    .B1(net80),
    .B2(net70),
    .X(_03770_));
 sky130_fd_sc_hd__xnor2_1 _10691_ (.A(net108),
    .B(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__and2_1 _10692_ (.A(_03769_),
    .B(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__nor2_1 _10693_ (.A(_03769_),
    .B(_03771_),
    .Y(_03773_));
 sky130_fd_sc_hd__nor2_1 _10694_ (.A(_03772_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__and3b_1 _10695_ (.A_N(_03761_),
    .B(_03762_),
    .C(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__o21ba_1 _10696_ (.A1(_03761_),
    .A2(_03763_),
    .B1_N(_03774_),
    .X(_03776_));
 sky130_fd_sc_hd__o21bai_2 _10697_ (.A1(_03624_),
    .A2(_03626_),
    .B1_N(_03622_),
    .Y(_03777_));
 sky130_fd_sc_hd__a21o_1 _10698_ (.A1(_03660_),
    .A2(_03663_),
    .B1(_03659_),
    .X(_03778_));
 sky130_fd_sc_hd__and2_1 _10699_ (.A(_03671_),
    .B(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__xor2_1 _10700_ (.A(_03671_),
    .B(_03778_),
    .X(_03780_));
 sky130_fd_sc_hd__xnor2_1 _10701_ (.A(_03777_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__or3_1 _10702_ (.A(_03775_),
    .B(_03776_),
    .C(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__o21ai_1 _10703_ (.A1(_03775_),
    .A2(_03776_),
    .B1(_03781_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _10704_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__a21oi_2 _10705_ (.A1(_03644_),
    .A2(_03646_),
    .B1(_03649_),
    .Y(_03785_));
 sky130_fd_sc_hd__o22a_1 _10706_ (.A1(net125),
    .A2(net13),
    .B1(net6),
    .B2(net121),
    .X(_03786_));
 sky130_fd_sc_hd__xnor2_2 _10707_ (.A(net153),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__o22a_1 _10708_ (.A1(net74),
    .A2(net56),
    .B1(net18),
    .B2(net115),
    .X(_03788_));
 sky130_fd_sc_hd__xnor2_2 _10709_ (.A(net149),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__xnor2_2 _10710_ (.A(net186),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__nand2b_1 _10711_ (.A_N(_03787_),
    .B(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__xnor2_2 _10712_ (.A(_03787_),
    .B(_03790_),
    .Y(_03792_));
 sky130_fd_sc_hd__a21o_1 _10713_ (.A1(_03635_),
    .A2(_03637_),
    .B1(_03641_),
    .X(_03793_));
 sky130_fd_sc_hd__xor2_2 _10714_ (.A(_03792_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__nand2b_1 _10715_ (.A_N(_03785_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__xnor2_2 _10716_ (.A(_03785_),
    .B(_03794_),
    .Y(_03796_));
 sky130_fd_sc_hd__xnor2_2 _10717_ (.A(_03784_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__o21a_1 _10718_ (.A1(_03632_),
    .A2(_03677_),
    .B1(_03676_),
    .X(_03798_));
 sky130_fd_sc_hd__a21o_1 _10719_ (.A1(_03680_),
    .A2(_03681_),
    .B1(_03683_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_03629_),
    .B(_03631_),
    .Y(_03800_));
 sky130_fd_sc_hd__o21ai_2 _10721_ (.A1(_03643_),
    .A2(_03666_),
    .B1(_03665_),
    .Y(_03801_));
 sky130_fd_sc_hd__nor2_1 _10722_ (.A(_03672_),
    .B(_03674_),
    .Y(_03802_));
 sky130_fd_sc_hd__o21a_1 _10723_ (.A1(_03672_),
    .A2(_03674_),
    .B1(_03801_),
    .X(_03803_));
 sky130_fd_sc_hd__xnor2_1 _10724_ (.A(_03801_),
    .B(_03802_),
    .Y(_03804_));
 sky130_fd_sc_hd__xnor2_1 _10725_ (.A(_03800_),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__and2b_1 _10726_ (.A_N(_03805_),
    .B(_03799_),
    .X(_03806_));
 sky130_fd_sc_hd__xnor2_2 _10727_ (.A(_03799_),
    .B(_03805_),
    .Y(_03807_));
 sky130_fd_sc_hd__and2b_1 _10728_ (.A_N(_03798_),
    .B(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__xnor2_2 _10729_ (.A(_03798_),
    .B(_03807_),
    .Y(_03809_));
 sky130_fd_sc_hd__nand2_1 _10730_ (.A(_03797_),
    .B(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__xnor2_2 _10731_ (.A(_03797_),
    .B(_03809_),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2b_1 _10732_ (.A_N(_03811_),
    .B(_03741_),
    .Y(_03812_));
 sky130_fd_sc_hd__xor2_4 _10733_ (.A(_03741_),
    .B(_03811_),
    .X(_03813_));
 sky130_fd_sc_hd__a21oi_4 _10734_ (.A1(_03616_),
    .A2(_03691_),
    .B1(_03690_),
    .Y(_03814_));
 sky130_fd_sc_hd__or2_1 _10735_ (.A(_03813_),
    .B(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _10736_ (.A(_03813_),
    .B(_03814_),
    .X(_03816_));
 sky130_fd_sc_hd__xnor2_4 _10737_ (.A(_03813_),
    .B(_03814_),
    .Y(_03817_));
 sky130_fd_sc_hd__a21o_1 _10738_ (.A1(_03573_),
    .A2(_03694_),
    .B1(_03695_),
    .X(_03818_));
 sky130_fd_sc_hd__or2_1 _10739_ (.A(_03575_),
    .B(_03696_),
    .X(_03819_));
 sky130_fd_sc_hd__o21a_1 _10740_ (.A1(_03576_),
    .A2(_03819_),
    .B1(_03818_),
    .X(_03820_));
 sky130_fd_sc_hd__or3_1 _10741_ (.A(_03315_),
    .B(_03447_),
    .C(_03819_),
    .X(_03821_));
 sky130_fd_sc_hd__a21o_1 _10742_ (.A1(_03317_),
    .A2(_03318_),
    .B1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__o311a_2 _10743_ (.A1(_02739_),
    .A2(_03316_),
    .A3(_03821_),
    .B1(_03822_),
    .C1(_03820_),
    .X(_03823_));
 sky130_fd_sc_hd__xnor2_4 _10744_ (.A(_03817_),
    .B(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__inv_2 _10745_ (.A(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__a21oi_1 _10746_ (.A1(_03740_),
    .A2(_03824_),
    .B1(net209),
    .Y(_03826_));
 sky130_fd_sc_hd__o21a_1 _10747_ (.A1(_03740_),
    .A2(_03824_),
    .B1(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__or3_1 _10748_ (.A(net157),
    .B(_02094_),
    .C(_02097_),
    .X(_03828_));
 sky130_fd_sc_hd__o21ai_1 _10749_ (.A1(net157),
    .A2(_02094_),
    .B1(_02097_),
    .Y(_03829_));
 sky130_fd_sc_hd__a21o_1 _10750_ (.A1(_06138_),
    .A2(_03708_),
    .B1(_06126_),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(_06362_),
    .A1(_03830_),
    .S(net303),
    .X(_03831_));
 sky130_fd_sc_hd__nand2_1 _10752_ (.A(_06102_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__o211a_1 _10753_ (.A1(_06102_),
    .A2(_03831_),
    .B1(_03832_),
    .C1(_02247_),
    .X(_03833_));
 sky130_fd_sc_hd__or2_1 _10754_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03834_));
 sky130_fd_sc_hd__and2_1 _10755_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03835_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .Y(_03836_));
 sky130_fd_sc_hd__a211o_1 _10757_ (.A1(_03834_),
    .A2(_03836_),
    .B1(_03713_),
    .C1(_03717_),
    .X(_03837_));
 sky130_fd_sc_hd__o211a_1 _10758_ (.A1(_03713_),
    .A2(_03717_),
    .B1(_03834_),
    .C1(_03836_),
    .X(_03838_));
 sky130_fd_sc_hd__or3b_1 _10759_ (.A(_03838_),
    .B(net243),
    .C_N(_03837_),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(_02752_),
    .A1(_02756_),
    .S(net237),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _10761_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(_02907_),
    .A1(_03841_),
    .S(net239),
    .X(_03842_));
 sky130_fd_sc_hd__o21ai_1 _10763_ (.A1(net268),
    .A2(_03842_),
    .B1(_03839_),
    .Y(_03843_));
 sky130_fd_sc_hd__or2_1 _10764_ (.A(\div_res[10] ),
    .B(_03722_),
    .X(_03844_));
 sky130_fd_sc_hd__a21oi_1 _10765_ (.A1(net163),
    .A2(_03844_),
    .B1(\div_res[11] ),
    .Y(_03845_));
 sky130_fd_sc_hd__a31o_1 _10766_ (.A1(\div_res[11] ),
    .A2(net162),
    .A3(_03844_),
    .B1(net204),
    .X(_03846_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(net253),
    .A1(net206),
    .S(_06087_),
    .X(_03847_));
 sky130_fd_sc_hd__a21o_1 _10768_ (.A1(net207),
    .A2(_03847_),
    .B1(_06096_),
    .X(_03848_));
 sky130_fd_sc_hd__or2_1 _10769_ (.A(\div_shifter[42] ),
    .B(_03727_),
    .X(_03849_));
 sky130_fd_sc_hd__a21oi_1 _10770_ (.A1(net249),
    .A2(_03849_),
    .B1(\div_shifter[43] ),
    .Y(_03850_));
 sky130_fd_sc_hd__a31o_1 _10771_ (.A1(\div_shifter[43] ),
    .A2(net248),
    .A3(_03849_),
    .B1(net250),
    .X(_03851_));
 sky130_fd_sc_hd__o2bb2a_1 _10772_ (.A1_N(_06065_),
    .A2_N(_06459_),
    .B1(_03850_),
    .B2(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__o211a_1 _10773_ (.A1(_03845_),
    .A2(_03846_),
    .B1(_03848_),
    .C1(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__o21ai_2 _10774_ (.A1(net241),
    .A2(_02914_),
    .B1(_02272_),
    .Y(_03854_));
 sky130_fd_sc_hd__o221ai_1 _10775_ (.A1(net188),
    .A2(_03842_),
    .B1(_03854_),
    .B2(net190),
    .C1(_03853_),
    .Y(_03855_));
 sky130_fd_sc_hd__a211o_1 _10776_ (.A1(net216),
    .A2(_03843_),
    .B1(_03855_),
    .C1(_03833_),
    .X(_03856_));
 sky130_fd_sc_hd__a311o_1 _10777_ (.A1(net252),
    .A2(_03828_),
    .A3(_03829_),
    .B1(_03856_),
    .C1(_03827_),
    .X(_03857_));
 sky130_fd_sc_hd__a31o_1 _10778_ (.A1(curr_PC[9]),
    .A2(curr_PC[10]),
    .A3(_03486_),
    .B1(curr_PC[11]),
    .X(_03858_));
 sky130_fd_sc_hd__and4_1 _10779_ (.A(curr_PC[9]),
    .B(curr_PC[10]),
    .C(curr_PC[11]),
    .D(_03486_),
    .X(_03859_));
 sky130_fd_sc_hd__nor2_1 _10780_ (.A(net262),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__a22o_4 _10781_ (.A1(net262),
    .A2(_03857_),
    .B1(_03858_),
    .B2(_03860_),
    .X(dest_val[11]));
 sky130_fd_sc_hd__and2_1 _10782_ (.A(_03739_),
    .B(_03824_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_1 _10783_ (.A(net155),
    .B(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__o22a_1 _10784_ (.A1(net68),
    .A2(net59),
    .B1(net57),
    .B2(net94),
    .X(_03863_));
 sky130_fd_sc_hd__xnor2_1 _10785_ (.A(net100),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__o32a_1 _10786_ (.A1(_00176_),
    .A2(_00177_),
    .A3(net45),
    .B1(net54),
    .B2(net66),
    .X(_03865_));
 sky130_fd_sc_hd__xnor2_1 _10787_ (.A(net102),
    .B(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _10788_ (.A(_03864_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__xor2_1 _10789_ (.A(_03864_),
    .B(_03866_),
    .X(_03868_));
 sky130_fd_sc_hd__o22a_1 _10790_ (.A1(net64),
    .A2(net61),
    .B1(net50),
    .B2(net20),
    .X(_03869_));
 sky130_fd_sc_hd__xnor2_1 _10791_ (.A(net91),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _10792_ (.A(_03868_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__xor2_1 _10793_ (.A(_03868_),
    .B(_03870_),
    .X(_03872_));
 sky130_fd_sc_hd__o22a_1 _10794_ (.A1(net113),
    .A2(net15),
    .B1(net37),
    .B2(net123),
    .X(_03873_));
 sky130_fd_sc_hd__xnor2_1 _10795_ (.A(net77),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__a21oi_1 _10796_ (.A1(_00599_),
    .A2(_00600_),
    .B1(_00269_),
    .Y(_03875_));
 sky130_fd_sc_hd__nor2_1 _10797_ (.A(net117),
    .B(net10),
    .Y(_03876_));
 sky130_fd_sc_hd__o21a_1 _10798_ (.A1(_03875_),
    .A2(_03876_),
    .B1(net33),
    .X(_03877_));
 sky130_fd_sc_hd__nor3_1 _10799_ (.A(net33),
    .B(_03875_),
    .C(_03876_),
    .Y(_03878_));
 sky130_fd_sc_hd__or3_2 _10800_ (.A(_03874_),
    .B(_03877_),
    .C(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__o21ai_1 _10801_ (.A1(_03877_),
    .A2(_03878_),
    .B1(_03874_),
    .Y(_03880_));
 sky130_fd_sc_hd__and3_1 _10802_ (.A(_03872_),
    .B(_03879_),
    .C(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__a21o_1 _10803_ (.A1(_03879_),
    .A2(_03880_),
    .B1(_03872_),
    .X(_03882_));
 sky130_fd_sc_hd__inv_2 _10804_ (.A(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__o22a_1 _10805_ (.A1(net72),
    .A2(net48),
    .B1(net39),
    .B2(net25),
    .X(_03884_));
 sky130_fd_sc_hd__xnor2_1 _10806_ (.A(net105),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__o22a_1 _10807_ (.A1(net119),
    .A2(net29),
    .B1(net27),
    .B2(net85),
    .X(_03886_));
 sky130_fd_sc_hd__xnor2_1 _10808_ (.A(net111),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__and2_1 _10809_ (.A(_03885_),
    .B(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__xor2_1 _10810_ (.A(_03885_),
    .B(_03887_),
    .X(_03889_));
 sky130_fd_sc_hd__o22a_1 _10811_ (.A1(net23),
    .A2(net80),
    .B1(net42),
    .B2(net70),
    .X(_03890_));
 sky130_fd_sc_hd__xnor2_1 _10812_ (.A(net108),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__xor2_1 _10813_ (.A(_03889_),
    .B(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__and3b_1 _10814_ (.A_N(_03881_),
    .B(_03882_),
    .C(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__o21ba_1 _10815_ (.A1(_03881_),
    .A2(_03883_),
    .B1_N(_03892_),
    .X(_03894_));
 sky130_fd_sc_hd__o21ai_1 _10816_ (.A1(_06470_),
    .A2(_03789_),
    .B1(_03791_),
    .Y(_03895_));
 sky130_fd_sc_hd__a21o_1 _10817_ (.A1(_03757_),
    .A2(_03759_),
    .B1(_03755_),
    .X(_03896_));
 sky130_fd_sc_hd__or2_1 _10818_ (.A(net96),
    .B(net32),
    .X(_03897_));
 sky130_fd_sc_hd__nand2b_1 _10819_ (.A_N(_03897_),
    .B(_03896_),
    .Y(_03898_));
 sky130_fd_sc_hd__xnor2_1 _10820_ (.A(_03896_),
    .B(_03897_),
    .Y(_03899_));
 sky130_fd_sc_hd__xnor2_1 _10821_ (.A(_03895_),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__or3_1 _10822_ (.A(_03893_),
    .B(_03894_),
    .C(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__inv_2 _10823_ (.A(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__o21a_1 _10824_ (.A1(_03893_),
    .A2(_03894_),
    .B1(_03900_),
    .X(_03903_));
 sky130_fd_sc_hd__nor2_1 _10825_ (.A(_03902_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__o21bai_1 _10826_ (.A1(_03743_),
    .A2(_03744_),
    .B1_N(_03749_),
    .Y(_03905_));
 sky130_fd_sc_hd__o22a_1 _10827_ (.A1(net74),
    .A2(net18),
    .B1(net13),
    .B2(net115),
    .X(_03906_));
 sky130_fd_sc_hd__xnor2_1 _10828_ (.A(_06499_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__o21ba_1 _10829_ (.A1(_06475_),
    .A2(net6),
    .B1_N(net153),
    .X(_03908_));
 sky130_fd_sc_hd__a31o_1 _10830_ (.A1(net153),
    .A2(_06473_),
    .A3(_00510_),
    .B1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__nor2_1 _10831_ (.A(_03907_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__and2_1 _10832_ (.A(_03907_),
    .B(_03909_),
    .X(_03911_));
 sky130_fd_sc_hd__or2_1 _10833_ (.A(_03910_),
    .B(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__o21ai_1 _10834_ (.A1(_03768_),
    .A2(_03772_),
    .B1(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__or3_1 _10835_ (.A(_03768_),
    .B(_03772_),
    .C(_03912_),
    .X(_03914_));
 sky130_fd_sc_hd__and2_1 _10836_ (.A(_03913_),
    .B(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__nand2_1 _10837_ (.A(_03905_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__xnor2_1 _10838_ (.A(_03905_),
    .B(_03915_),
    .Y(_03917_));
 sky130_fd_sc_hd__xnor2_1 _10839_ (.A(_03904_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a21bo_1 _10840_ (.A1(_03783_),
    .A2(_03796_),
    .B1_N(_03782_),
    .X(_03919_));
 sky130_fd_sc_hd__a21bo_1 _10841_ (.A1(_03792_),
    .A2(_03793_),
    .B1_N(_03795_),
    .X(_03920_));
 sky130_fd_sc_hd__a21oi_1 _10842_ (.A1(_03777_),
    .A2(_03780_),
    .B1(_03779_),
    .Y(_03921_));
 sky130_fd_sc_hd__o21ba_1 _10843_ (.A1(_03761_),
    .A2(_03775_),
    .B1_N(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__or3b_1 _10844_ (.A(_03761_),
    .B(_03775_),
    .C_N(_03921_),
    .X(_03923_));
 sky130_fd_sc_hd__and2b_1 _10845_ (.A_N(_03922_),
    .B(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__xnor2_1 _10846_ (.A(_03920_),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__a21oi_1 _10847_ (.A1(_03800_),
    .A2(_03804_),
    .B1(_03803_),
    .Y(_03926_));
 sky130_fd_sc_hd__xnor2_1 _10848_ (.A(_03925_),
    .B(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2b_1 _10849_ (.A_N(_03927_),
    .B(_03919_),
    .Y(_03928_));
 sky130_fd_sc_hd__xnor2_1 _10850_ (.A(_03919_),
    .B(_03927_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _10851_ (.A(_03918_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__xor2_1 _10852_ (.A(_03918_),
    .B(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__o21ai_2 _10853_ (.A1(_03806_),
    .A2(_03808_),
    .B1(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__or3_1 _10854_ (.A(_03806_),
    .B(_03808_),
    .C(_03931_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_2 _10855_ (.A(_03932_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand2_2 _10856_ (.A(_03810_),
    .B(_03812_),
    .Y(_03935_));
 sky130_fd_sc_hd__nand2b_1 _10857_ (.A_N(_03934_),
    .B(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__and3_1 _10858_ (.A(_03810_),
    .B(_03812_),
    .C(_03934_),
    .X(_03937_));
 sky130_fd_sc_hd__xor2_4 _10859_ (.A(_03934_),
    .B(_03935_),
    .X(_03938_));
 sky130_fd_sc_hd__nor2_1 _10860_ (.A(_03696_),
    .B(_03817_),
    .Y(_03939_));
 sky130_fd_sc_hd__and4b_1 _10861_ (.A_N(_03575_),
    .B(_03939_),
    .C(_03445_),
    .D(_03446_),
    .X(_03940_));
 sky130_fd_sc_hd__inv_2 _10862_ (.A(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__a211o_1 _10863_ (.A1(_02794_),
    .A2(_02796_),
    .B1(_03451_),
    .C1(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__or2_1 _10864_ (.A(_03450_),
    .B(_03941_),
    .X(_03943_));
 sky130_fd_sc_hd__a21oi_1 _10865_ (.A1(_03694_),
    .A2(_03815_),
    .B1(_03816_),
    .Y(_03944_));
 sky130_fd_sc_hd__inv_2 _10866_ (.A(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__a21o_1 _10867_ (.A1(_03700_),
    .A2(_03939_),
    .B1(_03944_),
    .X(_03946_));
 sky130_fd_sc_hd__inv_2 _10868_ (.A(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__a31o_1 _10869_ (.A1(_03942_),
    .A2(_03943_),
    .A3(_03947_),
    .B1(_03938_),
    .X(_03948_));
 sky130_fd_sc_hd__nand4_1 _10870_ (.A(_03938_),
    .B(_03942_),
    .C(_03943_),
    .D(_03947_),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_2 _10871_ (.A(_03948_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__o21ai_1 _10872_ (.A1(_03862_),
    .A2(_03950_),
    .B1(_02171_),
    .Y(_03951_));
 sky130_fd_sc_hd__a21oi_1 _10873_ (.A1(_03862_),
    .A2(_03950_),
    .B1(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__o21ai_1 _10874_ (.A1(net156),
    .A2(_02098_),
    .B1(_02099_),
    .Y(_03953_));
 sky130_fd_sc_hd__o31a_1 _10875_ (.A1(net156),
    .A2(_02098_),
    .A3(_02099_),
    .B1(net252),
    .X(_03954_));
 sky130_fd_sc_hd__a21o_1 _10876_ (.A1(_06102_),
    .A2(_03830_),
    .B1(_06087_),
    .X(_03955_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(_06363_),
    .A1(_03955_),
    .S(net303),
    .X(_03956_));
 sky130_fd_sc_hd__nand2_1 _10878_ (.A(_06043_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__or2_1 _10879_ (.A(_06043_),
    .B(_03956_),
    .X(_03958_));
 sky130_fd_sc_hd__or2_1 _10880_ (.A(net238),
    .B(_02913_),
    .X(_03959_));
 sky130_fd_sc_hd__o211a_1 _10881_ (.A1(net237),
    .A2(_02910_),
    .B1(_03959_),
    .C1(net239),
    .X(_03960_));
 sky130_fd_sc_hd__a21oi_2 _10882_ (.A1(net241),
    .A2(_02769_),
    .B1(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__inv_2 _10883_ (.A(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__or2_1 _10884_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .X(_03963_));
 sky130_fd_sc_hd__nand2_1 _10885_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .Y(_03964_));
 sky130_fd_sc_hd__o211a_1 _10886_ (.A1(_03835_),
    .A2(_03838_),
    .B1(_03963_),
    .C1(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__a211o_1 _10887_ (.A1(_03963_),
    .A2(_03964_),
    .B1(_03835_),
    .C1(_03838_),
    .X(_03966_));
 sky130_fd_sc_hd__or3b_1 _10888_ (.A(net243),
    .B(_03965_),
    .C_N(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__o21ai_1 _10889_ (.A1(net268),
    .A2(_03961_),
    .B1(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__or2_1 _10890_ (.A(\div_res[11] ),
    .B(_03844_),
    .X(_03969_));
 sky130_fd_sc_hd__a21o_1 _10891_ (.A1(net163),
    .A2(_03969_),
    .B1(\div_res[12] ),
    .X(_03970_));
 sky130_fd_sc_hd__a31oi_1 _10892_ (.A1(\div_res[12] ),
    .A2(net163),
    .A3(_03969_),
    .B1(net204),
    .Y(_03971_));
 sky130_fd_sc_hd__or2_1 _10893_ (.A(\div_shifter[43] ),
    .B(_03849_),
    .X(_03972_));
 sky130_fd_sc_hd__a21oi_1 _10894_ (.A1(net248),
    .A2(_03972_),
    .B1(\div_shifter[44] ),
    .Y(_03973_));
 sky130_fd_sc_hd__a31o_1 _10895_ (.A1(\div_shifter[44] ),
    .A2(net248),
    .A3(_03972_),
    .B1(net250),
    .X(_03974_));
 sky130_fd_sc_hd__nor2_2 _10896_ (.A(_03973_),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(net253),
    .A1(net206),
    .S(_06021_),
    .X(_03976_));
 sky130_fd_sc_hd__a21oi_1 _10898_ (.A1(net207),
    .A2(_03976_),
    .B1(_06032_),
    .Y(_03977_));
 sky130_fd_sc_hd__a211o_1 _10899_ (.A1(_05999_),
    .A2(_06459_),
    .B1(_03975_),
    .C1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__o21a_1 _10900_ (.A1(net240),
    .A2(_02759_),
    .B1(_02272_),
    .X(_03979_));
 sky130_fd_sc_hd__inv_2 _10901_ (.A(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__a221o_1 _10902_ (.A1(_03970_),
    .A2(_03971_),
    .B1(_03979_),
    .B2(net192),
    .C1(_03978_),
    .X(_03981_));
 sky130_fd_sc_hd__a221o_1 _10903_ (.A1(_02243_),
    .A2(_03962_),
    .B1(_03968_),
    .B2(net216),
    .C1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__a31o_1 _10904_ (.A1(_02247_),
    .A2(_03957_),
    .A3(_03958_),
    .B1(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__a211o_1 _10905_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03983_),
    .C1(_03952_),
    .X(_03984_));
 sky130_fd_sc_hd__and2_1 _10906_ (.A(curr_PC[12]),
    .B(_03859_),
    .X(_03985_));
 sky130_fd_sc_hd__o21ai_1 _10907_ (.A1(curr_PC[12]),
    .A2(_03859_),
    .B1(net267),
    .Y(_03986_));
 sky130_fd_sc_hd__a2bb2o_4 _10908_ (.A1_N(_03985_),
    .A2_N(_03986_),
    .B1(net262),
    .B2(_03984_),
    .X(dest_val[12]));
 sky130_fd_sc_hd__a31o_1 _10909_ (.A1(_03739_),
    .A2(_03824_),
    .A3(_03950_),
    .B1(net156),
    .X(_03987_));
 sky130_fd_sc_hd__o21ai_1 _10910_ (.A1(_03925_),
    .A2(_03926_),
    .B1(_03928_),
    .Y(_03988_));
 sky130_fd_sc_hd__a21oi_1 _10911_ (.A1(_03889_),
    .A2(_03891_),
    .B1(_03888_),
    .Y(_03989_));
 sky130_fd_sc_hd__a21o_1 _10912_ (.A1(_03867_),
    .A2(_03871_),
    .B1(_03879_),
    .X(_03990_));
 sky130_fd_sc_hd__nand3_1 _10913_ (.A(_03867_),
    .B(_03871_),
    .C(_03879_),
    .Y(_03991_));
 sky130_fd_sc_hd__and2_1 _10914_ (.A(_03990_),
    .B(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__nand2b_1 _10915_ (.A_N(_03989_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__xnor2_1 _10916_ (.A(_03989_),
    .B(_03992_),
    .Y(_03994_));
 sky130_fd_sc_hd__o22a_1 _10917_ (.A1(net20),
    .A2(net61),
    .B1(net59),
    .B2(net64),
    .X(_03995_));
 sky130_fd_sc_hd__xnor2_1 _10918_ (.A(net91),
    .B(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__o22a_1 _10919_ (.A1(net25),
    .A2(net48),
    .B1(net44),
    .B2(net72),
    .X(_03997_));
 sky130_fd_sc_hd__xnor2_1 _10920_ (.A(net105),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__and2_1 _10921_ (.A(_03996_),
    .B(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__nor2_1 _10922_ (.A(_03996_),
    .B(_03998_),
    .Y(_04000_));
 sky130_fd_sc_hd__nor2_1 _10923_ (.A(_03999_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__o22a_1 _10924_ (.A1(net22),
    .A2(net54),
    .B1(net51),
    .B2(net66),
    .X(_04002_));
 sky130_fd_sc_hd__xnor2_1 _10925_ (.A(net102),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xor2_1 _10926_ (.A(_04001_),
    .B(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__o32a_1 _10927_ (.A1(net124),
    .A2(_00351_),
    .A3(_00352_),
    .B1(net36),
    .B2(net120),
    .X(_04005_));
 sky130_fd_sc_hd__xnor2_1 _10928_ (.A(net77),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__a21o_1 _10929_ (.A1(_00137_),
    .A2(_00138_),
    .B1(net42),
    .X(_04007_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(net70),
    .B(net39),
    .X(_04008_));
 sky130_fd_sc_hd__nand3_1 _10931_ (.A(net109),
    .B(_04007_),
    .C(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__a21o_1 _10932_ (.A1(_04007_),
    .A2(_04008_),
    .B1(net109),
    .X(_04010_));
 sky130_fd_sc_hd__a21o_1 _10933_ (.A1(_04009_),
    .A2(_04010_),
    .B1(_04006_),
    .X(_04011_));
 sky130_fd_sc_hd__inv_2 _10934_ (.A(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__nand3_1 _10935_ (.A(_04006_),
    .B(_04009_),
    .C(_04010_),
    .Y(_04013_));
 sky130_fd_sc_hd__o22a_1 _10936_ (.A1(net30),
    .A2(net85),
    .B1(net80),
    .B2(net27),
    .X(_04014_));
 sky130_fd_sc_hd__xnor2_1 _10937_ (.A(net112),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__and3_1 _10938_ (.A(_04011_),
    .B(_04013_),
    .C(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__a21oi_1 _10939_ (.A1(_04011_),
    .A2(_04013_),
    .B1(_04015_),
    .Y(_04017_));
 sky130_fd_sc_hd__nor2_1 _10940_ (.A(_04016_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__or2_1 _10941_ (.A(net68),
    .B(net57),
    .X(_04019_));
 sky130_fd_sc_hd__a21o_1 _10942_ (.A1(_00243_),
    .A2(_00244_),
    .B1(net94),
    .X(_04020_));
 sky130_fd_sc_hd__nand3_1 _10943_ (.A(net100),
    .B(_04019_),
    .C(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21o_1 _10944_ (.A1(_04019_),
    .A2(_04020_),
    .B1(net100),
    .X(_04022_));
 sky130_fd_sc_hd__a21boi_1 _10945_ (.A1(_04021_),
    .A2(_04022_),
    .B1_N(net152),
    .Y(_04023_));
 sky130_fd_sc_hd__a21bo_1 _10946_ (.A1(_04021_),
    .A2(_04022_),
    .B1_N(net152),
    .X(_04024_));
 sky130_fd_sc_hd__nand3b_1 _10947_ (.A_N(net152),
    .B(_04021_),
    .C(_04022_),
    .Y(_04025_));
 sky130_fd_sc_hd__o22a_1 _10948_ (.A1(net74),
    .A2(net13),
    .B1(net6),
    .B2(net115),
    .X(_04026_));
 sky130_fd_sc_hd__xnor2_1 _10949_ (.A(net151),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__and3_1 _10950_ (.A(_04024_),
    .B(_04025_),
    .C(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__a21oi_1 _10951_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_04027_),
    .Y(_04029_));
 sky130_fd_sc_hd__nor2_1 _10952_ (.A(_04028_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _10953_ (.A(_04018_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__xor2_1 _10954_ (.A(_04018_),
    .B(_04030_),
    .X(_04032_));
 sky130_fd_sc_hd__nand2_1 _10955_ (.A(_04004_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__or2_1 _10956_ (.A(_04004_),
    .B(_04032_),
    .X(_04034_));
 sky130_fd_sc_hd__nand2_1 _10957_ (.A(_04033_),
    .B(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__o22a_1 _10958_ (.A1(net113),
    .A2(net10),
    .B1(net5),
    .B2(net117),
    .X(_04036_));
 sky130_fd_sc_hd__xnor2_1 _10959_ (.A(net33),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand2b_1 _10960_ (.A_N(_03910_),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__or3_1 _10961_ (.A(_03907_),
    .B(_03909_),
    .C(_04037_),
    .X(_04039_));
 sky130_fd_sc_hd__nand2_1 _10962_ (.A(_04038_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__or2_1 _10963_ (.A(net89),
    .B(net32),
    .X(_04041_));
 sky130_fd_sc_hd__xnor2_1 _10964_ (.A(_04040_),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__or2_1 _10965_ (.A(_04035_),
    .B(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__nand2_1 _10966_ (.A(_04035_),
    .B(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__and3_1 _10967_ (.A(_03994_),
    .B(_04043_),
    .C(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__a21oi_1 _10968_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_03994_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor2_1 _10969_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__o21ai_1 _10970_ (.A1(_03903_),
    .A2(_03917_),
    .B1(_03901_),
    .Y(_04048_));
 sky130_fd_sc_hd__nor2_1 _10971_ (.A(_03881_),
    .B(_03893_),
    .Y(_04049_));
 sky130_fd_sc_hd__a21boi_1 _10972_ (.A1(_03895_),
    .A2(_03899_),
    .B1_N(_03898_),
    .Y(_04050_));
 sky130_fd_sc_hd__or2_1 _10973_ (.A(_04049_),
    .B(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__xnor2_1 _10974_ (.A(_04049_),
    .B(_04050_),
    .Y(_04052_));
 sky130_fd_sc_hd__a21o_1 _10975_ (.A1(_03913_),
    .A2(_03916_),
    .B1(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__nand3_1 _10976_ (.A(_03913_),
    .B(_03916_),
    .C(_04052_),
    .Y(_04054_));
 sky130_fd_sc_hd__nand2_1 _10977_ (.A(_04053_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__a21oi_1 _10978_ (.A1(_03920_),
    .A2(_03923_),
    .B1(_03922_),
    .Y(_04056_));
 sky130_fd_sc_hd__xnor2_1 _10979_ (.A(_04055_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__and2b_1 _10980_ (.A_N(_04057_),
    .B(_04048_),
    .X(_04058_));
 sky130_fd_sc_hd__xnor2_1 _10981_ (.A(_04048_),
    .B(_04057_),
    .Y(_04059_));
 sky130_fd_sc_hd__and2_1 _10982_ (.A(_04047_),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__xnor2_1 _10983_ (.A(_04047_),
    .B(_04059_),
    .Y(_04061_));
 sky130_fd_sc_hd__and2b_1 _10984_ (.A_N(_04061_),
    .B(_03988_),
    .X(_04062_));
 sky130_fd_sc_hd__xor2_1 _10985_ (.A(_03988_),
    .B(_04061_),
    .X(_04063_));
 sky130_fd_sc_hd__a21o_1 _10986_ (.A1(_03930_),
    .A2(_03932_),
    .B1(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__nand3_2 _10987_ (.A(_03930_),
    .B(_03932_),
    .C(_04063_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_2 _10988_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__a21oi_1 _10989_ (.A1(_03815_),
    .A2(_03936_),
    .B1(_03937_),
    .Y(_04067_));
 sky130_fd_sc_hd__or2_1 _10990_ (.A(_03817_),
    .B(_03938_),
    .X(_04068_));
 sky130_fd_sc_hd__o21ba_1 _10991_ (.A1(_03818_),
    .A2(_04068_),
    .B1_N(_04067_),
    .X(_04069_));
 sky130_fd_sc_hd__or2_1 _10992_ (.A(_03819_),
    .B(_04068_),
    .X(_04070_));
 sky130_fd_sc_hd__a31o_1 _10993_ (.A1(_03577_),
    .A2(_03579_),
    .A3(_03580_),
    .B1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__a21o_1 _10994_ (.A1(_04069_),
    .A2(_04071_),
    .B1(_04066_),
    .X(_04072_));
 sky130_fd_sc_hd__nand3_1 _10995_ (.A(_04066_),
    .B(_04069_),
    .C(_04071_),
    .Y(_04073_));
 sky130_fd_sc_hd__nand2_2 _10996_ (.A(_04072_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__a21oi_1 _10997_ (.A1(_03987_),
    .A2(_04074_),
    .B1(net209),
    .Y(_04075_));
 sky130_fd_sc_hd__o21a_1 _10998_ (.A1(_03987_),
    .A2(_04074_),
    .B1(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__or3_1 _10999_ (.A(net155),
    .B(_02100_),
    .C(_02106_),
    .X(_04077_));
 sky130_fd_sc_hd__o21ai_1 _11000_ (.A1(net155),
    .A2(_02100_),
    .B1(_02106_),
    .Y(_04078_));
 sky130_fd_sc_hd__a21o_1 _11001_ (.A1(_06043_),
    .A2(_03955_),
    .B1(_06021_),
    .X(_04079_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(_06364_),
    .A1(_04079_),
    .S(net303),
    .X(_04080_));
 sky130_fd_sc_hd__nand2_1 _11003_ (.A(_05979_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__or2_1 _11004_ (.A(_05979_),
    .B(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__or2_1 _11005_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .X(_04083_));
 sky130_fd_sc_hd__nand2_1 _11006_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _11007_ (.A(_04083_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__a21oi_1 _11008_ (.A1(reg1_val[12]),
    .A2(curr_PC[12]),
    .B1(_03965_),
    .Y(_04086_));
 sky130_fd_sc_hd__xor2_1 _11009_ (.A(_04085_),
    .B(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(_03057_),
    .A1(_03061_),
    .S(net236),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_2 _11011_ (.A0(_02585_),
    .A1(_04088_),
    .S(net239),
    .X(_04089_));
 sky130_fd_sc_hd__nand2_1 _11012_ (.A(net244),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__o211a_1 _11013_ (.A1(net243),
    .A2(_04087_),
    .B1(_04090_),
    .C1(net216),
    .X(_04091_));
 sky130_fd_sc_hd__or2_1 _11014_ (.A(\div_res[12] ),
    .B(_03969_),
    .X(_04092_));
 sky130_fd_sc_hd__a21oi_1 _11015_ (.A1(net163),
    .A2(_04092_),
    .B1(\div_res[13] ),
    .Y(_04093_));
 sky130_fd_sc_hd__a31o_1 _11016_ (.A1(\div_res[13] ),
    .A2(net163),
    .A3(_04092_),
    .B1(net204),
    .X(_04094_));
 sky130_fd_sc_hd__or2_1 _11017_ (.A(\div_shifter[44] ),
    .B(_03972_),
    .X(_04095_));
 sky130_fd_sc_hd__a21oi_1 _11018_ (.A1(net248),
    .A2(_04095_),
    .B1(\div_shifter[45] ),
    .Y(_04096_));
 sky130_fd_sc_hd__a31o_1 _11019_ (.A1(\div_shifter[45] ),
    .A2(net248),
    .A3(_04095_),
    .B1(net250),
    .X(_04097_));
 sky130_fd_sc_hd__nand2_1 _11020_ (.A(_05955_),
    .B(_06459_),
    .Y(_04098_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(net253),
    .A1(net206),
    .S(_05967_),
    .X(_04099_));
 sky130_fd_sc_hd__a21o_1 _11022_ (.A1(net207),
    .A2(_04099_),
    .B1(_05973_),
    .X(_04100_));
 sky130_fd_sc_hd__o211a_1 _11023_ (.A1(_04096_),
    .A2(_04097_),
    .B1(_04098_),
    .C1(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__o21ai_2 _11024_ (.A1(net240),
    .A2(_02599_),
    .B1(_02272_),
    .Y(_04102_));
 sky130_fd_sc_hd__o221a_1 _11025_ (.A1(_04093_),
    .A2(_04094_),
    .B1(_04102_),
    .B2(net190),
    .C1(_04101_),
    .X(_04103_));
 sky130_fd_sc_hd__o21ai_1 _11026_ (.A1(net188),
    .A2(_04089_),
    .B1(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__a311o_1 _11027_ (.A1(_02247_),
    .A2(_04081_),
    .A3(_04082_),
    .B1(_04091_),
    .C1(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__a311o_1 _11028_ (.A1(net252),
    .A2(_04077_),
    .A3(_04078_),
    .B1(_04105_),
    .C1(_04076_),
    .X(_04106_));
 sky130_fd_sc_hd__or2_1 _11029_ (.A(curr_PC[13]),
    .B(_03985_),
    .X(_04107_));
 sky130_fd_sc_hd__a21oi_1 _11030_ (.A1(curr_PC[13]),
    .A2(_03985_),
    .B1(net262),
    .Y(_04108_));
 sky130_fd_sc_hd__a22o_4 _11031_ (.A1(net263),
    .A2(_04106_),
    .B1(_04107_),
    .B2(_04108_),
    .X(dest_val[13]));
 sky130_fd_sc_hd__a22o_1 _11032_ (.A1(_03948_),
    .A2(_03949_),
    .B1(_04072_),
    .B2(_04073_),
    .X(_04109_));
 sky130_fd_sc_hd__or4_2 _11033_ (.A(_03358_),
    .B(_03738_),
    .C(_03825_),
    .D(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__nand2_1 _11034_ (.A(net160),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__o22a_1 _11035_ (.A1(net29),
    .A2(net79),
    .B1(net42),
    .B2(net27),
    .X(_04112_));
 sky130_fd_sc_hd__xnor2_1 _11036_ (.A(net111),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__o22a_1 _11037_ (.A1(net70),
    .A2(net48),
    .B1(net39),
    .B2(net23),
    .X(_04114_));
 sky130_fd_sc_hd__xnor2_1 _11038_ (.A(net109),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__and2_1 _11039_ (.A(_04113_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__xnor2_1 _11040_ (.A(_04113_),
    .B(_04115_),
    .Y(_04117_));
 sky130_fd_sc_hd__o22a_1 _11041_ (.A1(net68),
    .A2(net17),
    .B1(net12),
    .B2(net94),
    .X(_04118_));
 sky130_fd_sc_hd__xnor2_1 _11042_ (.A(net100),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__a31o_1 _11043_ (.A1(net152),
    .A2(_06503_),
    .A3(_00510_),
    .B1(net149),
    .X(_04120_));
 sky130_fd_sc_hd__o21a_1 _11044_ (.A1(_06504_),
    .A2(net8),
    .B1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__and2b_1 _11045_ (.A_N(_04119_),
    .B(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__xnor2_1 _11046_ (.A(_04119_),
    .B(_04121_),
    .Y(_04123_));
 sky130_fd_sc_hd__nor2_1 _11047_ (.A(_04117_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _11048_ (.A(_04117_),
    .B(_04123_),
    .Y(_04125_));
 sky130_fd_sc_hd__and2b_1 _11049_ (.A_N(_04124_),
    .B(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__o22a_1 _11050_ (.A1(net20),
    .A2(net58),
    .B1(net56),
    .B2(net64),
    .X(_04127_));
 sky130_fd_sc_hd__xnor2_1 _11051_ (.A(net91),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__o22a_1 _11052_ (.A1(net72),
    .A2(net53),
    .B1(net45),
    .B2(net25),
    .X(_04129_));
 sky130_fd_sc_hd__xnor2_1 _11053_ (.A(net105),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__and2_1 _11054_ (.A(_04128_),
    .B(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__nor2_1 _11055_ (.A(_04128_),
    .B(_04130_),
    .Y(_04132_));
 sky130_fd_sc_hd__nor2_1 _11056_ (.A(_04131_),
    .B(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__o22a_1 _11057_ (.A1(net66),
    .A2(net61),
    .B1(net50),
    .B2(_00178_),
    .X(_04134_));
 sky130_fd_sc_hd__xnor2_1 _11058_ (.A(net102),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__xor2_1 _11059_ (.A(_04133_),
    .B(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__and2_1 _11060_ (.A(_04126_),
    .B(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__nor2_1 _11061_ (.A(_04126_),
    .B(_04136_),
    .Y(_04138_));
 sky130_fd_sc_hd__or2_1 _11062_ (.A(_04137_),
    .B(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__o22a_1 _11063_ (.A1(net123),
    .A2(net9),
    .B1(net4),
    .B2(net113),
    .X(_04140_));
 sky130_fd_sc_hd__xnor2_1 _11064_ (.A(net34),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__or2_1 _11065_ (.A(net117),
    .B(_00596_),
    .X(_04142_));
 sky130_fd_sc_hd__o22a_1 _11066_ (.A1(net119),
    .A2(net15),
    .B1(net36),
    .B2(net85),
    .X(_04143_));
 sky130_fd_sc_hd__xnor2_1 _11067_ (.A(_00348_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__and2b_1 _11068_ (.A_N(_04142_),
    .B(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__xnor2_1 _11069_ (.A(_04142_),
    .B(_04144_),
    .Y(_04146_));
 sky130_fd_sc_hd__xnor2_1 _11070_ (.A(_04141_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__nor2_1 _11071_ (.A(_04139_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__and2_1 _11072_ (.A(_04139_),
    .B(_04147_),
    .X(_04149_));
 sky130_fd_sc_hd__nor2_1 _11073_ (.A(_04148_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21o_1 _11074_ (.A1(_04001_),
    .A2(_04003_),
    .B1(_03999_),
    .X(_04151_));
 sky130_fd_sc_hd__o22a_1 _11075_ (.A1(_04012_),
    .A2(_04016_),
    .B1(_04023_),
    .B2(_04028_),
    .X(_04152_));
 sky130_fd_sc_hd__or4_1 _11076_ (.A(_04012_),
    .B(_04016_),
    .C(_04023_),
    .D(_04028_),
    .X(_04153_));
 sky130_fd_sc_hd__and2b_1 _11077_ (.A_N(_04152_),
    .B(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__xor2_1 _11078_ (.A(_04151_),
    .B(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__xnor2_1 _11079_ (.A(_04150_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__a21bo_1 _11080_ (.A1(_03994_),
    .A2(_04044_),
    .B1_N(_04043_),
    .X(_04157_));
 sky130_fd_sc_hd__nand2_1 _11081_ (.A(_03990_),
    .B(_03993_),
    .Y(_04158_));
 sky130_fd_sc_hd__a21bo_1 _11082_ (.A1(_04004_),
    .A2(_04032_),
    .B1_N(_04031_),
    .X(_04159_));
 sky130_fd_sc_hd__o21a_1 _11083_ (.A1(_04040_),
    .A2(_04041_),
    .B1(_04038_),
    .X(_04160_));
 sky130_fd_sc_hd__a21o_1 _11084_ (.A1(_04031_),
    .A2(_04033_),
    .B1(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__xnor2_1 _11085_ (.A(_04159_),
    .B(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__xnor2_1 _11086_ (.A(_04158_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_1 _11087_ (.A1(_04051_),
    .A2(_04053_),
    .B1(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__and3_1 _11088_ (.A(_04051_),
    .B(_04053_),
    .C(_04163_),
    .X(_04165_));
 sky130_fd_sc_hd__nor2_1 _11089_ (.A(_04164_),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__xnor2_1 _11090_ (.A(_04157_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__or2_1 _11091_ (.A(_04156_),
    .B(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__xor2_1 _11092_ (.A(_04156_),
    .B(_04167_),
    .X(_04169_));
 sky130_fd_sc_hd__o21ba_1 _11093_ (.A1(_04055_),
    .A2(_04056_),
    .B1_N(_04058_),
    .X(_04170_));
 sky130_fd_sc_hd__nand2b_1 _11094_ (.A_N(_04170_),
    .B(_04169_),
    .Y(_04171_));
 sky130_fd_sc_hd__xnor2_1 _11095_ (.A(_04169_),
    .B(_04170_),
    .Y(_04172_));
 sky130_fd_sc_hd__o21ai_2 _11096_ (.A1(_04060_),
    .A2(_04062_),
    .B1(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__or3_1 _11097_ (.A(_04060_),
    .B(_04062_),
    .C(_04172_),
    .X(_04174_));
 sky130_fd_sc_hd__and2_2 _11098_ (.A(_04173_),
    .B(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__a21bo_1 _11099_ (.A1(_03936_),
    .A2(_04064_),
    .B1_N(_04065_),
    .X(_04176_));
 sky130_fd_sc_hd__or2_1 _11100_ (.A(_03938_),
    .B(_04066_),
    .X(_04177_));
 sky130_fd_sc_hd__o21ai_1 _11101_ (.A1(_03945_),
    .A2(_04177_),
    .B1(_04176_),
    .Y(_04178_));
 sky130_fd_sc_hd__nor3_1 _11102_ (.A(_03696_),
    .B(_03817_),
    .C(_04177_),
    .Y(_04179_));
 sky130_fd_sc_hd__a21oi_2 _11103_ (.A1(_03702_),
    .A2(_04179_),
    .B1(_04178_),
    .Y(_04180_));
 sky130_fd_sc_hd__xor2_4 _11104_ (.A(_04175_),
    .B(_04180_),
    .X(_04181_));
 sky130_fd_sc_hd__o21ai_1 _11105_ (.A1(_04111_),
    .A2(_04181_),
    .B1(_02171_),
    .Y(_04182_));
 sky130_fd_sc_hd__a21oi_1 _11106_ (.A1(_04111_),
    .A2(_04181_),
    .B1(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__or3_1 _11107_ (.A(net156),
    .B(_02107_),
    .C(_02108_),
    .X(_04184_));
 sky130_fd_sc_hd__o21ai_1 _11108_ (.A1(net156),
    .A2(_02107_),
    .B1(_02108_),
    .Y(_04185_));
 sky130_fd_sc_hd__a21o_1 _11109_ (.A1(_05979_),
    .A2(_04079_),
    .B1(_05967_),
    .X(_04186_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(_06365_),
    .A1(_04186_),
    .S(net303),
    .X(_04187_));
 sky130_fd_sc_hd__nand2_1 _11111_ (.A(_05943_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__o211a_1 _11112_ (.A1(_05943_),
    .A2(_04187_),
    .B1(_04188_),
    .C1(_02247_),
    .X(_04189_));
 sky130_fd_sc_hd__or2_1 _11113_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .X(_04190_));
 sky130_fd_sc_hd__nand2_1 _11114_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _11115_ (.A(_04190_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__o21a_1 _11116_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_04084_),
    .X(_04193_));
 sky130_fd_sc_hd__xor2_1 _11117_ (.A(_04192_),
    .B(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__or2_1 _11118_ (.A(net238),
    .B(_03202_),
    .X(_04195_));
 sky130_fd_sc_hd__o211a_1 _11119_ (.A1(net236),
    .A2(_03200_),
    .B1(_04195_),
    .C1(net239),
    .X(_04196_));
 sky130_fd_sc_hd__a21oi_2 _11120_ (.A1(net240),
    .A2(_02458_),
    .B1(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _11121_ (.A(net244),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__o211a_1 _11122_ (.A1(net243),
    .A2(_04194_),
    .B1(_04198_),
    .C1(net216),
    .X(_04199_));
 sky130_fd_sc_hd__or2_1 _11123_ (.A(\div_shifter[45] ),
    .B(_04095_),
    .X(_04200_));
 sky130_fd_sc_hd__a21oi_1 _11124_ (.A1(net249),
    .A2(_04200_),
    .B1(\div_shifter[46] ),
    .Y(_04201_));
 sky130_fd_sc_hd__a31o_1 _11125_ (.A1(\div_shifter[46] ),
    .A2(net249),
    .A3(_04200_),
    .B1(net251),
    .X(_04202_));
 sky130_fd_sc_hd__or2_2 _11126_ (.A(_04201_),
    .B(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__or2_1 _11127_ (.A(\div_res[13] ),
    .B(_04092_),
    .X(_04204_));
 sky130_fd_sc_hd__a21oi_1 _11128_ (.A1(net162),
    .A2(_04204_),
    .B1(\div_res[14] ),
    .Y(_04205_));
 sky130_fd_sc_hd__a31o_1 _11129_ (.A1(\div_res[14] ),
    .A2(net162),
    .A3(_04204_),
    .B1(net204),
    .X(_04206_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(net253),
    .A1(net206),
    .S(_05925_),
    .X(_04207_));
 sky130_fd_sc_hd__a21oi_1 _11131_ (.A1(net207),
    .A2(_04207_),
    .B1(_05934_),
    .Y(_04208_));
 sky130_fd_sc_hd__a21oi_1 _11132_ (.A1(_05907_),
    .A2(_06459_),
    .B1(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__o211a_1 _11133_ (.A1(_04205_),
    .A2(_04206_),
    .B1(_04209_),
    .C1(_04203_),
    .X(_04210_));
 sky130_fd_sc_hd__o21a_1 _11134_ (.A1(net240),
    .A2(_02429_),
    .B1(_02272_),
    .X(_04211_));
 sky130_fd_sc_hd__inv_2 _11135_ (.A(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__o221a_1 _11136_ (.A1(net188),
    .A2(_04197_),
    .B1(_04212_),
    .B2(net190),
    .C1(_04210_),
    .X(_04213_));
 sky130_fd_sc_hd__or3b_1 _11137_ (.A(_04189_),
    .B(_04199_),
    .C_N(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__a311o_1 _11138_ (.A1(net252),
    .A2(_04184_),
    .A3(_04185_),
    .B1(_04214_),
    .C1(_04183_),
    .X(_04215_));
 sky130_fd_sc_hd__and3_1 _11139_ (.A(curr_PC[13]),
    .B(curr_PC[14]),
    .C(_03985_),
    .X(_04216_));
 sky130_fd_sc_hd__a21oi_1 _11140_ (.A1(curr_PC[13]),
    .A2(_03985_),
    .B1(curr_PC[14]),
    .Y(_04217_));
 sky130_fd_sc_hd__nor2_1 _11141_ (.A(_04216_),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__mux2_8 _11142_ (.A0(_04215_),
    .A1(_04218_),
    .S(net267),
    .X(dest_val[14]));
 sky130_fd_sc_hd__a41o_1 _11143_ (.A1(_03861_),
    .A2(_03950_),
    .A3(_04074_),
    .A4(_04181_),
    .B1(net155),
    .X(_04219_));
 sky130_fd_sc_hd__a21o_1 _11144_ (.A1(_04157_),
    .A2(_04166_),
    .B1(_04164_),
    .X(_04220_));
 sky130_fd_sc_hd__a21oi_1 _11145_ (.A1(_04133_),
    .A2(_04135_),
    .B1(_04131_),
    .Y(_04221_));
 sky130_fd_sc_hd__or2_1 _11146_ (.A(net113),
    .B(net31),
    .X(_04222_));
 sky130_fd_sc_hd__nor2_1 _11147_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__xnor2_1 _11148_ (.A(_04221_),
    .B(_04222_),
    .Y(_04224_));
 sky130_fd_sc_hd__nor2_1 _11149_ (.A(_04122_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__and2_1 _11150_ (.A(_04122_),
    .B(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__nor2_1 _11151_ (.A(_04225_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__o22a_1 _11152_ (.A1(net84),
    .A2(net15),
    .B1(net36),
    .B2(net79),
    .X(_04228_));
 sky130_fd_sc_hd__xnor2_1 _11153_ (.A(net76),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__o22a_1 _11154_ (.A1(net119),
    .A2(net9),
    .B1(net4),
    .B2(net123),
    .X(_04230_));
 sky130_fd_sc_hd__xnor2_1 _11155_ (.A(net34),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__o22a_1 _11156_ (.A1(net29),
    .A2(net41),
    .B1(net38),
    .B2(net27),
    .X(_04232_));
 sky130_fd_sc_hd__xnor2_1 _11157_ (.A(net111),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__xor2_1 _11158_ (.A(_04231_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__and2b_1 _11159_ (.A_N(_04229_),
    .B(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__xnor2_1 _11160_ (.A(_04229_),
    .B(_04234_),
    .Y(_04236_));
 sky130_fd_sc_hd__o22a_1 _11161_ (.A1(net21),
    .A2(net56),
    .B1(net17),
    .B2(net65),
    .X(_04237_));
 sky130_fd_sc_hd__xnor2_1 _11162_ (.A(net92),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__and2_1 _11163_ (.A(net149),
    .B(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__xnor2_1 _11164_ (.A(_06499_),
    .B(_04238_),
    .Y(_04240_));
 sky130_fd_sc_hd__o22a_1 _11165_ (.A1(net68),
    .A2(net12),
    .B1(net8),
    .B2(net94),
    .X(_04241_));
 sky130_fd_sc_hd__xnor2_1 _11166_ (.A(net100),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__and2_1 _11167_ (.A(_04240_),
    .B(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__nor2_1 _11168_ (.A(_04240_),
    .B(_04242_),
    .Y(_04244_));
 sky130_fd_sc_hd__nor2_1 _11169_ (.A(_04243_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__a21o_1 _11170_ (.A1(_00137_),
    .A2(_00138_),
    .B1(net48),
    .X(_04246_));
 sky130_fd_sc_hd__or2_1 _11171_ (.A(net70),
    .B(net44),
    .X(_04247_));
 sky130_fd_sc_hd__nand3_1 _11172_ (.A(net108),
    .B(_04246_),
    .C(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21o_1 _11173_ (.A1(_04246_),
    .A2(_04247_),
    .B1(net108),
    .X(_04249_));
 sky130_fd_sc_hd__o32a_1 _11174_ (.A1(_00176_),
    .A2(_00177_),
    .A3(net61),
    .B1(net58),
    .B2(net66),
    .X(_04250_));
 sky130_fd_sc_hd__xor2_1 _11175_ (.A(net102),
    .B(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__a21oi_1 _11176_ (.A1(_04248_),
    .A2(_04249_),
    .B1(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand3_1 _11177_ (.A(_04248_),
    .B(_04249_),
    .C(_04251_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand2b_1 _11178_ (.A_N(_04252_),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__o22a_1 _11179_ (.A1(net25),
    .A2(net53),
    .B1(net50),
    .B2(net72),
    .X(_04255_));
 sky130_fd_sc_hd__xnor2_1 _11180_ (.A(net105),
    .B(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__xnor2_1 _11181_ (.A(_04254_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__and2_1 _11182_ (.A(_04116_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__or2_1 _11183_ (.A(_04116_),
    .B(_04257_),
    .X(_04259_));
 sky130_fd_sc_hd__nand2b_1 _11184_ (.A_N(_04258_),
    .B(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__inv_2 _11185_ (.A(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__nand2_1 _11186_ (.A(_04245_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__or2_1 _11187_ (.A(_04245_),
    .B(_04261_),
    .X(_04263_));
 sky130_fd_sc_hd__and3_1 _11188_ (.A(_04236_),
    .B(_04262_),
    .C(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__a21o_1 _11189_ (.A1(_04262_),
    .A2(_04263_),
    .B1(_04236_),
    .X(_04265_));
 sky130_fd_sc_hd__nand2b_1 _11190_ (.A_N(_04264_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__xnor2_1 _11191_ (.A(_04227_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a21oi_1 _11192_ (.A1(_04150_),
    .A2(_04155_),
    .B1(_04148_),
    .Y(_04268_));
 sky130_fd_sc_hd__a21o_1 _11193_ (.A1(_04151_),
    .A2(_04153_),
    .B1(_04152_),
    .X(_04269_));
 sky130_fd_sc_hd__a21o_1 _11194_ (.A1(_04141_),
    .A2(_04146_),
    .B1(_04145_),
    .X(_04270_));
 sky130_fd_sc_hd__o21ai_1 _11195_ (.A1(_04124_),
    .A2(_04137_),
    .B1(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__or3_1 _11196_ (.A(_04124_),
    .B(_04137_),
    .C(_04270_),
    .X(_04272_));
 sky130_fd_sc_hd__and2_1 _11197_ (.A(_04271_),
    .B(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__xnor2_1 _11198_ (.A(_04269_),
    .B(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__a21bo_1 _11199_ (.A1(_04158_),
    .A2(_04162_),
    .B1_N(_04161_),
    .X(_04275_));
 sky130_fd_sc_hd__nand2b_1 _11200_ (.A_N(_04274_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__xnor2_1 _11201_ (.A(_04274_),
    .B(_04275_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2b_1 _11202_ (.A_N(_04268_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__xnor2_1 _11203_ (.A(_04268_),
    .B(_04277_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _11204_ (.A(_04267_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__xnor2_1 _11205_ (.A(_04267_),
    .B(_04279_),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2b_1 _11206_ (.A_N(_04281_),
    .B(_04220_),
    .Y(_04282_));
 sky130_fd_sc_hd__xor2_1 _11207_ (.A(_04220_),
    .B(_04281_),
    .X(_04283_));
 sky130_fd_sc_hd__a21oi_1 _11208_ (.A1(_04168_),
    .A2(_04171_),
    .B1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__a21o_1 _11209_ (.A1(_04168_),
    .A2(_04171_),
    .B1(_04283_),
    .X(_04285_));
 sky130_fd_sc_hd__and3_1 _11210_ (.A(_04168_),
    .B(_04171_),
    .C(_04283_),
    .X(_04286_));
 sky130_fd_sc_hd__nor2_2 _11211_ (.A(_04284_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__a21boi_1 _11212_ (.A1(_04064_),
    .A2(_04173_),
    .B1_N(_04174_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2b_1 _11213_ (.A_N(_04066_),
    .B(_04175_),
    .Y(_04289_));
 sky130_fd_sc_hd__a41o_1 _11214_ (.A1(_04064_),
    .A2(_04065_),
    .A3(_04067_),
    .A4(_04175_),
    .B1(_04288_),
    .X(_04290_));
 sky130_fd_sc_hd__or2_1 _11215_ (.A(_04068_),
    .B(_04289_),
    .X(_04291_));
 sky130_fd_sc_hd__o21ba_1 _11216_ (.A1(_03823_),
    .A2(_04291_),
    .B1_N(_04290_),
    .X(_04292_));
 sky130_fd_sc_hd__xor2_4 _11217_ (.A(_04287_),
    .B(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__nand2_1 _11218_ (.A(_04219_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__o21a_1 _11219_ (.A1(_04219_),
    .A2(_04293_),
    .B1(_02171_),
    .X(_04295_));
 sky130_fd_sc_hd__a21oi_1 _11220_ (.A1(_02107_),
    .A2(_02108_),
    .B1(net155),
    .Y(_04296_));
 sky130_fd_sc_hd__xnor2_1 _11221_ (.A(_02112_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a21o_1 _11222_ (.A1(_05943_),
    .A2(_04186_),
    .B1(_05925_),
    .X(_04298_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(_06366_),
    .A1(_04298_),
    .S(net303),
    .X(_04299_));
 sky130_fd_sc_hd__nand2_1 _11224_ (.A(_05889_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__o211a_1 _11225_ (.A1(_05889_),
    .A2(_04299_),
    .B1(_04300_),
    .C1(_02247_),
    .X(_04301_));
 sky130_fd_sc_hd__nor2_1 _11226_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _11227_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .Y(_04303_));
 sky130_fd_sc_hd__and2b_1 _11228_ (.A_N(_04302_),
    .B(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__o21a_1 _11229_ (.A1(_04192_),
    .A2(_04193_),
    .B1(_04191_),
    .X(_04305_));
 sky130_fd_sc_hd__xnor2_1 _11230_ (.A(_04304_),
    .B(_04305_),
    .Y(_04306_));
 sky130_fd_sc_hd__mux2_1 _11231_ (.A0(_03332_),
    .A1(_03334_),
    .S(net237),
    .X(_04307_));
 sky130_fd_sc_hd__inv_2 _11232_ (.A(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__mux2_2 _11233_ (.A0(_02270_),
    .A1(_04308_),
    .S(net239),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _11234_ (.A(net243),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__o211a_1 _11235_ (.A1(net243),
    .A2(_04306_),
    .B1(_04310_),
    .C1(net216),
    .X(_04311_));
 sky130_fd_sc_hd__or2_1 _11236_ (.A(\div_res[14] ),
    .B(_04204_),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(\div_res[15] ),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__a21o_1 _11238_ (.A1(net162),
    .A2(_04312_),
    .B1(\div_res[15] ),
    .X(_04314_));
 sky130_fd_sc_hd__o211a_1 _11239_ (.A1(_02071_),
    .A2(_04313_),
    .B1(_04314_),
    .C1(_02260_),
    .X(_04315_));
 sky130_fd_sc_hd__or2_1 _11240_ (.A(\div_shifter[46] ),
    .B(_04200_),
    .X(_04316_));
 sky130_fd_sc_hd__a21oi_1 _11241_ (.A1(net248),
    .A2(_04316_),
    .B1(\div_shifter[47] ),
    .Y(_04317_));
 sky130_fd_sc_hd__a31o_1 _11242_ (.A1(\div_shifter[47] ),
    .A2(net249),
    .A3(_04316_),
    .B1(net251),
    .X(_04318_));
 sky130_fd_sc_hd__nor2_2 _11243_ (.A(_04317_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(net253),
    .A1(net206),
    .S(_05872_),
    .X(_04320_));
 sky130_fd_sc_hd__a21oi_1 _11245_ (.A1(net207),
    .A2(_04320_),
    .B1(_05880_),
    .Y(_04321_));
 sky130_fd_sc_hd__a211o_1 _11246_ (.A1(_05854_),
    .A2(_06459_),
    .B1(_04319_),
    .C1(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__o21a_1 _11247_ (.A1(net240),
    .A2(_02237_),
    .B1(_02272_),
    .X(_04323_));
 sky130_fd_sc_hd__a2bb2o_1 _11248_ (.A1_N(net188),
    .A2_N(_04309_),
    .B1(_04323_),
    .B2(net192),
    .X(_04324_));
 sky130_fd_sc_hd__or3_1 _11249_ (.A(_04315_),
    .B(_04322_),
    .C(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__or3_2 _11250_ (.A(_04301_),
    .B(_04311_),
    .C(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__a221o_1 _11251_ (.A1(_04294_),
    .A2(_04295_),
    .B1(_04297_),
    .B2(net252),
    .C1(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__or2_1 _11252_ (.A(curr_PC[15]),
    .B(_04216_),
    .X(_04328_));
 sky130_fd_sc_hd__and2_1 _11253_ (.A(curr_PC[15]),
    .B(_04216_),
    .X(_04329_));
 sky130_fd_sc_hd__nor2_1 _11254_ (.A(net263),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__a22o_4 _11255_ (.A1(net263),
    .A2(_04327_),
    .B1(_04328_),
    .B2(_04330_),
    .X(dest_val[15]));
 sky130_fd_sc_hd__and3b_1 _11256_ (.A_N(_04110_),
    .B(_04181_),
    .C(_04293_),
    .X(_04331_));
 sky130_fd_sc_hd__a21o_1 _11257_ (.A1(_04253_),
    .A2(_04256_),
    .B1(_04252_),
    .X(_04332_));
 sky130_fd_sc_hd__o22a_1 _11258_ (.A1(net73),
    .A2(net61),
    .B1(net50),
    .B2(net26),
    .X(_04333_));
 sky130_fd_sc_hd__xor2_1 _11259_ (.A(net106),
    .B(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__o22a_1 _11260_ (.A1(net22),
    .A2(net58),
    .B1(net56),
    .B2(net67),
    .X(_04335_));
 sky130_fd_sc_hd__xor2_1 _11261_ (.A(net102),
    .B(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__nor2_1 _11262_ (.A(_04334_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__and2_1 _11263_ (.A(_04334_),
    .B(_04336_),
    .X(_04338_));
 sky130_fd_sc_hd__nor2_1 _11264_ (.A(_04337_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(_04332_),
    .B(_04339_),
    .Y(_04341_));
 sky130_fd_sc_hd__or2_1 _11266_ (.A(_04332_),
    .B(_04339_),
    .X(_04342_));
 sky130_fd_sc_hd__nand2_1 _11267_ (.A(_04341_),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__o22a_1 _11268_ (.A1(net20),
    .A2(net17),
    .B1(net12),
    .B2(net64),
    .X(_04344_));
 sky130_fd_sc_hd__xnor2_1 _11269_ (.A(net91),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__o31a_1 _11270_ (.A1(_06499_),
    .A2(_00159_),
    .A3(net6),
    .B1(net100),
    .X(_04346_));
 sky130_fd_sc_hd__nor2_1 _11271_ (.A(_00161_),
    .B(net8),
    .Y(_04347_));
 sky130_fd_sc_hd__nor3_2 _11272_ (.A(_04345_),
    .B(_04346_),
    .C(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__o21a_1 _11273_ (.A1(_04346_),
    .A2(_04347_),
    .B1(_04345_),
    .X(_04349_));
 sky130_fd_sc_hd__nor2_1 _11274_ (.A(_04348_),
    .B(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_1 _11275_ (.A(_04343_),
    .B(_04350_),
    .Y(_04352_));
 sky130_fd_sc_hd__o22a_1 _11276_ (.A1(net80),
    .A2(net15),
    .B1(net36),
    .B2(net41),
    .X(_04353_));
 sky130_fd_sc_hd__xnor2_1 _11277_ (.A(net76),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__o22a_1 _11278_ (.A1(net71),
    .A2(net53),
    .B1(net44),
    .B2(net24),
    .X(_04355_));
 sky130_fd_sc_hd__xnor2_1 _11279_ (.A(net109),
    .B(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__and2b_1 _11280_ (.A_N(_04354_),
    .B(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__and2b_1 _11281_ (.A_N(_04356_),
    .B(_04354_),
    .X(_04358_));
 sky130_fd_sc_hd__or2_1 _11282_ (.A(_04357_),
    .B(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__o22a_1 _11283_ (.A1(net27),
    .A2(net47),
    .B1(net38),
    .B2(net29),
    .X(_04360_));
 sky130_fd_sc_hd__xnor2_1 _11284_ (.A(net111),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__and2b_1 _11285_ (.A_N(_04359_),
    .B(_04361_),
    .X(_04363_));
 sky130_fd_sc_hd__and2b_1 _11286_ (.A_N(_04361_),
    .B(_04359_),
    .X(_04364_));
 sky130_fd_sc_hd__or2_1 _11287_ (.A(_04363_),
    .B(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__xnor2_1 _11288_ (.A(_04352_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__o22a_1 _11289_ (.A1(net85),
    .A2(net9),
    .B1(net4),
    .B2(net119),
    .X(_04367_));
 sky130_fd_sc_hd__xnor2_1 _11290_ (.A(net34),
    .B(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__o21a_1 _11291_ (.A1(_04239_),
    .A2(_04243_),
    .B1(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__nor3_1 _11292_ (.A(_04239_),
    .B(_04243_),
    .C(_04368_),
    .Y(_04370_));
 sky130_fd_sc_hd__nor2_1 _11293_ (.A(_04369_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__or2_1 _11294_ (.A(net123),
    .B(net31),
    .X(_04372_));
 sky130_fd_sc_hd__xnor2_1 _11295_ (.A(_04371_),
    .B(_04372_),
    .Y(_04374_));
 sky130_fd_sc_hd__and2b_1 _11296_ (.A_N(_04366_),
    .B(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__xnor2_1 _11297_ (.A(_04366_),
    .B(_04374_),
    .Y(_04376_));
 sky130_fd_sc_hd__a21oi_1 _11298_ (.A1(_04227_),
    .A2(_04265_),
    .B1(_04264_),
    .Y(_04377_));
 sky130_fd_sc_hd__a21o_1 _11299_ (.A1(_04231_),
    .A2(_04233_),
    .B1(_04235_),
    .X(_04378_));
 sky130_fd_sc_hd__a21o_1 _11300_ (.A1(_04245_),
    .A2(_04259_),
    .B1(_04258_),
    .X(_04379_));
 sky130_fd_sc_hd__xor2_1 _11301_ (.A(_04378_),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__o21ai_1 _11302_ (.A1(_04223_),
    .A2(_04225_),
    .B1(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__or3_1 _11303_ (.A(_04223_),
    .B(_04225_),
    .C(_04380_),
    .X(_04382_));
 sky130_fd_sc_hd__nand2_1 _11304_ (.A(_04381_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21bo_1 _11305_ (.A1(_04269_),
    .A2(_04272_),
    .B1_N(_04271_),
    .X(_04385_));
 sky130_fd_sc_hd__xnor2_1 _11306_ (.A(_04383_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__and2b_1 _11307_ (.A_N(_04377_),
    .B(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__xnor2_1 _11308_ (.A(_04377_),
    .B(_04386_),
    .Y(_04388_));
 sky130_fd_sc_hd__nand2_1 _11309_ (.A(_04376_),
    .B(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__xnor2_1 _11310_ (.A(_04376_),
    .B(_04388_),
    .Y(_04390_));
 sky130_fd_sc_hd__and2_1 _11311_ (.A(_04276_),
    .B(_04278_),
    .X(_04391_));
 sky130_fd_sc_hd__or2_1 _11312_ (.A(_04390_),
    .B(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__xnor2_1 _11313_ (.A(_04390_),
    .B(_04391_),
    .Y(_04393_));
 sky130_fd_sc_hd__a21o_1 _11314_ (.A1(_04280_),
    .A2(_04282_),
    .B1(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__nand3_1 _11315_ (.A(_04280_),
    .B(_04282_),
    .C(_04393_),
    .Y(_04396_));
 sky130_fd_sc_hd__and2_2 _11316_ (.A(_04394_),
    .B(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__a21oi_1 _11317_ (.A1(_04173_),
    .A2(_04285_),
    .B1(_04286_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _11318_ (.A(_04175_),
    .B(_04287_),
    .Y(_04399_));
 sky130_fd_sc_hd__nor2_1 _11319_ (.A(_04176_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__nor2_1 _11320_ (.A(_04177_),
    .B(_04399_),
    .Y(_04401_));
 sky130_fd_sc_hd__a211o_1 _11321_ (.A1(_03946_),
    .A2(_04401_),
    .B1(_04400_),
    .C1(_04398_),
    .X(_04402_));
 sky130_fd_sc_hd__a31o_4 _11322_ (.A1(_03453_),
    .A2(_03940_),
    .A3(_04401_),
    .B1(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__xnor2_4 _11323_ (.A(_04397_),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__o21ai_1 _11324_ (.A1(net155),
    .A2(_04331_),
    .B1(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__or3_1 _11325_ (.A(net155),
    .B(_04331_),
    .C(_04404_),
    .X(_04407_));
 sky130_fd_sc_hd__and3_1 _11326_ (.A(_02171_),
    .B(_04405_),
    .C(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__o21ai_1 _11327_ (.A1(net155),
    .A2(_02113_),
    .B1(_02114_),
    .Y(_04409_));
 sky130_fd_sc_hd__or3_1 _11328_ (.A(net155),
    .B(_02113_),
    .C(_02114_),
    .X(_04410_));
 sky130_fd_sc_hd__a21o_1 _11329_ (.A1(_05889_),
    .A2(_04298_),
    .B1(_05872_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(_06367_),
    .A1(_04411_),
    .S(net303),
    .X(_04412_));
 sky130_fd_sc_hd__or2_1 _11331_ (.A(_05835_),
    .B(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__nand2_1 _11332_ (.A(_05835_),
    .B(_04412_),
    .Y(_04414_));
 sky130_fd_sc_hd__o21a_1 _11333_ (.A1(_04302_),
    .A2(_04305_),
    .B1(_04303_),
    .X(_04415_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04416_));
 sky130_fd_sc_hd__nand2_1 _11335_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04418_));
 sky130_fd_sc_hd__and2b_1 _11336_ (.A_N(_04416_),
    .B(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__xnor2_1 _11337_ (.A(_04415_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(_04323_),
    .A1(_04420_),
    .S(net268),
    .X(_04421_));
 sky130_fd_sc_hd__or2_1 _11339_ (.A(\div_shifter[47] ),
    .B(_04316_),
    .X(_04422_));
 sky130_fd_sc_hd__a21o_1 _11340_ (.A1(net248),
    .A2(_04422_),
    .B1(\div_shifter[48] ),
    .X(_04423_));
 sky130_fd_sc_hd__nand3_1 _11341_ (.A(\div_shifter[48] ),
    .B(net248),
    .C(_04422_),
    .Y(_04424_));
 sky130_fd_sc_hd__o21ai_1 _11342_ (.A1(_05817_),
    .A2(net253),
    .B1(net207),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_1 _11343_ (.A(_05799_),
    .B(net215),
    .Y(_04426_));
 sky130_fd_sc_hd__a221o_2 _11344_ (.A1(_05817_),
    .A2(_02255_),
    .B1(_04425_),
    .B2(_05826_),
    .C1(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__a31o_2 _11345_ (.A1(_02258_),
    .A2(_04423_),
    .A3(_04424_),
    .B1(_04427_),
    .X(_04429_));
 sky130_fd_sc_hd__or2_1 _11346_ (.A(\div_res[15] ),
    .B(_04312_),
    .X(_04430_));
 sky130_fd_sc_hd__a21oi_1 _11347_ (.A1(net162),
    .A2(_04430_),
    .B1(\div_res[16] ),
    .Y(_04431_));
 sky130_fd_sc_hd__a31o_1 _11348_ (.A1(\div_res[16] ),
    .A2(net162),
    .A3(_04430_),
    .B1(net204),
    .X(_04432_));
 sky130_fd_sc_hd__o2bb2a_1 _11349_ (.A1_N(_02243_),
    .A2_N(_04323_),
    .B1(_04431_),
    .B2(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__o21ai_1 _11350_ (.A1(net190),
    .A2(_04309_),
    .B1(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__a211o_1 _11351_ (.A1(net216),
    .A2(_04421_),
    .B1(_04429_),
    .C1(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__a31o_1 _11352_ (.A1(_02247_),
    .A2(_04413_),
    .A3(_04414_),
    .B1(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__a311o_1 _11353_ (.A1(net252),
    .A2(_04409_),
    .A3(_04410_),
    .B1(_04436_),
    .C1(_04408_),
    .X(_04437_));
 sky130_fd_sc_hd__nand2_1 _11354_ (.A(curr_PC[16]),
    .B(_04329_),
    .Y(_04438_));
 sky130_fd_sc_hd__o21a_1 _11355_ (.A1(curr_PC[16]),
    .A2(_04329_),
    .B1(net267),
    .X(_04440_));
 sky130_fd_sc_hd__a22o_4 _11356_ (.A1(net263),
    .A2(_04437_),
    .B1(_04438_),
    .B2(_04440_),
    .X(dest_val[16]));
 sky130_fd_sc_hd__and3_1 _11357_ (.A(curr_PC[16]),
    .B(curr_PC[17]),
    .C(_04329_),
    .X(_04441_));
 sky130_fd_sc_hd__a21oi_1 _11358_ (.A1(curr_PC[16]),
    .A2(_04329_),
    .B1(curr_PC[17]),
    .Y(_04442_));
 sky130_fd_sc_hd__o21ai_1 _11359_ (.A1(_04441_),
    .A2(_04442_),
    .B1(net267),
    .Y(_04443_));
 sky130_fd_sc_hd__nand2_1 _11360_ (.A(_04331_),
    .B(_04404_),
    .Y(_04444_));
 sky130_fd_sc_hd__nand2_1 _11361_ (.A(net159),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__a31o_1 _11362_ (.A1(_04381_),
    .A2(_04382_),
    .A3(_04385_),
    .B1(_04387_),
    .X(_04446_));
 sky130_fd_sc_hd__o22a_1 _11363_ (.A1(net79),
    .A2(net9),
    .B1(net4),
    .B2(net84),
    .X(_04447_));
 sky130_fd_sc_hd__xnor2_2 _11364_ (.A(net34),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__o22a_1 _11365_ (.A1(net41),
    .A2(net15),
    .B1(net36),
    .B2(net38),
    .X(_04450_));
 sky130_fd_sc_hd__xnor2_1 _11366_ (.A(net76),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__or2_1 _11367_ (.A(net120),
    .B(net31),
    .X(_04452_));
 sky130_fd_sc_hd__nor2_1 _11368_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__and2_1 _11369_ (.A(_04451_),
    .B(_04452_),
    .X(_04454_));
 sky130_fd_sc_hd__nor2_1 _11370_ (.A(_04453_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__xnor2_2 _11371_ (.A(_04448_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__o22a_1 _11372_ (.A1(net29),
    .A2(net47),
    .B1(net44),
    .B2(net27),
    .X(_04457_));
 sky130_fd_sc_hd__xnor2_1 _11373_ (.A(net111),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__o22a_1 _11374_ (.A1(net26),
    .A2(net61),
    .B1(net58),
    .B2(net73),
    .X(_04459_));
 sky130_fd_sc_hd__xnor2_1 _11375_ (.A(net106),
    .B(_04459_),
    .Y(_04461_));
 sky130_fd_sc_hd__and2_1 _11376_ (.A(_04458_),
    .B(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__nor2_1 _11377_ (.A(_04458_),
    .B(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__nor2_1 _11378_ (.A(_04462_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__o22a_1 _11379_ (.A1(net24),
    .A2(net53),
    .B1(net50),
    .B2(net71),
    .X(_04465_));
 sky130_fd_sc_hd__xnor2_1 _11380_ (.A(net109),
    .B(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__xor2_1 _11381_ (.A(_04464_),
    .B(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__o22a_1 _11382_ (.A1(net22),
    .A2(net56),
    .B1(net17),
    .B2(net67),
    .X(_04468_));
 sky130_fd_sc_hd__xnor2_1 _11383_ (.A(net104),
    .B(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__and2_1 _11384_ (.A(_00153_),
    .B(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__xnor2_1 _11385_ (.A(net101),
    .B(_04469_),
    .Y(_04472_));
 sky130_fd_sc_hd__o22a_1 _11386_ (.A1(net21),
    .A2(net12),
    .B1(net8),
    .B2(net65),
    .X(_04473_));
 sky130_fd_sc_hd__xnor2_1 _11387_ (.A(net92),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__and2_1 _11388_ (.A(_04472_),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__nor2_1 _11389_ (.A(_04472_),
    .B(_04474_),
    .Y(_04476_));
 sky130_fd_sc_hd__or2_1 _11390_ (.A(_04475_),
    .B(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__nor2_1 _11391_ (.A(_04348_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__nand2_1 _11392_ (.A(_04348_),
    .B(_04477_),
    .Y(_04479_));
 sky130_fd_sc_hd__and2b_1 _11393_ (.A_N(_04478_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__xor2_1 _11394_ (.A(_04337_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__and2_1 _11395_ (.A(_04467_),
    .B(_04481_),
    .X(_04483_));
 sky130_fd_sc_hd__nor2_1 _11396_ (.A(_04467_),
    .B(_04481_),
    .Y(_04484_));
 sky130_fd_sc_hd__nor2_1 _11397_ (.A(_04483_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__xnor2_2 _11398_ (.A(_04456_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__o21ba_1 _11399_ (.A1(_04352_),
    .A2(_04365_),
    .B1_N(_04375_),
    .X(_04487_));
 sky130_fd_sc_hd__o21bai_2 _11400_ (.A1(_04370_),
    .A2(_04372_),
    .B1_N(_04369_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21ai_2 _11401_ (.A1(_04343_),
    .A2(_04350_),
    .B1(_04341_),
    .Y(_04489_));
 sky130_fd_sc_hd__nor2_1 _11402_ (.A(_04357_),
    .B(_04363_),
    .Y(_04490_));
 sky130_fd_sc_hd__o21ai_1 _11403_ (.A1(_04357_),
    .A2(_04363_),
    .B1(_04489_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_2 _11404_ (.A(_04489_),
    .B(_04490_),
    .Y(_04492_));
 sky130_fd_sc_hd__xnor2_2 _11405_ (.A(_04488_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__a21bo_1 _11406_ (.A1(_04378_),
    .A2(_04379_),
    .B1_N(_04381_),
    .X(_04494_));
 sky130_fd_sc_hd__nand2b_1 _11407_ (.A_N(_04493_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__xnor2_2 _11408_ (.A(_04493_),
    .B(_04494_),
    .Y(_04496_));
 sky130_fd_sc_hd__nand2b_1 _11409_ (.A_N(_04487_),
    .B(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__xnor2_2 _11410_ (.A(_04487_),
    .B(_04496_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _11411_ (.A(_04486_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__xor2_2 _11412_ (.A(_04486_),
    .B(_04498_),
    .X(_04500_));
 sky130_fd_sc_hd__nand2_1 _11413_ (.A(_04446_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__xnor2_2 _11414_ (.A(_04446_),
    .B(_04500_),
    .Y(_04502_));
 sky130_fd_sc_hd__a21oi_2 _11415_ (.A1(_04389_),
    .A2(_04392_),
    .B1(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__a21o_1 _11416_ (.A1(_04389_),
    .A2(_04392_),
    .B1(_04502_),
    .X(_04504_));
 sky130_fd_sc_hd__and3_1 _11417_ (.A(_04389_),
    .B(_04392_),
    .C(_04502_),
    .X(_04505_));
 sky130_fd_sc_hd__or2_2 _11418_ (.A(_04503_),
    .B(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__a21boi_1 _11419_ (.A1(_04285_),
    .A2(_04394_),
    .B1_N(_04396_),
    .Y(_04507_));
 sky130_fd_sc_hd__inv_2 _11420_ (.A(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__nand2_1 _11421_ (.A(_04287_),
    .B(_04397_),
    .Y(_04509_));
 sky130_fd_sc_hd__a31o_1 _11422_ (.A1(_04287_),
    .A2(_04288_),
    .A3(_04397_),
    .B1(_04507_),
    .X(_04510_));
 sky130_fd_sc_hd__or2_1 _11423_ (.A(_04289_),
    .B(_04509_),
    .X(_04511_));
 sky130_fd_sc_hd__nor2_1 _11424_ (.A(_04069_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__a311o_1 _11425_ (.A1(_03577_),
    .A2(_03579_),
    .A3(_03580_),
    .B1(_04070_),
    .C1(_04511_),
    .X(_04514_));
 sky130_fd_sc_hd__or3b_4 _11426_ (.A(_04510_),
    .B(_04512_),
    .C_N(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__xor2_4 _11427_ (.A(_04506_),
    .B(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__inv_2 _11428_ (.A(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__a31o_1 _11429_ (.A1(net159),
    .A2(_04444_),
    .A3(_04517_),
    .B1(net209),
    .X(_04518_));
 sky130_fd_sc_hd__a21oi_1 _11430_ (.A1(_04445_),
    .A2(_04516_),
    .B1(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__a21o_1 _11431_ (.A1(_02113_),
    .A2(_02114_),
    .B1(net155),
    .X(_04520_));
 sky130_fd_sc_hd__o21a_1 _11432_ (.A1(_02117_),
    .A2(_04520_),
    .B1(net252),
    .X(_04521_));
 sky130_fd_sc_hd__a21boi_1 _11433_ (.A1(_02117_),
    .A2(_04520_),
    .B1_N(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__a21o_1 _11434_ (.A1(_05826_),
    .A2(_04411_),
    .B1(_05817_),
    .X(_04523_));
 sky130_fd_sc_hd__inv_2 _11435_ (.A(_04523_),
    .Y(_04525_));
 sky130_fd_sc_hd__mux2_1 _11436_ (.A0(_06368_),
    .A1(_04525_),
    .S(net303),
    .X(_04526_));
 sky130_fd_sc_hd__xor2_1 _11437_ (.A(_05772_),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__o21a_1 _11438_ (.A1(_04415_),
    .A2(_04416_),
    .B1(_04418_),
    .X(_04528_));
 sky130_fd_sc_hd__nor2_1 _11439_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04529_));
 sky130_fd_sc_hd__nand2_1 _11440_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04530_));
 sky130_fd_sc_hd__nand2b_1 _11441_ (.A_N(_04529_),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__xor2_1 _11442_ (.A(_04528_),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__or2_1 _11443_ (.A(net268),
    .B(_04211_),
    .X(_04533_));
 sky130_fd_sc_hd__o211a_1 _11444_ (.A1(net244),
    .A2(_04532_),
    .B1(_04533_),
    .C1(net216),
    .X(_04534_));
 sky130_fd_sc_hd__o21ai_1 _11445_ (.A1(_05754_),
    .A2(net253),
    .B1(net207),
    .Y(_04536_));
 sky130_fd_sc_hd__o21ai_1 _11446_ (.A1(_05734_),
    .A2(net215),
    .B1(net266),
    .Y(_04537_));
 sky130_fd_sc_hd__a221o_1 _11447_ (.A1(_05754_),
    .A2(_02255_),
    .B1(_04536_),
    .B2(_05763_),
    .C1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__a21oi_1 _11448_ (.A1(_02243_),
    .A2(_04211_),
    .B1(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__or2_1 _11449_ (.A(\div_res[16] ),
    .B(_04430_),
    .X(_04540_));
 sky130_fd_sc_hd__and3_1 _11450_ (.A(\div_res[17] ),
    .B(net162),
    .C(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__a21oi_1 _11451_ (.A1(net162),
    .A2(_04540_),
    .B1(\div_res[17] ),
    .Y(_04542_));
 sky130_fd_sc_hd__o21a_1 _11452_ (.A1(\div_shifter[48] ),
    .A2(_04422_),
    .B1(net249),
    .X(_04543_));
 sky130_fd_sc_hd__o21ai_1 _11453_ (.A1(\div_shifter[49] ),
    .A2(_04543_),
    .B1(_02258_),
    .Y(_04544_));
 sky130_fd_sc_hd__a21o_1 _11454_ (.A1(\div_shifter[49] ),
    .A2(_04543_),
    .B1(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__o31a_1 _11455_ (.A1(net204),
    .A2(_04541_),
    .A3(_04542_),
    .B1(_04545_),
    .X(_04547_));
 sky130_fd_sc_hd__o211ai_1 _11456_ (.A1(net190),
    .A2(_04197_),
    .B1(_04539_),
    .C1(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__a211o_1 _11457_ (.A1(_02247_),
    .A2(_04527_),
    .B1(_04534_),
    .C1(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__o31a_4 _11458_ (.A1(_04519_),
    .A2(_04522_),
    .A3(_04549_),
    .B1(_04443_),
    .X(dest_val[17]));
 sky130_fd_sc_hd__a31o_1 _11459_ (.A1(_04331_),
    .A2(_04404_),
    .A3(_04516_),
    .B1(net156),
    .X(_04550_));
 sky130_fd_sc_hd__o22a_1 _11460_ (.A1(net71),
    .A2(net61),
    .B1(net50),
    .B2(net24),
    .X(_04551_));
 sky130_fd_sc_hd__xnor2_1 _11461_ (.A(net109),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__o22a_1 _11462_ (.A1(net22),
    .A2(net17),
    .B1(net12),
    .B2(net67),
    .X(_04553_));
 sky130_fd_sc_hd__xnor2_1 _11463_ (.A(net104),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__and2_1 _11464_ (.A(_04552_),
    .B(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__nor2_1 _11465_ (.A(_04552_),
    .B(_04554_),
    .Y(_04557_));
 sky130_fd_sc_hd__nor2_1 _11466_ (.A(_04555_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__o22a_1 _11467_ (.A1(net26),
    .A2(net58),
    .B1(net56),
    .B2(net73),
    .X(_04559_));
 sky130_fd_sc_hd__xnor2_1 _11468_ (.A(net106),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__xor2_1 _11469_ (.A(_04558_),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__or3_1 _11470_ (.A(net100),
    .B(_00187_),
    .C(net6),
    .X(_04562_));
 sky130_fd_sc_hd__a2bb2o_4 _11471_ (.A1_N(_00188_),
    .A2_N(net6),
    .B1(_04562_),
    .B2(net91),
    .X(_04563_));
 sky130_fd_sc_hd__nor2_1 _11472_ (.A(net84),
    .B(net31),
    .Y(_04564_));
 sky130_fd_sc_hd__xnor2_1 _11473_ (.A(_04563_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__o21ai_1 _11474_ (.A1(_04470_),
    .A2(_04475_),
    .B1(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__or3_1 _11475_ (.A(_04470_),
    .B(_04475_),
    .C(_04565_),
    .X(_04568_));
 sky130_fd_sc_hd__and2_1 _11476_ (.A(_04566_),
    .B(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__nand2_1 _11477_ (.A(_04561_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__or2_1 _11478_ (.A(_04561_),
    .B(_04569_),
    .X(_04571_));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_04570_),
    .B(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__o22a_1 _11480_ (.A1(net38),
    .A2(net15),
    .B1(net36),
    .B2(net47),
    .X(_04573_));
 sky130_fd_sc_hd__xnor2_1 _11481_ (.A(net76),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__o22a_1 _11482_ (.A1(net41),
    .A2(net9),
    .B1(net4),
    .B2(net79),
    .X(_04575_));
 sky130_fd_sc_hd__xnor2_1 _11483_ (.A(net34),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__o22a_1 _11484_ (.A1(net27),
    .A2(net53),
    .B1(net44),
    .B2(net29),
    .X(_04577_));
 sky130_fd_sc_hd__xnor2_1 _11485_ (.A(net111),
    .B(_04577_),
    .Y(_04579_));
 sky130_fd_sc_hd__xor2_1 _11486_ (.A(_04576_),
    .B(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__and2b_1 _11487_ (.A_N(_04574_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__xor2_1 _11488_ (.A(_04574_),
    .B(_04580_),
    .X(_04582_));
 sky130_fd_sc_hd__xor2_1 _11489_ (.A(_04572_),
    .B(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__o21ba_1 _11490_ (.A1(_04456_),
    .A2(_04484_),
    .B1_N(_04483_),
    .X(_04584_));
 sky130_fd_sc_hd__a21bo_1 _11491_ (.A1(_04488_),
    .A2(_04492_),
    .B1_N(_04491_),
    .X(_04585_));
 sky130_fd_sc_hd__a21o_1 _11492_ (.A1(_04448_),
    .A2(_04455_),
    .B1(_04453_),
    .X(_04586_));
 sky130_fd_sc_hd__a21o_1 _11493_ (.A1(_04464_),
    .A2(_04466_),
    .B1(_04462_),
    .X(_04587_));
 sky130_fd_sc_hd__a21o_1 _11494_ (.A1(_04337_),
    .A2(_04479_),
    .B1(_04478_),
    .X(_04588_));
 sky130_fd_sc_hd__xor2_1 _11495_ (.A(_04587_),
    .B(_04588_),
    .X(_04590_));
 sky130_fd_sc_hd__nand2_1 _11496_ (.A(_04586_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__xnor2_1 _11497_ (.A(_04586_),
    .B(_04590_),
    .Y(_04592_));
 sky130_fd_sc_hd__and2b_1 _11498_ (.A_N(_04592_),
    .B(_04585_),
    .X(_04593_));
 sky130_fd_sc_hd__xnor2_1 _11499_ (.A(_04585_),
    .B(_04592_),
    .Y(_04594_));
 sky130_fd_sc_hd__and2b_1 _11500_ (.A_N(_04584_),
    .B(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__xnor2_1 _11501_ (.A(_04584_),
    .B(_04594_),
    .Y(_04596_));
 sky130_fd_sc_hd__and2_1 _11502_ (.A(_04583_),
    .B(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__xnor2_1 _11503_ (.A(_04583_),
    .B(_04596_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _11504_ (.A(_04495_),
    .B(_04497_),
    .Y(_04599_));
 sky130_fd_sc_hd__and2b_1 _11505_ (.A_N(_04598_),
    .B(_04599_),
    .X(_04601_));
 sky130_fd_sc_hd__xor2_1 _11506_ (.A(_04598_),
    .B(_04599_),
    .X(_04602_));
 sky130_fd_sc_hd__a21oi_2 _11507_ (.A1(_04499_),
    .A2(_04501_),
    .B1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand3_2 _11508_ (.A(_04499_),
    .B(_04501_),
    .C(_04602_),
    .Y(_04604_));
 sky130_fd_sc_hd__nand2b_2 _11509_ (.A_N(_04603_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__a21o_1 _11510_ (.A1(_04394_),
    .A2(_04504_),
    .B1(_04505_),
    .X(_04606_));
 sky130_fd_sc_hd__or3b_2 _11511_ (.A(_04503_),
    .B(_04505_),
    .C_N(_04397_),
    .X(_04607_));
 sky130_fd_sc_hd__inv_2 _11512_ (.A(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__a21bo_1 _11513_ (.A1(_04398_),
    .A2(_04608_),
    .B1_N(_04606_),
    .X(_04609_));
 sky130_fd_sc_hd__nor2_1 _11514_ (.A(_04399_),
    .B(_04607_),
    .Y(_04610_));
 sky130_fd_sc_hd__and2_1 _11515_ (.A(_04178_),
    .B(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__a311o_4 _11516_ (.A1(_03702_),
    .A2(_04179_),
    .A3(_04610_),
    .B1(_04612_),
    .C1(_04609_),
    .X(_04613_));
 sky130_fd_sc_hd__xor2_4 _11517_ (.A(_04605_),
    .B(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__inv_2 _11518_ (.A(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _11519_ (.A(_04550_),
    .B(_04614_),
    .Y(_04616_));
 sky130_fd_sc_hd__a21o_1 _11520_ (.A1(_04550_),
    .A2(_04614_),
    .B1(net209),
    .X(_04617_));
 sky130_fd_sc_hd__or3_1 _11521_ (.A(net155),
    .B(_02118_),
    .C(_02119_),
    .X(_04618_));
 sky130_fd_sc_hd__o21ai_1 _11522_ (.A1(net155),
    .A2(_02118_),
    .B1(_02119_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_04618_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__or2_1 _11524_ (.A(net303),
    .B(_06369_),
    .X(_04621_));
 sky130_fd_sc_hd__a21o_1 _11525_ (.A1(_05763_),
    .A2(_04523_),
    .B1(_05754_),
    .X(_04623_));
 sky130_fd_sc_hd__nand2_1 _11526_ (.A(net303),
    .B(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__a21oi_1 _11527_ (.A1(_04621_),
    .A2(_04624_),
    .B1(_05706_),
    .Y(_04625_));
 sky130_fd_sc_hd__a31o_1 _11528_ (.A1(_05706_),
    .A2(_04621_),
    .A3(_04624_),
    .B1(net255),
    .X(_04626_));
 sky130_fd_sc_hd__or2_1 _11529_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .X(_04627_));
 sky130_fd_sc_hd__nand2_1 _11530_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04628_));
 sky130_fd_sc_hd__o21ai_1 _11531_ (.A1(_04528_),
    .A2(_04529_),
    .B1(_04530_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand3_1 _11532_ (.A(_04627_),
    .B(_04628_),
    .C(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21o_1 _11533_ (.A1(_04627_),
    .A2(_04628_),
    .B1(_04629_),
    .X(_04631_));
 sky130_fd_sc_hd__a21oi_1 _11534_ (.A1(_04630_),
    .A2(_04631_),
    .B1(net243),
    .Y(_04632_));
 sky130_fd_sc_hd__a211o_1 _11535_ (.A1(net244),
    .A2(_04102_),
    .B1(_04632_),
    .C1(_06447_),
    .X(_04634_));
 sky130_fd_sc_hd__or3_1 _11536_ (.A(\div_shifter[49] ),
    .B(\div_shifter[48] ),
    .C(_04422_),
    .X(_04635_));
 sky130_fd_sc_hd__a21oi_1 _11537_ (.A1(net248),
    .A2(_04635_),
    .B1(\div_shifter[50] ),
    .Y(_04636_));
 sky130_fd_sc_hd__a31o_1 _11538_ (.A1(\div_shifter[50] ),
    .A2(net248),
    .A3(_04635_),
    .B1(net250),
    .X(_04637_));
 sky130_fd_sc_hd__or2_2 _11539_ (.A(_04636_),
    .B(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__nand2_1 _11540_ (.A(_05677_),
    .B(_02255_),
    .Y(_04639_));
 sky130_fd_sc_hd__o211a_1 _11541_ (.A1(_05677_),
    .A2(net253),
    .B1(_04639_),
    .C1(net207),
    .X(_04640_));
 sky130_fd_sc_hd__o22a_1 _11542_ (.A1(_05649_),
    .A2(net215),
    .B1(_04640_),
    .B2(_05687_),
    .X(_04641_));
 sky130_fd_sc_hd__o221a_1 _11543_ (.A1(net190),
    .A2(_04089_),
    .B1(_04102_),
    .B2(net188),
    .C1(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__or2_1 _11544_ (.A(\div_res[17] ),
    .B(_04540_),
    .X(_04643_));
 sky130_fd_sc_hd__a21oi_1 _11545_ (.A1(net162),
    .A2(_04643_),
    .B1(\div_res[18] ),
    .Y(_04645_));
 sky130_fd_sc_hd__a31o_1 _11546_ (.A1(\div_res[18] ),
    .A2(net162),
    .A3(_04643_),
    .B1(net204),
    .X(_04646_));
 sky130_fd_sc_hd__o211a_1 _11547_ (.A1(_04645_),
    .A2(_04646_),
    .B1(_04638_),
    .C1(_04642_),
    .X(_04647_));
 sky130_fd_sc_hd__o211a_1 _11548_ (.A1(_04625_),
    .A2(_04626_),
    .B1(_04634_),
    .C1(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__o221a_1 _11549_ (.A1(_04616_),
    .A2(_04617_),
    .B1(_04620_),
    .B2(_02254_),
    .C1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__and2_2 _11550_ (.A(curr_PC[18]),
    .B(_04441_),
    .X(_04650_));
 sky130_fd_sc_hd__o21ai_1 _11551_ (.A1(curr_PC[18]),
    .A2(_04441_),
    .B1(net267),
    .Y(_04651_));
 sky130_fd_sc_hd__o22ai_4 _11552_ (.A1(net267),
    .A2(_04649_),
    .B1(_04650_),
    .B2(_04651_),
    .Y(dest_val[18]));
 sky130_fd_sc_hd__o31a_1 _11553_ (.A1(_04444_),
    .A2(_04517_),
    .A3(_04615_),
    .B1(net159),
    .X(_04652_));
 sky130_fd_sc_hd__o22a_1 _11554_ (.A1(net38),
    .A2(net9),
    .B1(net4),
    .B2(net41),
    .X(_04653_));
 sky130_fd_sc_hd__xnor2_1 _11555_ (.A(net34),
    .B(_04653_),
    .Y(_04655_));
 sky130_fd_sc_hd__nand2_1 _11556_ (.A(_04563_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__xnor2_1 _11557_ (.A(_04563_),
    .B(_04655_),
    .Y(_04657_));
 sky130_fd_sc_hd__or3_1 _11558_ (.A(net79),
    .B(net31),
    .C(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__o21ai_1 _11559_ (.A1(net79),
    .A2(net31),
    .B1(_04657_),
    .Y(_04659_));
 sky130_fd_sc_hd__and2_1 _11560_ (.A(_04658_),
    .B(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__inv_2 _11561_ (.A(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__o22a_1 _11562_ (.A1(net26),
    .A2(net56),
    .B1(net17),
    .B2(net73),
    .X(_04662_));
 sky130_fd_sc_hd__xor2_1 _11563_ (.A(net106),
    .B(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__xnor2_1 _11564_ (.A(net92),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__o22a_1 _11565_ (.A1(net22),
    .A2(net12),
    .B1(net8),
    .B2(net67),
    .X(_04666_));
 sky130_fd_sc_hd__xor2_1 _11566_ (.A(net104),
    .B(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__or2_1 _11567_ (.A(_04664_),
    .B(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__nand2_1 _11568_ (.A(_04664_),
    .B(_04667_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_1 _11569_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__xor2_1 _11570_ (.A(_04660_),
    .B(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__o22a_1 _11571_ (.A1(net47),
    .A2(net15),
    .B1(net36),
    .B2(net44),
    .X(_04672_));
 sky130_fd_sc_hd__xnor2_1 _11572_ (.A(net76),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__o22a_1 _11573_ (.A1(net24),
    .A2(net61),
    .B1(net58),
    .B2(net71),
    .X(_04674_));
 sky130_fd_sc_hd__xor2_1 _11574_ (.A(net109),
    .B(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__xnor2_1 _11575_ (.A(_04673_),
    .B(_04675_),
    .Y(_04677_));
 sky130_fd_sc_hd__o22a_1 _11576_ (.A1(net29),
    .A2(net53),
    .B1(net50),
    .B2(net27),
    .X(_04678_));
 sky130_fd_sc_hd__xnor2_1 _11577_ (.A(net111),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__and2b_1 _11578_ (.A_N(_04677_),
    .B(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__and2b_1 _11579_ (.A_N(_04679_),
    .B(_04677_),
    .X(_04681_));
 sky130_fd_sc_hd__or2_1 _11580_ (.A(_04680_),
    .B(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__or2_1 _11581_ (.A(_04671_),
    .B(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__nand2_1 _11582_ (.A(_04671_),
    .B(_04682_),
    .Y(_04684_));
 sky130_fd_sc_hd__and2_1 _11583_ (.A(_04683_),
    .B(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__o21ai_1 _11584_ (.A1(_04572_),
    .A2(_04582_),
    .B1(_04570_),
    .Y(_04686_));
 sky130_fd_sc_hd__a21o_1 _11585_ (.A1(_04576_),
    .A2(_04579_),
    .B1(_04581_),
    .X(_04688_));
 sky130_fd_sc_hd__a21o_1 _11586_ (.A1(_04558_),
    .A2(_04560_),
    .B1(_04555_),
    .X(_04689_));
 sky130_fd_sc_hd__o31ai_2 _11587_ (.A1(net84),
    .A2(net31),
    .A3(_04563_),
    .B1(_04566_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_04689_),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__xor2_1 _11589_ (.A(_04689_),
    .B(_04690_),
    .X(_04692_));
 sky130_fd_sc_hd__nand2_1 _11590_ (.A(_04688_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__xnor2_1 _11591_ (.A(_04688_),
    .B(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__a21boi_1 _11592_ (.A1(_04587_),
    .A2(_04588_),
    .B1_N(_04591_),
    .Y(_04695_));
 sky130_fd_sc_hd__or2_1 _11593_ (.A(_04694_),
    .B(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__xnor2_1 _11594_ (.A(_04694_),
    .B(_04695_),
    .Y(_04697_));
 sky130_fd_sc_hd__nand2b_1 _11595_ (.A_N(_04697_),
    .B(_04686_),
    .Y(_04699_));
 sky130_fd_sc_hd__xnor2_1 _11596_ (.A(_04686_),
    .B(_04697_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand2_1 _11597_ (.A(_04685_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__xor2_1 _11598_ (.A(_04685_),
    .B(_04700_),
    .X(_04702_));
 sky130_fd_sc_hd__nor2_1 _11599_ (.A(_04593_),
    .B(_04595_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand2b_1 _11600_ (.A_N(_04703_),
    .B(_04702_),
    .Y(_04704_));
 sky130_fd_sc_hd__xnor2_1 _11601_ (.A(_04702_),
    .B(_04703_),
    .Y(_04705_));
 sky130_fd_sc_hd__o21a_1 _11602_ (.A1(_04597_),
    .A2(_04601_),
    .B1(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__nor3_1 _11603_ (.A(_04597_),
    .B(_04601_),
    .C(_04705_),
    .Y(_04707_));
 sky130_fd_sc_hd__nor2_1 _11604_ (.A(_04706_),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__o21ai_2 _11605_ (.A1(_04503_),
    .A2(_04603_),
    .B1(_04604_),
    .Y(_04710_));
 sky130_fd_sc_hd__or2_2 _11606_ (.A(_04506_),
    .B(_04605_),
    .X(_04711_));
 sky130_fd_sc_hd__o21ai_1 _11607_ (.A1(_04508_),
    .A2(_04711_),
    .B1(_04710_),
    .Y(_04712_));
 sky130_fd_sc_hd__nor2_1 _11608_ (.A(_04509_),
    .B(_04711_),
    .Y(_04713_));
 sky130_fd_sc_hd__inv_2 _11609_ (.A(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__a21oi_1 _11610_ (.A1(_04290_),
    .A2(_04713_),
    .B1(_04712_),
    .Y(_04715_));
 sky130_fd_sc_hd__o31a_2 _11611_ (.A1(_03823_),
    .A2(_04291_),
    .A3(_04714_),
    .B1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__xnor2_1 _11612_ (.A(_04708_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__xor2_1 _11613_ (.A(_04708_),
    .B(_04716_),
    .X(_04718_));
 sky130_fd_sc_hd__or2_1 _11614_ (.A(_04652_),
    .B(_04717_),
    .X(_04719_));
 sky130_fd_sc_hd__a21oi_1 _11615_ (.A1(_04652_),
    .A2(_04717_),
    .B1(net209),
    .Y(_04721_));
 sky130_fd_sc_hd__and3_1 _11616_ (.A(net159),
    .B(_02120_),
    .C(_02123_),
    .X(_04722_));
 sky130_fd_sc_hd__a21oi_1 _11617_ (.A1(net159),
    .A2(_02120_),
    .B1(_02123_),
    .Y(_04723_));
 sky130_fd_sc_hd__nor2_1 _11618_ (.A(_04722_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__or2_1 _11619_ (.A(net303),
    .B(_06370_),
    .X(_04725_));
 sky130_fd_sc_hd__a21oi_1 _11620_ (.A1(_05696_),
    .A2(_04623_),
    .B1(_05677_),
    .Y(_04726_));
 sky130_fd_sc_hd__or2_1 _11621_ (.A(net309),
    .B(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__a21oi_1 _11622_ (.A1(_04725_),
    .A2(_04727_),
    .B1(_05620_),
    .Y(_04728_));
 sky130_fd_sc_hd__and3_1 _11623_ (.A(_05620_),
    .B(_04725_),
    .C(_04727_),
    .X(_04729_));
 sky130_fd_sc_hd__or3_1 _11624_ (.A(net255),
    .B(_04728_),
    .C(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__or2_1 _11625_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .X(_04732_));
 sky130_fd_sc_hd__nand2_1 _11626_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04733_));
 sky130_fd_sc_hd__nand2_1 _11627_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__a21bo_1 _11628_ (.A1(_04627_),
    .A2(_04629_),
    .B1_N(_04628_),
    .X(_04735_));
 sky130_fd_sc_hd__xnor2_1 _11629_ (.A(_04734_),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__or2_1 _11630_ (.A(net268),
    .B(_03979_),
    .X(_04737_));
 sky130_fd_sc_hd__o211a_1 _11631_ (.A1(net244),
    .A2(_04736_),
    .B1(_04737_),
    .C1(net216),
    .X(_04738_));
 sky130_fd_sc_hd__or2_1 _11632_ (.A(\div_res[18] ),
    .B(_04643_),
    .X(_04739_));
 sky130_fd_sc_hd__and3_1 _11633_ (.A(\div_res[19] ),
    .B(net163),
    .C(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__a21oi_1 _11634_ (.A1(net163),
    .A2(_04739_),
    .B1(\div_res[19] ),
    .Y(_04741_));
 sky130_fd_sc_hd__or2_1 _11635_ (.A(\div_shifter[50] ),
    .B(_04635_),
    .X(_04743_));
 sky130_fd_sc_hd__and3_1 _11636_ (.A(\div_shifter[51] ),
    .B(net246),
    .C(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__a21oi_1 _11637_ (.A1(net246),
    .A2(_04743_),
    .B1(\div_shifter[51] ),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(_05588_),
    .B(_02255_),
    .Y(_04746_));
 sky130_fd_sc_hd__o211a_1 _11639_ (.A1(_05588_),
    .A2(net253),
    .B1(_04746_),
    .C1(net207),
    .X(_04747_));
 sky130_fd_sc_hd__o22a_1 _11640_ (.A1(_05567_),
    .A2(net215),
    .B1(_04747_),
    .B2(_05599_),
    .X(_04748_));
 sky130_fd_sc_hd__o221a_1 _11641_ (.A1(net190),
    .A2(_03961_),
    .B1(_03980_),
    .B2(net188),
    .C1(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__o31a_1 _11642_ (.A1(net251),
    .A2(_04744_),
    .A3(_04745_),
    .B1(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__o31ai_1 _11643_ (.A1(net204),
    .A2(_04740_),
    .A3(_04741_),
    .B1(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__or3b_2 _11644_ (.A(_04751_),
    .B(_04738_),
    .C_N(_04730_),
    .X(_04752_));
 sky130_fd_sc_hd__a221o_1 _11645_ (.A1(_04719_),
    .A2(_04721_),
    .B1(_04724_),
    .B2(net252),
    .C1(_04752_),
    .X(_04754_));
 sky130_fd_sc_hd__or2_1 _11646_ (.A(curr_PC[19]),
    .B(_04650_),
    .X(_04755_));
 sky130_fd_sc_hd__a21oi_1 _11647_ (.A1(curr_PC[19]),
    .A2(_04650_),
    .B1(net263),
    .Y(_04756_));
 sky130_fd_sc_hd__a22o_4 _11648_ (.A1(net263),
    .A2(_04754_),
    .B1(_04755_),
    .B2(_04756_),
    .X(dest_val[19]));
 sky130_fd_sc_hd__and4_1 _11649_ (.A(_04404_),
    .B(_04516_),
    .C(_04614_),
    .D(_04718_),
    .X(_04757_));
 sky130_fd_sc_hd__nand4b_4 _11650_ (.A_N(_04110_),
    .B(_04181_),
    .C(_04293_),
    .D(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__o22a_1 _11651_ (.A1(net26),
    .A2(net17),
    .B1(net12),
    .B2(net73),
    .X(_04759_));
 sky130_fd_sc_hd__xnor2_1 _11652_ (.A(net106),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nor2_1 _11653_ (.A(net22),
    .B(net8),
    .Y(_04761_));
 sky130_fd_sc_hd__xnor2_1 _11654_ (.A(net104),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__and2b_1 _11655_ (.A_N(_04760_),
    .B(_04762_),
    .X(_04764_));
 sky130_fd_sc_hd__inv_2 _11656_ (.A(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__and2b_1 _11657_ (.A_N(_04762_),
    .B(_04760_),
    .X(_04766_));
 sky130_fd_sc_hd__nor2_1 _11658_ (.A(_04764_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__o22a_1 _11659_ (.A1(net47),
    .A2(net9),
    .B1(net4),
    .B2(net38),
    .X(_04768_));
 sky130_fd_sc_hd__nand2_1 _11660_ (.A(net41),
    .B(net34),
    .Y(_04769_));
 sky130_fd_sc_hd__xnor2_1 _11661_ (.A(_04768_),
    .B(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__or2_1 _11662_ (.A(_04767_),
    .B(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_04767_),
    .B(_04770_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand2_1 _11664_ (.A(_04771_),
    .B(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__o22a_1 _11665_ (.A1(net44),
    .A2(net15),
    .B1(net36),
    .B2(net53),
    .X(_04775_));
 sky130_fd_sc_hd__xnor2_1 _11666_ (.A(net76),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__o22a_1 _11667_ (.A1(net24),
    .A2(net58),
    .B1(net56),
    .B2(net71),
    .X(_04777_));
 sky130_fd_sc_hd__xor2_1 _11668_ (.A(net109),
    .B(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__nor2_1 _11669_ (.A(_04776_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__and2_1 _11670_ (.A(_04776_),
    .B(_04778_),
    .X(_04780_));
 sky130_fd_sc_hd__or2_1 _11671_ (.A(_04779_),
    .B(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__o22a_1 _11672_ (.A1(net27),
    .A2(net61),
    .B1(net50),
    .B2(net29),
    .X(_04782_));
 sky130_fd_sc_hd__xnor2_1 _11673_ (.A(_06524_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__nor2_1 _11674_ (.A(_04781_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__and2_1 _11675_ (.A(_04781_),
    .B(_04783_),
    .X(_04786_));
 sky130_fd_sc_hd__or2_1 _11676_ (.A(_04784_),
    .B(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__xor2_1 _11677_ (.A(_04773_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__o21a_1 _11678_ (.A1(_04661_),
    .A2(_04670_),
    .B1(_04683_),
    .X(_04789_));
 sky130_fd_sc_hd__o21bai_2 _11679_ (.A1(_04673_),
    .A2(_04675_),
    .B1_N(_04680_),
    .Y(_04790_));
 sky130_fd_sc_hd__o21a_1 _11680_ (.A1(net92),
    .A2(_04663_),
    .B1(_04668_),
    .X(_04791_));
 sky130_fd_sc_hd__a21oi_1 _11681_ (.A1(_04656_),
    .A2(_04658_),
    .B1(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__and3_1 _11682_ (.A(_04656_),
    .B(_04658_),
    .C(_04791_),
    .X(_04793_));
 sky130_fd_sc_hd__nor2_1 _11683_ (.A(_04792_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__and2_1 _11684_ (.A(_04790_),
    .B(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__xnor2_1 _11685_ (.A(_04790_),
    .B(_04794_),
    .Y(_04797_));
 sky130_fd_sc_hd__a21o_1 _11686_ (.A1(_04691_),
    .A2(_04693_),
    .B1(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__nand3_1 _11687_ (.A(_04691_),
    .B(_04693_),
    .C(_04797_),
    .Y(_04799_));
 sky130_fd_sc_hd__nand2_1 _11688_ (.A(_04798_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__xor2_1 _11689_ (.A(_04789_),
    .B(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__nand2_1 _11690_ (.A(_04788_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__xnor2_1 _11691_ (.A(_04788_),
    .B(_04801_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21o_1 _11692_ (.A1(_04696_),
    .A2(_04699_),
    .B1(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__nand3_1 _11693_ (.A(_04696_),
    .B(_04699_),
    .C(_04803_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand2_1 _11694_ (.A(_04804_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__a21o_1 _11695_ (.A1(_04701_),
    .A2(_04704_),
    .B1(_04806_),
    .X(_04808_));
 sky130_fd_sc_hd__inv_2 _11696_ (.A(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__nand3_1 _11697_ (.A(_04701_),
    .B(_04704_),
    .C(_04806_),
    .Y(_04810_));
 sky130_fd_sc_hd__and2_1 _11698_ (.A(_04808_),
    .B(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__o21bai_1 _11699_ (.A1(_04603_),
    .A2(_04706_),
    .B1_N(_04707_),
    .Y(_04812_));
 sky130_fd_sc_hd__or3_1 _11700_ (.A(_04605_),
    .B(_04706_),
    .C(_04707_),
    .X(_04813_));
 sky130_fd_sc_hd__o21ai_1 _11701_ (.A1(_04606_),
    .A2(_04813_),
    .B1(_04812_),
    .Y(_04814_));
 sky130_fd_sc_hd__nor2_2 _11702_ (.A(_04607_),
    .B(_04813_),
    .Y(_04815_));
 sky130_fd_sc_hd__a21oi_2 _11703_ (.A1(_04403_),
    .A2(_04815_),
    .B1(_04814_),
    .Y(_04816_));
 sky130_fd_sc_hd__xnor2_2 _11704_ (.A(_04811_),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__and3_1 _11705_ (.A(net159),
    .B(_04758_),
    .C(_04817_),
    .X(_04819_));
 sky130_fd_sc_hd__a21o_1 _11706_ (.A1(net159),
    .A2(_04758_),
    .B1(_04817_),
    .X(_04820_));
 sky130_fd_sc_hd__nand2_1 _11707_ (.A(_02171_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__o21a_1 _11708_ (.A1(_02120_),
    .A2(_02123_),
    .B1(net159),
    .X(_04822_));
 sky130_fd_sc_hd__xor2_1 _11709_ (.A(_02124_),
    .B(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__o21bai_1 _11710_ (.A1(_05620_),
    .A2(_04726_),
    .B1_N(_05588_),
    .Y(_04824_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(_06371_),
    .A1(_04824_),
    .S(net303),
    .X(_04825_));
 sky130_fd_sc_hd__o21ai_1 _11712_ (.A1(_05459_),
    .A2(_04825_),
    .B1(_02247_),
    .Y(_04826_));
 sky130_fd_sc_hd__a21o_1 _11713_ (.A1(_05459_),
    .A2(_04825_),
    .B1(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__or2_1 _11714_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_1 _11715_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .Y(_04830_));
 sky130_fd_sc_hd__nand2_1 _11716_ (.A(_04828_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__a21boi_1 _11717_ (.A1(_04732_),
    .A2(_04735_),
    .B1_N(_04733_),
    .Y(_04832_));
 sky130_fd_sc_hd__xnor2_1 _11718_ (.A(_04831_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(_03854_),
    .A1(_04833_),
    .S(net268),
    .X(_04834_));
 sky130_fd_sc_hd__or2_1 _11720_ (.A(\div_res[19] ),
    .B(_04739_),
    .X(_04835_));
 sky130_fd_sc_hd__a21oi_1 _11721_ (.A1(net162),
    .A2(_04835_),
    .B1(\div_res[20] ),
    .Y(_04836_));
 sky130_fd_sc_hd__a31o_1 _11722_ (.A1(\div_res[20] ),
    .A2(net162),
    .A3(_04835_),
    .B1(net204),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _11723_ (.A(_04836_),
    .B(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__or2_1 _11724_ (.A(\div_shifter[51] ),
    .B(_04743_),
    .X(_04839_));
 sky130_fd_sc_hd__a21oi_1 _11725_ (.A1(net246),
    .A2(_04839_),
    .B1(\div_shifter[52] ),
    .Y(_04841_));
 sky130_fd_sc_hd__a31o_1 _11726_ (.A1(\div_shifter[52] ),
    .A2(net246),
    .A3(_04839_),
    .B1(net251),
    .X(_04842_));
 sky130_fd_sc_hd__nand2_1 _11727_ (.A(_05437_),
    .B(_02255_),
    .Y(_04843_));
 sky130_fd_sc_hd__o211a_1 _11728_ (.A1(_05437_),
    .A2(net253),
    .B1(_04843_),
    .C1(net207),
    .X(_04844_));
 sky130_fd_sc_hd__o22a_1 _11729_ (.A1(_05416_),
    .A2(net215),
    .B1(_04844_),
    .B2(_05448_),
    .X(_04845_));
 sky130_fd_sc_hd__o221a_1 _11730_ (.A1(net190),
    .A2(_03842_),
    .B1(_03854_),
    .B2(net188),
    .C1(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__o211a_1 _11731_ (.A1(_04841_),
    .A2(_04842_),
    .B1(_04846_),
    .C1(_04838_),
    .X(_04847_));
 sky130_fd_sc_hd__o211a_1 _11732_ (.A1(_06447_),
    .A2(_04834_),
    .B1(_04847_),
    .C1(_04827_),
    .X(_04848_));
 sky130_fd_sc_hd__o221a_1 _11733_ (.A1(_04819_),
    .A2(_04821_),
    .B1(_04823_),
    .B2(_02254_),
    .C1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__and3_1 _11734_ (.A(curr_PC[19]),
    .B(curr_PC[20]),
    .C(_04650_),
    .X(_04850_));
 sky130_fd_sc_hd__a21oi_1 _11735_ (.A1(curr_PC[19]),
    .A2(_04650_),
    .B1(curr_PC[20]),
    .Y(_04852_));
 sky130_fd_sc_hd__or3_1 _11736_ (.A(net263),
    .B(_04850_),
    .C(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__o21ai_4 _11737_ (.A1(net267),
    .A2(_04849_),
    .B1(_04853_),
    .Y(dest_val[20]));
 sky130_fd_sc_hd__o21a_1 _11738_ (.A1(_04758_),
    .A2(_04817_),
    .B1(net159),
    .X(_04854_));
 sky130_fd_sc_hd__o21ai_1 _11739_ (.A1(_04789_),
    .A2(_04800_),
    .B1(_04798_),
    .Y(_04855_));
 sky130_fd_sc_hd__o22a_1 _11740_ (.A1(net44),
    .A2(net9),
    .B1(net4),
    .B2(net47),
    .X(_04856_));
 sky130_fd_sc_hd__xnor2_1 _11741_ (.A(net34),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__o22a_1 _11742_ (.A1(net29),
    .A2(net61),
    .B1(net58),
    .B2(net27),
    .X(_04858_));
 sky130_fd_sc_hd__xnor2_1 _11743_ (.A(net111),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__nand2_1 _11744_ (.A(_04857_),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__or2_1 _11745_ (.A(_04857_),
    .B(_04859_),
    .X(_04862_));
 sky130_fd_sc_hd__and2_1 _11746_ (.A(_04860_),
    .B(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__inv_2 _11747_ (.A(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__o22a_1 _11748_ (.A1(net53),
    .A2(net15),
    .B1(net36),
    .B2(net50),
    .X(_04865_));
 sky130_fd_sc_hd__xnor2_1 _11749_ (.A(net76),
    .B(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__xor2_1 _11750_ (.A(_04863_),
    .B(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__or3b_1 _11751_ (.A(net41),
    .B(net31),
    .C_N(_04768_),
    .X(_04868_));
 sky130_fd_sc_hd__or2_1 _11752_ (.A(_04867_),
    .B(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__inv_2 _11753_ (.A(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__and2_1 _11754_ (.A(_04867_),
    .B(_04868_),
    .X(_04871_));
 sky130_fd_sc_hd__nor2_1 _11755_ (.A(_04870_),
    .B(_04871_),
    .Y(_04873_));
 sky130_fd_sc_hd__o22a_1 _11756_ (.A1(net24),
    .A2(net56),
    .B1(net17),
    .B2(net71),
    .X(_04874_));
 sky130_fd_sc_hd__xor2_2 _11757_ (.A(net109),
    .B(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__xnor2_1 _11758_ (.A(net104),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__o22a_1 _11759_ (.A1(net26),
    .A2(net12),
    .B1(net8),
    .B2(net73),
    .X(_04877_));
 sky130_fd_sc_hd__xnor2_1 _11760_ (.A(net106),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__and2b_1 _11761_ (.A_N(_04876_),
    .B(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__and2b_1 _11762_ (.A_N(_04878_),
    .B(_04876_),
    .X(_04880_));
 sky130_fd_sc_hd__or2_1 _11763_ (.A(_04879_),
    .B(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__xnor2_1 _11764_ (.A(_04873_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21a_1 _11765_ (.A1(_04773_),
    .A2(_04787_),
    .B1(_04771_),
    .X(_04884_));
 sky130_fd_sc_hd__or2_1 _11766_ (.A(net38),
    .B(net31),
    .X(_04885_));
 sky130_fd_sc_hd__o21ba_1 _11767_ (.A1(_04779_),
    .A2(_04784_),
    .B1_N(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__or3b_1 _11768_ (.A(_04779_),
    .B(_04784_),
    .C_N(_04885_),
    .X(_04887_));
 sky130_fd_sc_hd__and2b_1 _11769_ (.A_N(_04886_),
    .B(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__xnor2_1 _11770_ (.A(_04764_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__o21ai_1 _11771_ (.A1(_04792_),
    .A2(_04795_),
    .B1(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__or3_1 _11772_ (.A(_04792_),
    .B(_04795_),
    .C(_04889_),
    .X(_04891_));
 sky130_fd_sc_hd__and2_1 _11773_ (.A(_04890_),
    .B(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__nand2b_1 _11774_ (.A_N(_04884_),
    .B(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__xnor2_1 _11775_ (.A(_04884_),
    .B(_04892_),
    .Y(_04895_));
 sky130_fd_sc_hd__nand2_1 _11776_ (.A(_04882_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__xnor2_1 _11777_ (.A(_04882_),
    .B(_04895_),
    .Y(_04897_));
 sky130_fd_sc_hd__nand2b_1 _11778_ (.A_N(_04897_),
    .B(_04855_),
    .Y(_04898_));
 sky130_fd_sc_hd__xor2_1 _11779_ (.A(_04855_),
    .B(_04897_),
    .X(_04899_));
 sky130_fd_sc_hd__a21o_1 _11780_ (.A1(_04802_),
    .A2(_04804_),
    .B1(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__inv_2 _11781_ (.A(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__and3_1 _11782_ (.A(_04802_),
    .B(_04804_),
    .C(_04899_),
    .X(_04902_));
 sky130_fd_sc_hd__nor2_2 _11783_ (.A(_04901_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__o21ai_1 _11784_ (.A1(_04706_),
    .A2(_04809_),
    .B1(_04810_),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_04708_),
    .B(_04811_),
    .Y(_04906_));
 sky130_fd_sc_hd__o21ai_1 _11786_ (.A1(_04710_),
    .A2(_04906_),
    .B1(_04904_),
    .Y(_04907_));
 sky130_fd_sc_hd__nor2_1 _11787_ (.A(_04711_),
    .B(_04906_),
    .Y(_04908_));
 sky130_fd_sc_hd__a21oi_1 _11788_ (.A1(_04515_),
    .A2(_04908_),
    .B1(_04907_),
    .Y(_04909_));
 sky130_fd_sc_hd__xnor2_2 _11789_ (.A(_04903_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__nor2_1 _11790_ (.A(_04854_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__a21o_1 _11791_ (.A1(_04854_),
    .A2(_04910_),
    .B1(net209),
    .X(_04912_));
 sky130_fd_sc_hd__nor2_1 _11792_ (.A(net155),
    .B(_02125_),
    .Y(_04913_));
 sky130_fd_sc_hd__xnor2_1 _11793_ (.A(_02129_),
    .B(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__a21o_1 _11794_ (.A1(_05459_),
    .A2(_04824_),
    .B1(_05437_),
    .X(_04915_));
 sky130_fd_sc_hd__o21a_1 _11795_ (.A1(_05459_),
    .A2(_06371_),
    .B1(_06374_),
    .X(_04917_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(_04915_),
    .A1(_04917_),
    .S(net309),
    .X(_04918_));
 sky130_fd_sc_hd__xnor2_1 _11797_ (.A(_05524_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__or2_1 _11798_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .X(_04920_));
 sky130_fd_sc_hd__nand2_1 _11799_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_1 _11800_ (.A(_04920_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21ai_1 _11801_ (.A1(_04831_),
    .A2(_04832_),
    .B1(_04830_),
    .Y(_04923_));
 sky130_fd_sc_hd__xnor2_1 _11802_ (.A(_04922_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__nor2_1 _11803_ (.A(net243),
    .B(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__a211o_1 _11804_ (.A1(net243),
    .A2(_03732_),
    .B1(_04925_),
    .C1(_06447_),
    .X(_04926_));
 sky130_fd_sc_hd__or2_1 _11805_ (.A(\div_res[20] ),
    .B(_04835_),
    .X(_04928_));
 sky130_fd_sc_hd__a21oi_1 _11806_ (.A1(net162),
    .A2(_04928_),
    .B1(\div_res[21] ),
    .Y(_04929_));
 sky130_fd_sc_hd__a31o_1 _11807_ (.A1(\div_res[21] ),
    .A2(net162),
    .A3(_04928_),
    .B1(net204),
    .X(_04930_));
 sky130_fd_sc_hd__or2_1 _11808_ (.A(\div_shifter[52] ),
    .B(_04839_),
    .X(_04931_));
 sky130_fd_sc_hd__a21oi_1 _11809_ (.A1(net246),
    .A2(_04931_),
    .B1(\div_shifter[53] ),
    .Y(_04932_));
 sky130_fd_sc_hd__a311o_1 _11810_ (.A1(\div_shifter[53] ),
    .A2(net246),
    .A3(_04931_),
    .B1(_04932_),
    .C1(net251),
    .X(_04933_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(net253),
    .A1(net206),
    .S(_05502_),
    .X(_04934_));
 sky130_fd_sc_hd__a21o_1 _11812_ (.A1(net207),
    .A2(_04934_),
    .B1(_05513_),
    .X(_04935_));
 sky130_fd_sc_hd__o221a_1 _11813_ (.A1(_05491_),
    .A2(net215),
    .B1(net188),
    .B2(_03732_),
    .C1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__a21boi_1 _11814_ (.A1(net192),
    .A2(_03719_),
    .B1_N(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__o211a_1 _11815_ (.A1(_04929_),
    .A2(_04930_),
    .B1(_04933_),
    .C1(_04937_),
    .X(_04939_));
 sky130_fd_sc_hd__o211a_1 _11816_ (.A1(net255),
    .A2(_04919_),
    .B1(_04926_),
    .C1(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__o221a_1 _11817_ (.A1(_04911_),
    .A2(_04912_),
    .B1(_04914_),
    .B2(_02254_),
    .C1(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_1 _11818_ (.A(curr_PC[21]),
    .B(_04850_),
    .Y(_04942_));
 sky130_fd_sc_hd__and2_1 _11819_ (.A(curr_PC[21]),
    .B(_04850_),
    .X(_04943_));
 sky130_fd_sc_hd__or3_1 _11820_ (.A(net263),
    .B(_04942_),
    .C(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__o21ai_4 _11821_ (.A1(net267),
    .A2(_04941_),
    .B1(_04944_),
    .Y(dest_val[21]));
 sky130_fd_sc_hd__or2_1 _11822_ (.A(_04817_),
    .B(_04910_),
    .X(_04945_));
 sky130_fd_sc_hd__or2_1 _11823_ (.A(_04758_),
    .B(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__nand2_1 _11824_ (.A(_04890_),
    .B(_04893_),
    .Y(_04947_));
 sky130_fd_sc_hd__o21a_1 _11825_ (.A1(_04864_),
    .A2(_04866_),
    .B1(_04860_),
    .X(_04949_));
 sky130_fd_sc_hd__o22a_1 _11826_ (.A1(net50),
    .A2(net15),
    .B1(net36),
    .B2(net61),
    .X(_04950_));
 sky130_fd_sc_hd__xnor2_1 _11827_ (.A(net76),
    .B(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__o22a_1 _11828_ (.A1(net29),
    .A2(net58),
    .B1(net56),
    .B2(net27),
    .X(_04952_));
 sky130_fd_sc_hd__xnor2_1 _11829_ (.A(net111),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__and2b_1 _11830_ (.A_N(_04951_),
    .B(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__and2b_1 _11831_ (.A_N(_04953_),
    .B(_04951_),
    .X(_04955_));
 sky130_fd_sc_hd__or2_1 _11832_ (.A(_04954_),
    .B(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__xnor2_1 _11833_ (.A(_04949_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__o22a_1 _11834_ (.A1(net24),
    .A2(net17),
    .B1(net12),
    .B2(net71),
    .X(_04958_));
 sky130_fd_sc_hd__xnor2_1 _11835_ (.A(net109),
    .B(_04958_),
    .Y(_04960_));
 sky130_fd_sc_hd__o31a_1 _11836_ (.A1(net102),
    .A2(_06551_),
    .A3(net6),
    .B1(net105),
    .X(_04961_));
 sky130_fd_sc_hd__o21ba_2 _11837_ (.A1(_06552_),
    .A2(net6),
    .B1_N(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__and2b_1 _11838_ (.A_N(_04960_),
    .B(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__xnor2_1 _11839_ (.A(_04960_),
    .B(_04962_),
    .Y(_04964_));
 sky130_fd_sc_hd__xor2_1 _11840_ (.A(_04957_),
    .B(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__o21a_1 _11841_ (.A1(_04871_),
    .A2(_04881_),
    .B1(_04869_),
    .X(_04966_));
 sky130_fd_sc_hd__o21bai_2 _11842_ (.A1(net104),
    .A2(_04875_),
    .B1_N(_04879_),
    .Y(_04967_));
 sky130_fd_sc_hd__o22a_1 _11843_ (.A1(net53),
    .A2(net9),
    .B1(net4),
    .B2(net44),
    .X(_04968_));
 sky130_fd_sc_hd__xnor2_1 _11844_ (.A(net34),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand2_1 _11845_ (.A(_04967_),
    .B(_04969_),
    .Y(_04971_));
 sky130_fd_sc_hd__xnor2_1 _11846_ (.A(_04967_),
    .B(_04969_),
    .Y(_04972_));
 sky130_fd_sc_hd__or3_1 _11847_ (.A(net47),
    .B(net31),
    .C(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__o21ai_1 _11848_ (.A1(net47),
    .A2(net31),
    .B1(_04972_),
    .Y(_04974_));
 sky130_fd_sc_hd__and2_1 _11849_ (.A(_04973_),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__a21oi_1 _11850_ (.A1(_04765_),
    .A2(_04887_),
    .B1(_04886_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2b_1 _11851_ (.A_N(_04976_),
    .B(_04975_),
    .Y(_04977_));
 sky130_fd_sc_hd__and2b_1 _11852_ (.A_N(_04975_),
    .B(_04976_),
    .X(_04978_));
 sky130_fd_sc_hd__xnor2_1 _11853_ (.A(_04975_),
    .B(_04976_),
    .Y(_04979_));
 sky130_fd_sc_hd__xnor2_1 _11854_ (.A(_04966_),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _11855_ (.A(_04965_),
    .B(_04980_),
    .Y(_04982_));
 sky130_fd_sc_hd__or2_1 _11856_ (.A(_04965_),
    .B(_04980_),
    .X(_04983_));
 sky130_fd_sc_hd__nand2_1 _11857_ (.A(_04982_),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2b_1 _11858_ (.A_N(_04984_),
    .B(_04947_),
    .Y(_04985_));
 sky130_fd_sc_hd__xor2_1 _11859_ (.A(_04947_),
    .B(_04984_),
    .X(_04986_));
 sky130_fd_sc_hd__a21o_1 _11860_ (.A1(_04896_),
    .A2(_04898_),
    .B1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__and3_1 _11861_ (.A(_04896_),
    .B(_04898_),
    .C(_04986_),
    .X(_04988_));
 sky130_fd_sc_hd__inv_2 _11862_ (.A(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_2 _11863_ (.A(_04987_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__inv_2 _11864_ (.A(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__a21oi_1 _11865_ (.A1(_04808_),
    .A2(_04900_),
    .B1(_04902_),
    .Y(_04993_));
 sky130_fd_sc_hd__nand2_1 _11866_ (.A(_04811_),
    .B(_04903_),
    .Y(_04994_));
 sky130_fd_sc_hd__o21bai_1 _11867_ (.A1(_04812_),
    .A2(_04994_),
    .B1_N(_04993_),
    .Y(_04995_));
 sky130_fd_sc_hd__nor2_1 _11868_ (.A(_04813_),
    .B(_04994_),
    .Y(_04996_));
 sky130_fd_sc_hd__a21oi_2 _11869_ (.A1(_04613_),
    .A2(_04996_),
    .B1(_04995_),
    .Y(_04997_));
 sky130_fd_sc_hd__xnor2_2 _11870_ (.A(_04990_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__inv_2 _11871_ (.A(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__and3_1 _11872_ (.A(net159),
    .B(_04946_),
    .C(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__a21oi_1 _11873_ (.A1(net159),
    .A2(_04946_),
    .B1(_04999_),
    .Y(_05001_));
 sky130_fd_sc_hd__nand2_1 _11874_ (.A(net159),
    .B(_02130_),
    .Y(_05002_));
 sky130_fd_sc_hd__xnor2_1 _11875_ (.A(_02131_),
    .B(_05002_),
    .Y(_05004_));
 sky130_fd_sc_hd__nand2_1 _11876_ (.A(net252),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__a21o_1 _11877_ (.A1(_05524_),
    .A2(_04915_),
    .B1(_05502_),
    .X(_05006_));
 sky130_fd_sc_hd__o21a_1 _11878_ (.A1(_05524_),
    .A2(_04917_),
    .B1(_06373_),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_1 _11879_ (.A0(_05006_),
    .A1(_05007_),
    .S(net310),
    .X(_05008_));
 sky130_fd_sc_hd__xnor2_1 _11880_ (.A(_05383_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__or2_1 _11881_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .X(_05010_));
 sky130_fd_sc_hd__nand2_1 _11882_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _11883_ (.A(_05010_),
    .B(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__a21bo_1 _11884_ (.A1(_04920_),
    .A2(_04923_),
    .B1_N(_04921_),
    .X(_05013_));
 sky130_fd_sc_hd__xnor2_1 _11885_ (.A(_05012_),
    .B(_05013_),
    .Y(_05015_));
 sky130_fd_sc_hd__nor2_1 _11886_ (.A(net243),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__a211o_1 _11887_ (.A1(net243),
    .A2(_03610_),
    .B1(_05016_),
    .C1(_06447_),
    .X(_05017_));
 sky130_fd_sc_hd__or2_1 _11888_ (.A(\div_shifter[53] ),
    .B(_04931_),
    .X(_05018_));
 sky130_fd_sc_hd__a21oi_1 _11889_ (.A1(net246),
    .A2(_05018_),
    .B1(\div_shifter[54] ),
    .Y(_05019_));
 sky130_fd_sc_hd__a311o_1 _11890_ (.A1(\div_shifter[54] ),
    .A2(net246),
    .A3(_05018_),
    .B1(_05019_),
    .C1(net251),
    .X(_05020_));
 sky130_fd_sc_hd__or2_1 _11891_ (.A(\div_res[21] ),
    .B(_04928_),
    .X(_05021_));
 sky130_fd_sc_hd__a21oi_1 _11892_ (.A1(net162),
    .A2(_05021_),
    .B1(\div_res[22] ),
    .Y(_05022_));
 sky130_fd_sc_hd__a31o_1 _11893_ (.A1(\div_res[22] ),
    .A2(net162),
    .A3(_05021_),
    .B1(net204),
    .X(_05023_));
 sky130_fd_sc_hd__nand2_1 _11894_ (.A(_05361_),
    .B(_02255_),
    .Y(_05024_));
 sky130_fd_sc_hd__o211a_1 _11895_ (.A1(_05361_),
    .A2(net253),
    .B1(_05024_),
    .C1(net207),
    .X(_05026_));
 sky130_fd_sc_hd__o22a_1 _11896_ (.A1(_05340_),
    .A2(net215),
    .B1(_05026_),
    .B2(_05372_),
    .X(_05027_));
 sky130_fd_sc_hd__o221a_1 _11897_ (.A1(net190),
    .A2(_03598_),
    .B1(_03610_),
    .B2(net188),
    .C1(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__o211a_1 _11898_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_05028_),
    .C1(_05020_),
    .X(_05029_));
 sky130_fd_sc_hd__o211a_1 _11899_ (.A1(net255),
    .A2(_05009_),
    .B1(_05017_),
    .C1(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__o311a_1 _11900_ (.A1(net209),
    .A2(_05000_),
    .A3(_05001_),
    .B1(_05005_),
    .C1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__a21oi_1 _11901_ (.A1(curr_PC[22]),
    .A2(_04943_),
    .B1(net263),
    .Y(_05032_));
 sky130_fd_sc_hd__o21ai_2 _11902_ (.A1(curr_PC[22]),
    .A2(_04943_),
    .B1(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__o21ai_4 _11903_ (.A1(net267),
    .A2(_05031_),
    .B1(_05033_),
    .Y(dest_val[22]));
 sky130_fd_sc_hd__o21a_1 _11904_ (.A1(_04946_),
    .A2(_04999_),
    .B1(net159),
    .X(_05034_));
 sky130_fd_sc_hd__o22a_1 _11905_ (.A1(net29),
    .A2(net56),
    .B1(net17),
    .B2(net27),
    .X(_05036_));
 sky130_fd_sc_hd__xnor2_1 _11906_ (.A(net111),
    .B(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__and2b_1 _11907_ (.A_N(net106),
    .B(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__xnor2_1 _11908_ (.A(net106),
    .B(_05037_),
    .Y(_05039_));
 sky130_fd_sc_hd__o22a_1 _11909_ (.A1(net24),
    .A2(net12),
    .B1(net8),
    .B2(net71),
    .X(_05040_));
 sky130_fd_sc_hd__xnor2_1 _11910_ (.A(net109),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__and2_1 _11911_ (.A(_05039_),
    .B(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__nor2_1 _11912_ (.A(_05039_),
    .B(_05041_),
    .Y(_05043_));
 sky130_fd_sc_hd__or2_1 _11913_ (.A(_05042_),
    .B(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__or2_1 _11914_ (.A(_04963_),
    .B(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__nand2_1 _11915_ (.A(_04963_),
    .B(_05044_),
    .Y(_05047_));
 sky130_fd_sc_hd__and2_1 _11916_ (.A(_05045_),
    .B(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_04954_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__or2_1 _11918_ (.A(_04954_),
    .B(_05048_),
    .X(_05050_));
 sky130_fd_sc_hd__and2_1 _11919_ (.A(_05049_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__o32a_1 _11920_ (.A1(_04949_),
    .A2(_04954_),
    .A3(_04955_),
    .B1(_04957_),
    .B2(_04964_),
    .X(_05052_));
 sky130_fd_sc_hd__o22a_1 _11921_ (.A1(net50),
    .A2(net9),
    .B1(net4),
    .B2(net53),
    .X(_05053_));
 sky130_fd_sc_hd__xnor2_1 _11922_ (.A(net34),
    .B(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__or2_1 _11923_ (.A(net44),
    .B(_00596_),
    .X(_05055_));
 sky130_fd_sc_hd__o22a_1 _11924_ (.A1(net61),
    .A2(net15),
    .B1(net36),
    .B2(net58),
    .X(_05056_));
 sky130_fd_sc_hd__xnor2_1 _11925_ (.A(net76),
    .B(_05056_),
    .Y(_05058_));
 sky130_fd_sc_hd__nor2_1 _11926_ (.A(_05055_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _11927_ (.A(_05055_),
    .B(_05058_),
    .Y(_05060_));
 sky130_fd_sc_hd__and2b_1 _11928_ (.A_N(_05059_),
    .B(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__xnor2_1 _11929_ (.A(_05054_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__a21oi_2 _11930_ (.A1(_04971_),
    .A2(_04973_),
    .B1(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__and3_1 _11931_ (.A(_04971_),
    .B(_04973_),
    .C(_05062_),
    .X(_05064_));
 sky130_fd_sc_hd__nor2_1 _11932_ (.A(_05063_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__and2b_1 _11933_ (.A_N(_05052_),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__xnor2_1 _11934_ (.A(_05052_),
    .B(_05065_),
    .Y(_05067_));
 sky130_fd_sc_hd__and2_1 _11935_ (.A(_05051_),
    .B(_05067_),
    .X(_05069_));
 sky130_fd_sc_hd__xnor2_1 _11936_ (.A(_05051_),
    .B(_05067_),
    .Y(_05070_));
 sky130_fd_sc_hd__o21a_1 _11937_ (.A1(_04966_),
    .A2(_04978_),
    .B1(_04977_),
    .X(_05071_));
 sky130_fd_sc_hd__nor2_1 _11938_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__and2_1 _11939_ (.A(_05070_),
    .B(_05071_),
    .X(_05073_));
 sky130_fd_sc_hd__or2_1 _11940_ (.A(_05072_),
    .B(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__a21o_1 _11941_ (.A1(_04982_),
    .A2(_04985_),
    .B1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__inv_2 _11942_ (.A(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__and3_1 _11943_ (.A(_04982_),
    .B(_04985_),
    .C(_05074_),
    .X(_05077_));
 sky130_fd_sc_hd__or2_2 _11944_ (.A(_05076_),
    .B(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a21oi_1 _11945_ (.A1(_04900_),
    .A2(_04987_),
    .B1(_04988_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_04903_),
    .B(_04991_),
    .Y(_05081_));
 sky130_fd_sc_hd__o21ba_1 _11947_ (.A1(_04904_),
    .A2(_05081_),
    .B1_N(_05080_),
    .X(_05082_));
 sky130_fd_sc_hd__o31a_1 _11948_ (.A1(_04716_),
    .A2(_04906_),
    .A3(_05081_),
    .B1(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__xnor2_2 _11949_ (.A(_05078_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand2b_1 _11950_ (.A_N(_05034_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__nand2b_1 _11951_ (.A_N(_05084_),
    .B(_05034_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21ai_1 _11952_ (.A1(_02130_),
    .A2(_02131_),
    .B1(net159),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_1 _11953_ (.A(_02136_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__o211a_1 _11954_ (.A1(_02136_),
    .A2(_05087_),
    .B1(_05088_),
    .C1(net252),
    .X(_05089_));
 sky130_fd_sc_hd__o211a_1 _11955_ (.A1(_05383_),
    .A2(_05007_),
    .B1(_06372_),
    .C1(net309),
    .X(_05091_));
 sky130_fd_sc_hd__a21o_1 _11956_ (.A1(_05383_),
    .A2(_05006_),
    .B1(_05361_),
    .X(_05092_));
 sky130_fd_sc_hd__a21o_1 _11957_ (.A1(net303),
    .A2(_05092_),
    .B1(_05091_),
    .X(_05093_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_05307_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__or2_1 _11959_ (.A(_05307_),
    .B(_05093_),
    .X(_05095_));
 sky130_fd_sc_hd__or2_1 _11960_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .X(_05096_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .Y(_05097_));
 sky130_fd_sc_hd__nand2_1 _11962_ (.A(_05096_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__a21boi_1 _11963_ (.A1(_05010_),
    .A2(_05013_),
    .B1_N(_05011_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_1 _11964_ (.A(_05098_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(_03481_),
    .A1(_05100_),
    .S(net268),
    .X(_05102_));
 sky130_fd_sc_hd__or2_1 _11966_ (.A(\div_res[22] ),
    .B(_05021_),
    .X(_05103_));
 sky130_fd_sc_hd__a21oi_1 _11967_ (.A1(net164),
    .A2(_05103_),
    .B1(\div_res[23] ),
    .Y(_05104_));
 sky130_fd_sc_hd__a31o_1 _11968_ (.A1(\div_res[23] ),
    .A2(net164),
    .A3(_05103_),
    .B1(net204),
    .X(_05105_));
 sky130_fd_sc_hd__or2_1 _11969_ (.A(_05104_),
    .B(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__or2_1 _11970_ (.A(\div_shifter[54] ),
    .B(_05018_),
    .X(_05107_));
 sky130_fd_sc_hd__a21oi_1 _11971_ (.A1(net246),
    .A2(_05107_),
    .B1(\div_shifter[55] ),
    .Y(_05108_));
 sky130_fd_sc_hd__a31o_1 _11972_ (.A1(\div_shifter[55] ),
    .A2(net246),
    .A3(_05107_),
    .B1(net251),
    .X(_05109_));
 sky130_fd_sc_hd__nand2_1 _11973_ (.A(_05286_),
    .B(_02255_),
    .Y(_05110_));
 sky130_fd_sc_hd__o211a_1 _11974_ (.A1(_05286_),
    .A2(net253),
    .B1(_05110_),
    .C1(net207),
    .X(_05111_));
 sky130_fd_sc_hd__o22a_1 _11975_ (.A1(_05275_),
    .A2(net215),
    .B1(_05111_),
    .B2(_05296_),
    .X(_05113_));
 sky130_fd_sc_hd__o221a_1 _11976_ (.A1(net190),
    .A2(_03470_),
    .B1(_03481_),
    .B2(net188),
    .C1(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__o211a_1 _11977_ (.A1(_05108_),
    .A2(_05109_),
    .B1(_05114_),
    .C1(_05106_),
    .X(_05115_));
 sky130_fd_sc_hd__o21ai_1 _11978_ (.A1(_06447_),
    .A2(_05102_),
    .B1(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__a311o_1 _11979_ (.A1(_02247_),
    .A2(_05094_),
    .A3(_05095_),
    .B1(_05116_),
    .C1(_05089_),
    .X(_05117_));
 sky130_fd_sc_hd__a31o_1 _11980_ (.A1(_02171_),
    .A2(_05085_),
    .A3(_05086_),
    .B1(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__a31o_1 _11981_ (.A1(curr_PC[21]),
    .A2(curr_PC[22]),
    .A3(_04850_),
    .B1(curr_PC[23]),
    .X(_05119_));
 sky130_fd_sc_hd__and3_1 _11982_ (.A(curr_PC[22]),
    .B(curr_PC[23]),
    .C(_04943_),
    .X(_05120_));
 sky130_fd_sc_hd__nor2_1 _11983_ (.A(net263),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__a22o_4 _11984_ (.A1(net262),
    .A2(_05118_),
    .B1(_05119_),
    .B2(_05121_),
    .X(dest_val[23]));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(_04998_),
    .B(_05084_),
    .Y(_05123_));
 sky130_fd_sc_hd__or3_1 _11986_ (.A(_04758_),
    .B(_04945_),
    .C(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__or3_1 _11987_ (.A(net107),
    .B(_00136_),
    .C(net6),
    .X(_05125_));
 sky130_fd_sc_hd__a2bb2o_2 _11988_ (.A1_N(_00137_),
    .A2_N(net6),
    .B1(_05125_),
    .B2(net108),
    .X(_05126_));
 sky130_fd_sc_hd__nor2_1 _11989_ (.A(net53),
    .B(net31),
    .Y(_05127_));
 sky130_fd_sc_hd__xnor2_1 _11990_ (.A(_05126_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__o21ai_1 _11991_ (.A1(_05038_),
    .A2(_05042_),
    .B1(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__or3_1 _11992_ (.A(_05038_),
    .B(_05042_),
    .C(_05128_),
    .X(_05130_));
 sky130_fd_sc_hd__and2_1 _11993_ (.A(_05129_),
    .B(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__a21o_1 _11994_ (.A1(_05054_),
    .A2(_05060_),
    .B1(_05059_),
    .X(_05132_));
 sky130_fd_sc_hd__o22a_1 _11995_ (.A1(net58),
    .A2(net15),
    .B1(net36),
    .B2(net56),
    .X(_05134_));
 sky130_fd_sc_hd__xnor2_1 _11996_ (.A(net76),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o22a_1 _11997_ (.A1(net61),
    .A2(net9),
    .B1(net4),
    .B2(net50),
    .X(_05136_));
 sky130_fd_sc_hd__xnor2_1 _11998_ (.A(net34),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__o22a_1 _11999_ (.A1(net29),
    .A2(net17),
    .B1(net12),
    .B2(net27),
    .X(_05138_));
 sky130_fd_sc_hd__xnor2_1 _12000_ (.A(net111),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__and2_1 _12001_ (.A(_05137_),
    .B(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__nor2_1 _12002_ (.A(_05137_),
    .B(_05139_),
    .Y(_05141_));
 sky130_fd_sc_hd__or2_1 _12003_ (.A(_05140_),
    .B(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__nor2_1 _12004_ (.A(_05135_),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__and2_1 _12005_ (.A(_05135_),
    .B(_05142_),
    .X(_05145_));
 sky130_fd_sc_hd__nor2_1 _12006_ (.A(_05143_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__and2_1 _12007_ (.A(_05132_),
    .B(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__inv_2 _12008_ (.A(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__nor2_1 _12009_ (.A(_05132_),
    .B(_05146_),
    .Y(_05149_));
 sky130_fd_sc_hd__or2_1 _12010_ (.A(_05147_),
    .B(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a21o_1 _12011_ (.A1(_05045_),
    .A2(_05049_),
    .B1(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__nand3_1 _12012_ (.A(_05045_),
    .B(_05049_),
    .C(_05150_),
    .Y(_05152_));
 sky130_fd_sc_hd__nand3_2 _12013_ (.A(_05131_),
    .B(_05151_),
    .C(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21o_1 _12014_ (.A1(_05151_),
    .A2(_05152_),
    .B1(_05131_),
    .X(_05154_));
 sky130_fd_sc_hd__o211ai_4 _12015_ (.A1(_05063_),
    .A2(_05066_),
    .B1(_05153_),
    .C1(_05154_),
    .Y(_05156_));
 sky130_fd_sc_hd__a211o_1 _12016_ (.A1(_05153_),
    .A2(_05154_),
    .B1(_05063_),
    .C1(_05066_),
    .X(_05157_));
 sky130_fd_sc_hd__o211a_1 _12017_ (.A1(_05069_),
    .A2(_05072_),
    .B1(_05156_),
    .C1(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__a211o_1 _12018_ (.A1(_05156_),
    .A2(_05157_),
    .B1(_05069_),
    .C1(_05072_),
    .X(_05159_));
 sky130_fd_sc_hd__nand2b_2 _12019_ (.A_N(_05158_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__a21oi_2 _12020_ (.A1(_04987_),
    .A2(_05075_),
    .B1(_05077_),
    .Y(_05161_));
 sky130_fd_sc_hd__inv_2 _12021_ (.A(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__nor2_1 _12022_ (.A(_04990_),
    .B(_05078_),
    .Y(_05163_));
 sky130_fd_sc_hd__a21o_1 _12023_ (.A1(_04993_),
    .A2(_05163_),
    .B1(_05161_),
    .X(_05164_));
 sky130_fd_sc_hd__or3_1 _12024_ (.A(_04990_),
    .B(_04994_),
    .C(_05078_),
    .X(_05165_));
 sky130_fd_sc_hd__inv_2 _12025_ (.A(_05165_),
    .Y(_05167_));
 sky130_fd_sc_hd__and2b_1 _12026_ (.A_N(_05165_),
    .B(_04814_),
    .X(_05168_));
 sky130_fd_sc_hd__a311oi_4 _12027_ (.A1(_04403_),
    .A2(_04815_),
    .A3(_05167_),
    .B1(_05168_),
    .C1(_05164_),
    .Y(_05169_));
 sky130_fd_sc_hd__xor2_2 _12028_ (.A(_05160_),
    .B(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__a21o_1 _12029_ (.A1(net160),
    .A2(_05124_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nand3_1 _12030_ (.A(net160),
    .B(_05124_),
    .C(_05170_),
    .Y(_05172_));
 sky130_fd_sc_hd__or3_1 _12031_ (.A(net156),
    .B(_02137_),
    .C(_02138_),
    .X(_05173_));
 sky130_fd_sc_hd__o21ai_1 _12032_ (.A1(net156),
    .A2(_02137_),
    .B1(_02138_),
    .Y(_05174_));
 sky130_fd_sc_hd__a21oi_1 _12033_ (.A1(_05307_),
    .A2(_05092_),
    .B1(_05286_),
    .Y(_05175_));
 sky130_fd_sc_hd__mux2_1 _12034_ (.A0(_06379_),
    .A1(_05175_),
    .S(net304),
    .X(_05176_));
 sky130_fd_sc_hd__a21oi_1 _12035_ (.A1(_05209_),
    .A2(_05176_),
    .B1(net255),
    .Y(_05178_));
 sky130_fd_sc_hd__o21a_1 _12036_ (.A1(_05209_),
    .A2(_05176_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__o21a_1 _12037_ (.A1(_05098_),
    .A2(_05099_),
    .B1(_05097_),
    .X(_05180_));
 sky130_fd_sc_hd__nor2_1 _12038_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _12039_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05182_));
 sky130_fd_sc_hd__and2b_1 _12040_ (.A_N(_05181_),
    .B(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__xnor2_1 _12041_ (.A(_05180_),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__mux2_1 _12042_ (.A0(_03330_),
    .A1(_05184_),
    .S(net268),
    .X(_05185_));
 sky130_fd_sc_hd__or2_1 _12043_ (.A(\div_res[23] ),
    .B(_05103_),
    .X(_05186_));
 sky130_fd_sc_hd__a21oi_1 _12044_ (.A1(net164),
    .A2(_05186_),
    .B1(\div_res[24] ),
    .Y(_05187_));
 sky130_fd_sc_hd__a31o_1 _12045_ (.A1(\div_res[24] ),
    .A2(net164),
    .A3(_05186_),
    .B1(net205),
    .X(_05189_));
 sky130_fd_sc_hd__or2_1 _12046_ (.A(\div_shifter[55] ),
    .B(_05107_),
    .X(_05190_));
 sky130_fd_sc_hd__a21oi_1 _12047_ (.A1(net246),
    .A2(_05190_),
    .B1(\div_shifter[56] ),
    .Y(_05191_));
 sky130_fd_sc_hd__a311o_1 _12048_ (.A1(\div_shifter[56] ),
    .A2(net246),
    .A3(_05190_),
    .B1(_05191_),
    .C1(net251),
    .X(_05192_));
 sky130_fd_sc_hd__mux2_1 _12049_ (.A0(_02255_),
    .A1(_02249_),
    .S(_05188_),
    .X(_05193_));
 sky130_fd_sc_hd__o22a_1 _12050_ (.A1(reg1_val[24]),
    .A2(_05177_),
    .B1(_02245_),
    .B2(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__a221o_1 _12051_ (.A1(_05177_),
    .A2(_06459_),
    .B1(_02243_),
    .B2(_03330_),
    .C1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__a21oi_1 _12052_ (.A1(net192),
    .A2(_03336_),
    .B1(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__o211ai_2 _12053_ (.A1(_05187_),
    .A2(_05189_),
    .B1(_05192_),
    .C1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a211o_1 _12054_ (.A1(net216),
    .A2(_05185_),
    .B1(_05197_),
    .C1(_05179_),
    .X(_05198_));
 sky130_fd_sc_hd__a31o_1 _12055_ (.A1(net252),
    .A2(_05173_),
    .A3(_05174_),
    .B1(_05198_),
    .X(_05200_));
 sky130_fd_sc_hd__a31o_1 _12056_ (.A1(_02171_),
    .A2(_05171_),
    .A3(_05172_),
    .B1(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(curr_PC[24]),
    .B(_05120_),
    .X(_05202_));
 sky130_fd_sc_hd__and2_2 _12058_ (.A(curr_PC[24]),
    .B(_05120_),
    .X(_05203_));
 sky130_fd_sc_hd__nor2_1 _12059_ (.A(net266),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__a22o_4 _12060_ (.A1(net266),
    .A2(_05201_),
    .B1(_05202_),
    .B2(_05204_),
    .X(dest_val[24]));
 sky130_fd_sc_hd__o21a_1 _12061_ (.A1(_05124_),
    .A2(_05170_),
    .B1(net160),
    .X(_05205_));
 sky130_fd_sc_hd__o22a_1 _12062_ (.A1(net58),
    .A2(net9),
    .B1(net4),
    .B2(net61),
    .X(_05206_));
 sky130_fd_sc_hd__xnor2_1 _12063_ (.A(net34),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__nand2_1 _12064_ (.A(_05126_),
    .B(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__or2_1 _12065_ (.A(_05126_),
    .B(_05207_),
    .X(_05210_));
 sky130_fd_sc_hd__nand2_1 _12066_ (.A(_05208_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__nor2_1 _12067_ (.A(net50),
    .B(net31),
    .Y(_05212_));
 sky130_fd_sc_hd__xnor2_1 _12068_ (.A(_05211_),
    .B(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__o31a_1 _12069_ (.A1(net53),
    .A2(net31),
    .A3(_05126_),
    .B1(_05129_),
    .X(_05214_));
 sky130_fd_sc_hd__o22a_1 _12070_ (.A1(net56),
    .A2(net15),
    .B1(net36),
    .B2(net17),
    .X(_05215_));
 sky130_fd_sc_hd__xnor2_1 _12071_ (.A(net76),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nor2_1 _12072_ (.A(net109),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__and2_1 _12073_ (.A(net109),
    .B(_05216_),
    .X(_05218_));
 sky130_fd_sc_hd__nor2_1 _12074_ (.A(_05217_),
    .B(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__o22a_1 _12075_ (.A1(net29),
    .A2(net12),
    .B1(net8),
    .B2(net27),
    .X(_05221_));
 sky130_fd_sc_hd__xnor2_1 _12076_ (.A(net112),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__and2_1 _12077_ (.A(_05219_),
    .B(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__nor2_1 _12078_ (.A(_05219_),
    .B(_05222_),
    .Y(_05224_));
 sky130_fd_sc_hd__nor2_1 _12079_ (.A(_05223_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__o21ai_1 _12080_ (.A1(_05140_),
    .A2(_05143_),
    .B1(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__or3_1 _12081_ (.A(_05140_),
    .B(_05143_),
    .C(_05225_),
    .X(_05227_));
 sky130_fd_sc_hd__and2_1 _12082_ (.A(_05226_),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__nand2b_1 _12083_ (.A_N(_05214_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__xnor2_1 _12084_ (.A(_05214_),
    .B(_05228_),
    .Y(_05230_));
 sky130_fd_sc_hd__nand2_1 _12085_ (.A(_05213_),
    .B(_05230_),
    .Y(_05232_));
 sky130_fd_sc_hd__or2_1 _12086_ (.A(_05213_),
    .B(_05230_),
    .X(_05233_));
 sky130_fd_sc_hd__nand2_1 _12087_ (.A(_05232_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__a21o_1 _12088_ (.A1(_05148_),
    .A2(_05151_),
    .B1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__nand3_1 _12089_ (.A(_05148_),
    .B(_05151_),
    .C(_05234_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _12090_ (.A(_05235_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__a21o_1 _12091_ (.A1(_05153_),
    .A2(_05156_),
    .B1(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__inv_2 _12092_ (.A(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__nand3_1 _12093_ (.A(_05153_),
    .B(_05156_),
    .C(_05237_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_2 _12094_ (.A(_05238_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__o21a_1 _12095_ (.A1(_05076_),
    .A2(_05158_),
    .B1(_05159_),
    .X(_05243_));
 sky130_fd_sc_hd__nor2_1 _12096_ (.A(_05078_),
    .B(_05160_),
    .Y(_05244_));
 sky130_fd_sc_hd__a21o_1 _12097_ (.A1(_05080_),
    .A2(_05244_),
    .B1(_05243_),
    .X(_05245_));
 sky130_fd_sc_hd__and3_1 _12098_ (.A(_04903_),
    .B(_04991_),
    .C(_05244_),
    .X(_05246_));
 sky130_fd_sc_hd__and2_1 _12099_ (.A(_04907_),
    .B(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__a311oi_4 _12100_ (.A1(_04515_),
    .A2(_04908_),
    .A3(_05246_),
    .B1(_05247_),
    .C1(_05245_),
    .Y(_05248_));
 sky130_fd_sc_hd__xnor2_2 _12101_ (.A(_05241_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__inv_2 _12102_ (.A(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__nor2_1 _12103_ (.A(_05205_),
    .B(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__a21o_1 _12104_ (.A1(_05205_),
    .A2(_05250_),
    .B1(net209),
    .X(_05252_));
 sky130_fd_sc_hd__a21oi_1 _12105_ (.A1(_02137_),
    .A2(_02138_),
    .B1(net156),
    .Y(_05254_));
 sky130_fd_sc_hd__nor2_1 _12106_ (.A(_02142_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__a211o_1 _12107_ (.A1(_02142_),
    .A2(_05254_),
    .B1(_05255_),
    .C1(_02254_),
    .X(_05256_));
 sky130_fd_sc_hd__o21a_1 _12108_ (.A1(_05209_),
    .A2(_05175_),
    .B1(_05188_),
    .X(_05257_));
 sky130_fd_sc_hd__mux2_1 _12109_ (.A0(_06398_),
    .A1(_05257_),
    .S(net303),
    .X(_05258_));
 sky130_fd_sc_hd__nor2_1 _12110_ (.A(_05068_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__a211o_1 _12111_ (.A1(_05068_),
    .A2(_05258_),
    .B1(_05259_),
    .C1(net255),
    .X(_05260_));
 sky130_fd_sc_hd__o21ai_2 _12112_ (.A1(_05180_),
    .A2(_05181_),
    .B1(_05182_),
    .Y(_05261_));
 sky130_fd_sc_hd__nor2_1 _12113_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05262_));
 sky130_fd_sc_hd__or2_1 _12114_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .X(_05263_));
 sky130_fd_sc_hd__and2_1 _12115_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .X(_05265_));
 sky130_fd_sc_hd__o21ai_1 _12116_ (.A1(_05262_),
    .A2(_05265_),
    .B1(_05261_),
    .Y(_05266_));
 sky130_fd_sc_hd__o31a_1 _12117_ (.A1(_05261_),
    .A2(_05262_),
    .A3(_05265_),
    .B1(net268),
    .X(_05267_));
 sky130_fd_sc_hd__a22o_1 _12118_ (.A1(net244),
    .A2(_03197_),
    .B1(_05266_),
    .B2(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__or2_1 _12119_ (.A(\div_shifter[56] ),
    .B(_05190_),
    .X(_05269_));
 sky130_fd_sc_hd__a21oi_1 _12120_ (.A1(net246),
    .A2(_05269_),
    .B1(\div_shifter[57] ),
    .Y(_05270_));
 sky130_fd_sc_hd__a31o_1 _12121_ (.A1(\div_shifter[57] ),
    .A2(net246),
    .A3(_05269_),
    .B1(net251),
    .X(_05271_));
 sky130_fd_sc_hd__or2_1 _12122_ (.A(_05270_),
    .B(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__or2_1 _12123_ (.A(\div_res[24] ),
    .B(_05186_),
    .X(_05273_));
 sky130_fd_sc_hd__a21oi_1 _12124_ (.A1(net164),
    .A2(_05273_),
    .B1(\div_res[25] ),
    .Y(_05274_));
 sky130_fd_sc_hd__a31o_1 _12125_ (.A1(\div_res[25] ),
    .A2(net164),
    .A3(_05273_),
    .B1(net205),
    .X(_05276_));
 sky130_fd_sc_hd__mux2_1 _12126_ (.A0(net254),
    .A1(net206),
    .S(_05046_),
    .X(_05277_));
 sky130_fd_sc_hd__a21o_1 _12127_ (.A1(net207),
    .A2(_05277_),
    .B1(_05057_),
    .X(_05278_));
 sky130_fd_sc_hd__o221a_1 _12128_ (.A1(_05035_),
    .A2(net215),
    .B1(net188),
    .B2(_03197_),
    .C1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__a21boi_1 _12129_ (.A1(net192),
    .A2(_03204_),
    .B1_N(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__o211a_1 _12130_ (.A1(_05274_),
    .A2(_05276_),
    .B1(_05280_),
    .C1(_05272_),
    .X(_05281_));
 sky130_fd_sc_hd__o211a_1 _12131_ (.A1(_06447_),
    .A2(_05268_),
    .B1(_05281_),
    .C1(_05260_),
    .X(_05282_));
 sky130_fd_sc_hd__o211a_1 _12132_ (.A1(_05251_),
    .A2(_05252_),
    .B1(_05256_),
    .C1(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__a21oi_1 _12133_ (.A1(curr_PC[25]),
    .A2(_05203_),
    .B1(net266),
    .Y(_05284_));
 sky130_fd_sc_hd__o21ai_1 _12134_ (.A1(curr_PC[25]),
    .A2(_05203_),
    .B1(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__o21ai_4 _12135_ (.A1(_06424_),
    .A2(_05283_),
    .B1(_05285_),
    .Y(dest_val[25]));
 sky130_fd_sc_hd__a21bo_1 _12136_ (.A1(_05210_),
    .A2(_05212_),
    .B1_N(_05208_),
    .X(_05287_));
 sky130_fd_sc_hd__o22a_1 _12137_ (.A1(net17),
    .A2(net15),
    .B1(net36),
    .B2(net12),
    .X(_05288_));
 sky130_fd_sc_hd__xnor2_1 _12138_ (.A(_00348_),
    .B(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_1 _12139_ (.A(_06534_),
    .B(_00510_),
    .Y(_05290_));
 sky130_fd_sc_hd__a22o_1 _12140_ (.A1(_06533_),
    .A2(_00510_),
    .B1(_05290_),
    .B2(net112),
    .X(_05291_));
 sky130_fd_sc_hd__nor2_1 _12141_ (.A(_05289_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__and2_1 _12142_ (.A(_05289_),
    .B(_05291_),
    .X(_05293_));
 sky130_fd_sc_hd__or2_1 _12143_ (.A(_05292_),
    .B(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__o21ai_2 _12144_ (.A1(_05217_),
    .A2(_05223_),
    .B1(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__or3_1 _12145_ (.A(_05217_),
    .B(_05223_),
    .C(_05294_),
    .X(_05297_));
 sky130_fd_sc_hd__and2_1 _12146_ (.A(_05295_),
    .B(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_05287_),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__xnor2_1 _12148_ (.A(_05287_),
    .B(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__o22ai_2 _12149_ (.A1(net56),
    .A2(net9),
    .B1(net4),
    .B2(net58),
    .Y(_05301_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(net61),
    .B(net34),
    .Y(_05302_));
 sky130_fd_sc_hd__xor2_1 _12151_ (.A(_05301_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__or2_1 _12152_ (.A(_05300_),
    .B(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__nand2_1 _12153_ (.A(_05300_),
    .B(_05303_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_1 _12154_ (.A(_05304_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__a21o_1 _12155_ (.A1(_05226_),
    .A2(_05229_),
    .B1(_05306_),
    .X(_05308_));
 sky130_fd_sc_hd__nand3_1 _12156_ (.A(_05226_),
    .B(_05229_),
    .C(_05306_),
    .Y(_05309_));
 sky130_fd_sc_hd__nand2_1 _12157_ (.A(_05308_),
    .B(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__a21oi_1 _12158_ (.A1(_05232_),
    .A2(_05235_),
    .B1(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__and3_1 _12159_ (.A(_05232_),
    .B(_05235_),
    .C(_05310_),
    .X(_05312_));
 sky130_fd_sc_hd__or2_2 _12160_ (.A(_05311_),
    .B(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__o21ai_1 _12161_ (.A1(_05158_),
    .A2(_05239_),
    .B1(_05240_),
    .Y(_05314_));
 sky130_fd_sc_hd__or2_1 _12162_ (.A(_05160_),
    .B(_05241_),
    .X(_05315_));
 sky130_fd_sc_hd__o21ai_1 _12163_ (.A1(_05162_),
    .A2(_05315_),
    .B1(_05314_),
    .Y(_05316_));
 sky130_fd_sc_hd__inv_2 _12164_ (.A(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__or3_1 _12165_ (.A(_04990_),
    .B(_05078_),
    .C(_05315_),
    .X(_05319_));
 sky130_fd_sc_hd__o21ai_1 _12166_ (.A1(_04997_),
    .A2(_05319_),
    .B1(_05317_),
    .Y(_05320_));
 sky130_fd_sc_hd__xnor2_2 _12167_ (.A(_05313_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__nand2b_1 _12168_ (.A_N(_05170_),
    .B(_05249_),
    .Y(_05322_));
 sky130_fd_sc_hd__or4_4 _12169_ (.A(_04758_),
    .B(_04945_),
    .C(_05123_),
    .D(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__and3_1 _12170_ (.A(net160),
    .B(_05321_),
    .C(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__a21oi_1 _12171_ (.A1(net160),
    .A2(_05323_),
    .B1(_05321_),
    .Y(_05325_));
 sky130_fd_sc_hd__or3_1 _12172_ (.A(net209),
    .B(_05324_),
    .C(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__o21ba_1 _12173_ (.A1(_05068_),
    .A2(_05257_),
    .B1_N(_05046_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(_06399_),
    .A1(_05327_),
    .S(net303),
    .X(_05328_));
 sky130_fd_sc_hd__nor2_1 _12175_ (.A(_05133_),
    .B(_05328_),
    .Y(_05330_));
 sky130_fd_sc_hd__nor2_1 _12176_ (.A(_05133_),
    .B(_05327_),
    .Y(_05331_));
 sky130_fd_sc_hd__a211o_1 _12177_ (.A1(_05133_),
    .A2(_05328_),
    .B1(_05330_),
    .C1(net255),
    .X(_05332_));
 sky130_fd_sc_hd__a21oi_1 _12178_ (.A1(net160),
    .A2(_02143_),
    .B1(_02144_),
    .Y(_05333_));
 sky130_fd_sc_hd__a31o_1 _12179_ (.A1(net160),
    .A2(_02143_),
    .A3(_02144_),
    .B1(_02254_),
    .X(_05334_));
 sky130_fd_sc_hd__or2_1 _12180_ (.A(_05333_),
    .B(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(_05261_),
    .A2(_05263_),
    .B1(_05265_),
    .Y(_05336_));
 sky130_fd_sc_hd__nor2_1 _12182_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_1 _12183_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2b_1 _12184_ (.A_N(_05337_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__xnor2_1 _12185_ (.A(_05336_),
    .B(_05339_),
    .Y(_05341_));
 sky130_fd_sc_hd__mux2_1 _12186_ (.A0(_03053_),
    .A1(_05341_),
    .S(net269),
    .X(_05342_));
 sky130_fd_sc_hd__or2_1 _12187_ (.A(\div_shifter[57] ),
    .B(_05269_),
    .X(_05343_));
 sky130_fd_sc_hd__a21oi_1 _12188_ (.A1(net246),
    .A2(_05343_),
    .B1(\div_shifter[58] ),
    .Y(_05344_));
 sky130_fd_sc_hd__a31o_1 _12189_ (.A1(\div_shifter[58] ),
    .A2(net246),
    .A3(_05343_),
    .B1(net251),
    .X(_05345_));
 sky130_fd_sc_hd__or2_1 _12190_ (.A(_05344_),
    .B(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__or2_1 _12191_ (.A(\div_res[25] ),
    .B(_05273_),
    .X(_05347_));
 sky130_fd_sc_hd__a21oi_1 _12192_ (.A1(net164),
    .A2(_05347_),
    .B1(\div_res[26] ),
    .Y(_05348_));
 sky130_fd_sc_hd__a31o_1 _12193_ (.A1(\div_res[26] ),
    .A2(net164),
    .A3(_05347_),
    .B1(net205),
    .X(_05349_));
 sky130_fd_sc_hd__nor2_1 _12194_ (.A(_05348_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__mux2_1 _12195_ (.A0(net254),
    .A1(net206),
    .S(_05112_),
    .X(_05352_));
 sky130_fd_sc_hd__a21o_1 _12196_ (.A1(net208),
    .A2(_05352_),
    .B1(_05122_),
    .X(_05353_));
 sky130_fd_sc_hd__o221ai_1 _12197_ (.A1(_05101_),
    .A2(net215),
    .B1(net188),
    .B2(_03053_),
    .C1(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__a211oi_1 _12198_ (.A1(net192),
    .A2(_03064_),
    .B1(_05350_),
    .C1(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__o211a_1 _12199_ (.A1(_06447_),
    .A2(_05342_),
    .B1(_05346_),
    .C1(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__a41o_1 _12200_ (.A1(_05326_),
    .A2(_05332_),
    .A3(_05335_),
    .A4(_05356_),
    .B1(_06424_),
    .X(_05357_));
 sky130_fd_sc_hd__and3_1 _12201_ (.A(curr_PC[25]),
    .B(curr_PC[26]),
    .C(_05203_),
    .X(_05358_));
 sky130_fd_sc_hd__a21oi_2 _12202_ (.A1(curr_PC[25]),
    .A2(_05203_),
    .B1(curr_PC[26]),
    .Y(_05359_));
 sky130_fd_sc_hd__o31ai_4 _12203_ (.A1(net266),
    .A2(_05358_),
    .A3(_05359_),
    .B1(_05357_),
    .Y(dest_val[26]));
 sky130_fd_sc_hd__xor2_1 _12204_ (.A(curr_PC[27]),
    .B(_05358_),
    .X(_05360_));
 sky130_fd_sc_hd__o21ai_1 _12205_ (.A1(_05321_),
    .A2(_05323_),
    .B1(net160),
    .Y(_05362_));
 sky130_fd_sc_hd__o22a_1 _12206_ (.A1(net16),
    .A2(net12),
    .B1(net8),
    .B2(net37),
    .X(_05363_));
 sky130_fd_sc_hd__xnor2_1 _12207_ (.A(net76),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__o22a_1 _12208_ (.A1(net17),
    .A2(net9),
    .B1(net4),
    .B2(net56),
    .X(_05365_));
 sky130_fd_sc_hd__xnor2_1 _12209_ (.A(net34),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__xnor2_1 _12210_ (.A(net111),
    .B(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__and2b_1 _12211_ (.A_N(_05364_),
    .B(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__xnor2_1 _12212_ (.A(_05364_),
    .B(_05367_),
    .Y(_05369_));
 sky130_fd_sc_hd__nor2_1 _12213_ (.A(net58),
    .B(net31),
    .Y(_05370_));
 sky130_fd_sc_hd__or3_1 _12214_ (.A(net62),
    .B(net31),
    .C(_05301_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _12215_ (.A0(net58),
    .A1(_05370_),
    .S(_05371_),
    .X(_05373_));
 sky130_fd_sc_hd__inv_2 _12216_ (.A(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__xnor2_1 _12217_ (.A(_05292_),
    .B(_05373_),
    .Y(_05375_));
 sky130_fd_sc_hd__and2_1 _12218_ (.A(_05369_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__nor2_1 _12219_ (.A(_05369_),
    .B(_05375_),
    .Y(_05377_));
 sky130_fd_sc_hd__a211oi_2 _12220_ (.A1(_05295_),
    .A2(_05299_),
    .B1(_05376_),
    .C1(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__o211a_1 _12221_ (.A1(_05376_),
    .A2(_05377_),
    .B1(_05295_),
    .C1(_05299_),
    .X(_05379_));
 sky130_fd_sc_hd__a211oi_1 _12222_ (.A1(_05304_),
    .A2(_05308_),
    .B1(_05378_),
    .C1(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__o211ai_2 _12223_ (.A1(_05378_),
    .A2(_05379_),
    .B1(_05304_),
    .C1(_05308_),
    .Y(_05381_));
 sky130_fd_sc_hd__nand2b_2 _12224_ (.A_N(_05380_),
    .B(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__o21ba_1 _12225_ (.A1(_05239_),
    .A2(_05311_),
    .B1_N(_05312_),
    .X(_05384_));
 sky130_fd_sc_hd__nor2_1 _12226_ (.A(_05241_),
    .B(_05313_),
    .Y(_05385_));
 sky130_fd_sc_hd__a21oi_1 _12227_ (.A1(_05243_),
    .A2(_05385_),
    .B1(_05384_),
    .Y(_05386_));
 sky130_fd_sc_hd__nand2_1 _12228_ (.A(_05244_),
    .B(_05385_),
    .Y(_05387_));
 sky130_fd_sc_hd__o21a_1 _12229_ (.A1(_05083_),
    .A2(_05387_),
    .B1(_05386_),
    .X(_05388_));
 sky130_fd_sc_hd__xnor2_2 _12230_ (.A(_05382_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__o21ai_1 _12231_ (.A1(_05362_),
    .A2(_05389_),
    .B1(_02171_),
    .Y(_05390_));
 sky130_fd_sc_hd__a21oi_1 _12232_ (.A1(_05362_),
    .A2(_05389_),
    .B1(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _12233_ (.A(net310),
    .B(_06400_),
    .Y(_05392_));
 sky130_fd_sc_hd__o31ai_1 _12234_ (.A1(net309),
    .A2(_05112_),
    .A3(_05331_),
    .B1(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__a21oi_1 _12235_ (.A1(_04774_),
    .A2(_05393_),
    .B1(net255),
    .Y(_05395_));
 sky130_fd_sc_hd__o21a_1 _12236_ (.A1(_04774_),
    .A2(_05393_),
    .B1(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__o21ai_1 _12237_ (.A1(_02143_),
    .A2(_02144_),
    .B1(net160),
    .Y(_05397_));
 sky130_fd_sc_hd__xnor2_1 _12238_ (.A(_02149_),
    .B(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__o21a_1 _12239_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_05338_),
    .X(_05399_));
 sky130_fd_sc_hd__nor2_1 _12240_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _12241_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05401_));
 sky130_fd_sc_hd__nand2b_1 _12242_ (.A_N(_05400_),
    .B(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__xnor2_1 _12243_ (.A(_05399_),
    .B(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(_02908_),
    .A1(_05403_),
    .S(net268),
    .X(_05404_));
 sky130_fd_sc_hd__or2_1 _12245_ (.A(\div_shifter[58] ),
    .B(_05343_),
    .X(_05406_));
 sky130_fd_sc_hd__a21oi_1 _12246_ (.A1(_02445_),
    .A2(_05406_),
    .B1(\div_shifter[59] ),
    .Y(_05407_));
 sky130_fd_sc_hd__a311o_1 _12247_ (.A1(\div_shifter[59] ),
    .A2(_02445_),
    .A3(_05406_),
    .B1(_05407_),
    .C1(net251),
    .X(_05408_));
 sky130_fd_sc_hd__or2_1 _12248_ (.A(\div_res[26] ),
    .B(_05347_),
    .X(_05409_));
 sky130_fd_sc_hd__a21oi_1 _12249_ (.A1(net164),
    .A2(_05409_),
    .B1(\div_res[27] ),
    .Y(_05410_));
 sky130_fd_sc_hd__a31o_1 _12250_ (.A1(\div_res[27] ),
    .A2(net164),
    .A3(_05409_),
    .B1(net205),
    .X(_05411_));
 sky130_fd_sc_hd__a21o_1 _12251_ (.A1(_04753_),
    .A2(_02249_),
    .B1(_02245_),
    .X(_05412_));
 sky130_fd_sc_hd__o221a_1 _12252_ (.A1(_04731_),
    .A2(net215),
    .B1(net206),
    .B2(_04753_),
    .C1(net266),
    .X(_05413_));
 sky130_fd_sc_hd__a21boi_1 _12253_ (.A1(_04742_),
    .A2(_05412_),
    .B1_N(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__o221a_1 _12254_ (.A1(net188),
    .A2(_02908_),
    .B1(_02915_),
    .B2(net190),
    .C1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__o211a_1 _12255_ (.A1(_05410_),
    .A2(_05411_),
    .B1(_05415_),
    .C1(_05408_),
    .X(_05417_));
 sky130_fd_sc_hd__o21ai_1 _12256_ (.A1(_06447_),
    .A2(_05404_),
    .B1(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a211o_1 _12257_ (.A1(_02253_),
    .A2(_05398_),
    .B1(_05418_),
    .C1(_05396_),
    .X(_05419_));
 sky130_fd_sc_hd__o22a_4 _12258_ (.A1(_06425_),
    .A2(_05360_),
    .B1(_05391_),
    .B2(_05419_),
    .X(dest_val[27]));
 sky130_fd_sc_hd__a21o_1 _12259_ (.A1(_06524_),
    .A2(_05366_),
    .B1(_05368_),
    .X(_05420_));
 sky130_fd_sc_hd__o22a_1 _12260_ (.A1(net12),
    .A2(net11),
    .B1(net5),
    .B2(net17),
    .X(_05421_));
 sky130_fd_sc_hd__xnor2_1 _12261_ (.A(net34),
    .B(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand2_1 _12262_ (.A(_05420_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__xnor2_1 _12263_ (.A(_05420_),
    .B(_05422_),
    .Y(_05424_));
 sky130_fd_sc_hd__nand2_1 _12264_ (.A(_00242_),
    .B(net35),
    .Y(_05425_));
 sky130_fd_sc_hd__or2_1 _12265_ (.A(_05424_),
    .B(_05425_),
    .X(_05427_));
 sky130_fd_sc_hd__nand2_1 _12266_ (.A(_05424_),
    .B(_05425_),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_1 _12267_ (.A(_05427_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__o21a_1 _12268_ (.A1(net16),
    .A2(net8),
    .B1(_00348_),
    .X(_05430_));
 sky130_fd_sc_hd__a41o_1 _12269_ (.A1(net111),
    .A2(net76),
    .A3(_00350_),
    .A4(_00510_),
    .B1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__or2_1 _12270_ (.A(_05429_),
    .B(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__nand2_1 _12271_ (.A(_05429_),
    .B(_05431_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand2_1 _12272_ (.A(_05432_),
    .B(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__o22ai_2 _12273_ (.A1(net59),
    .A2(_05371_),
    .B1(_05374_),
    .B2(_05292_),
    .Y(_05435_));
 sky130_fd_sc_hd__nand2b_1 _12274_ (.A_N(_05434_),
    .B(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__xnor2_1 _12275_ (.A(_05434_),
    .B(_05435_),
    .Y(_05438_));
 sky130_fd_sc_hd__o21a_1 _12276_ (.A1(_05376_),
    .A2(_05378_),
    .B1(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__or3_1 _12277_ (.A(_05376_),
    .B(_05378_),
    .C(_05438_),
    .X(_05440_));
 sky130_fd_sc_hd__nand2b_1 _12278_ (.A_N(_05439_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__inv_2 _12279_ (.A(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__or2_1 _12280_ (.A(_05313_),
    .B(_05382_),
    .X(_05443_));
 sky130_fd_sc_hd__nor2_1 _12281_ (.A(_05315_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__inv_2 _12282_ (.A(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_1 _12283_ (.A1(_05311_),
    .A2(_05380_),
    .B1(_05381_),
    .Y(_05446_));
 sky130_fd_sc_hd__o221a_1 _12284_ (.A1(_05314_),
    .A2(_05443_),
    .B1(_05445_),
    .B2(_05169_),
    .C1(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__xnor2_2 _12285_ (.A(_05442_),
    .B(_05447_),
    .Y(_05449_));
 sky130_fd_sc_hd__nand2b_2 _12286_ (.A_N(_05321_),
    .B(_05389_),
    .Y(_05450_));
 sky130_fd_sc_hd__or2_1 _12287_ (.A(_05323_),
    .B(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__a21oi_1 _12288_ (.A1(net160),
    .A2(_05451_),
    .B1(_05449_),
    .Y(_05452_));
 sky130_fd_sc_hd__o211a_1 _12289_ (.A1(_05323_),
    .A2(_05450_),
    .B1(_05449_),
    .C1(net160),
    .X(_05453_));
 sky130_fd_sc_hd__or3_1 _12290_ (.A(net209),
    .B(_05452_),
    .C(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__o31a_1 _12291_ (.A1(_04763_),
    .A2(_05112_),
    .A3(_05331_),
    .B1(_04742_),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(_06401_),
    .A1(_05455_),
    .S(net304),
    .X(_05456_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_05003_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__o211a_1 _12294_ (.A1(_05003_),
    .A2(_05456_),
    .B1(_05457_),
    .C1(_02247_),
    .X(_05458_));
 sky130_fd_sc_hd__a21oi_1 _12295_ (.A1(net161),
    .A2(_02150_),
    .B1(_02151_),
    .Y(_05460_));
 sky130_fd_sc_hd__a31o_1 _12296_ (.A1(net161),
    .A2(_02150_),
    .A3(_02151_),
    .B1(_02254_),
    .X(_05461_));
 sky130_fd_sc_hd__o21ai_2 _12297_ (.A1(_05399_),
    .A2(_05400_),
    .B1(_05401_),
    .Y(_05462_));
 sky130_fd_sc_hd__xnor2_1 _12298_ (.A(reg1_val[28]),
    .B(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__nor2_1 _12299_ (.A(net269),
    .B(_02770_),
    .Y(_05464_));
 sky130_fd_sc_hd__a211o_1 _12300_ (.A1(net269),
    .A2(_05463_),
    .B1(_05464_),
    .C1(_06447_),
    .X(_05465_));
 sky130_fd_sc_hd__or2_1 _12301_ (.A(\div_shifter[59] ),
    .B(_05406_),
    .X(_05466_));
 sky130_fd_sc_hd__a21oi_1 _12302_ (.A1(net248),
    .A2(_05466_),
    .B1(\div_shifter[60] ),
    .Y(_05467_));
 sky130_fd_sc_hd__a311o_1 _12303_ (.A1(\div_shifter[60] ),
    .A2(net248),
    .A3(_05466_),
    .B1(_05467_),
    .C1(net250),
    .X(_05468_));
 sky130_fd_sc_hd__or2_1 _12304_ (.A(\div_res[27] ),
    .B(_05409_),
    .X(_05469_));
 sky130_fd_sc_hd__a21oi_1 _12305_ (.A1(net164),
    .A2(_05469_),
    .B1(\div_res[28] ),
    .Y(_05471_));
 sky130_fd_sc_hd__a31o_1 _12306_ (.A1(\div_res[28] ),
    .A2(net164),
    .A3(_05469_),
    .B1(net205),
    .X(_05472_));
 sky130_fd_sc_hd__o21ai_1 _12307_ (.A1(_04981_),
    .A2(net254),
    .B1(net207),
    .Y(_05473_));
 sky130_fd_sc_hd__a221o_1 _12308_ (.A1(_04981_),
    .A2(_02255_),
    .B1(_05473_),
    .B2(_04992_),
    .C1(_06459_),
    .X(_05474_));
 sky130_fd_sc_hd__a221oi_2 _12309_ (.A1(net192),
    .A2(_02760_),
    .B1(_02770_),
    .B2(_02243_),
    .C1(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__o211a_1 _12310_ (.A1(_05471_),
    .A2(_05472_),
    .B1(_05475_),
    .C1(_05468_),
    .X(_05476_));
 sky130_fd_sc_hd__o211ai_1 _12311_ (.A1(_05460_),
    .A2(_05461_),
    .B1(_05465_),
    .C1(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__nor2_1 _12312_ (.A(_05458_),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__a221oi_4 _12313_ (.A1(_04970_),
    .A2(_06459_),
    .B1(_05454_),
    .B2(_05478_),
    .C1(_06424_),
    .Y(dest_val[28]));
 sky130_fd_sc_hd__o22a_1 _12314_ (.A1(net9),
    .A2(net8),
    .B1(net4),
    .B2(net12),
    .X(_05479_));
 sky130_fd_sc_hd__xnor2_1 _12315_ (.A(net32),
    .B(_05479_),
    .Y(_05481_));
 sky130_fd_sc_hd__nor2_1 _12316_ (.A(net17),
    .B(net32),
    .Y(_05482_));
 sky130_fd_sc_hd__xnor2_1 _12317_ (.A(net76),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__nor2_1 _12318_ (.A(_05481_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__and2_1 _12319_ (.A(_05481_),
    .B(_05483_),
    .X(_05485_));
 sky130_fd_sc_hd__or2_1 _12320_ (.A(_05484_),
    .B(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__and2b_1 _12321_ (.A_N(_05486_),
    .B(_05431_),
    .X(_05487_));
 sky130_fd_sc_hd__and2b_1 _12322_ (.A_N(_05431_),
    .B(_05486_),
    .X(_05488_));
 sky130_fd_sc_hd__or2_1 _12323_ (.A(_05487_),
    .B(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__a21oi_1 _12324_ (.A1(_05423_),
    .A2(_05427_),
    .B1(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__and3_1 _12325_ (.A(_05423_),
    .B(_05427_),
    .C(_05489_),
    .X(_05492_));
 sky130_fd_sc_hd__or2_1 _12326_ (.A(_05490_),
    .B(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__nand3_1 _12327_ (.A(_05432_),
    .B(_05436_),
    .C(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__inv_2 _12328_ (.A(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__a21oi_2 _12329_ (.A1(_05432_),
    .A2(_05436_),
    .B1(_05493_),
    .Y(_05496_));
 sky130_fd_sc_hd__nor2_2 _12330_ (.A(_05495_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__nor2_1 _12331_ (.A(_05382_),
    .B(_05441_),
    .Y(_05498_));
 sky130_fd_sc_hd__nand2_1 _12332_ (.A(_05385_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__o21ai_1 _12333_ (.A1(_05380_),
    .A2(_05439_),
    .B1(_05440_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_1 _12334_ (.A(_05384_),
    .B(_05498_),
    .Y(_05501_));
 sky130_fd_sc_hd__o211a_1 _12335_ (.A1(_05248_),
    .A2(_05499_),
    .B1(_05500_),
    .C1(_05501_),
    .X(_05503_));
 sky130_fd_sc_hd__xnor2_2 _12336_ (.A(_05497_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__o31a_1 _12337_ (.A1(_05323_),
    .A2(_05449_),
    .A3(_05450_),
    .B1(net160),
    .X(_05505_));
 sky130_fd_sc_hd__o21ai_1 _12338_ (.A1(_05504_),
    .A2(_05505_),
    .B1(_02171_),
    .Y(_05506_));
 sky130_fd_sc_hd__a21oi_1 _12339_ (.A1(_05504_),
    .A2(_05505_),
    .B1(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__a21o_1 _12340_ (.A1(_04992_),
    .A2(_05455_),
    .B1(_04981_),
    .X(_05508_));
 sky130_fd_sc_hd__or2_1 _12341_ (.A(net310),
    .B(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__nand2_1 _12342_ (.A(net309),
    .B(_06402_),
    .Y(_05510_));
 sky130_fd_sc_hd__a21oi_1 _12343_ (.A1(_05509_),
    .A2(_05510_),
    .B1(_04927_),
    .Y(_05511_));
 sky130_fd_sc_hd__a31o_1 _12344_ (.A1(_04927_),
    .A2(_05509_),
    .A3(_05510_),
    .B1(net255),
    .X(_05512_));
 sky130_fd_sc_hd__nor2_1 _12345_ (.A(_05511_),
    .B(_05512_),
    .Y(_05514_));
 sky130_fd_sc_hd__o21ai_1 _12346_ (.A1(net158),
    .A2(_02152_),
    .B1(_02158_),
    .Y(_05515_));
 sky130_fd_sc_hd__o311a_1 _12347_ (.A1(net158),
    .A2(_02152_),
    .A3(_02158_),
    .B1(_02253_),
    .C1(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__and3_1 _12348_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_05462_),
    .X(_05517_));
 sky130_fd_sc_hd__a21oi_1 _12349_ (.A1(reg1_val[28]),
    .A2(_05462_),
    .B1(reg1_val[29]),
    .Y(_05518_));
 sky130_fd_sc_hd__o21a_1 _12350_ (.A1(_05517_),
    .A2(_05518_),
    .B1(net269),
    .X(_05519_));
 sky130_fd_sc_hd__a211oi_1 _12351_ (.A1(net244),
    .A2(_02586_),
    .B1(_05519_),
    .C1(_06447_),
    .Y(_05520_));
 sky130_fd_sc_hd__or2_1 _12352_ (.A(\div_shifter[60] ),
    .B(_05466_),
    .X(_05521_));
 sky130_fd_sc_hd__a21oi_1 _12353_ (.A1(net248),
    .A2(_05521_),
    .B1(\div_shifter[61] ),
    .Y(_05522_));
 sky130_fd_sc_hd__a311o_1 _12354_ (.A1(\div_shifter[61] ),
    .A2(net248),
    .A3(_05521_),
    .B1(_05522_),
    .C1(net250),
    .X(_05523_));
 sky130_fd_sc_hd__or2_1 _12355_ (.A(\div_res[28] ),
    .B(_05469_),
    .X(_05525_));
 sky130_fd_sc_hd__a21oi_1 _12356_ (.A1(net164),
    .A2(_05525_),
    .B1(\div_res[29] ),
    .Y(_05526_));
 sky130_fd_sc_hd__a31o_1 _12357_ (.A1(\div_res[29] ),
    .A2(net164),
    .A3(_05525_),
    .B1(net205),
    .X(_05527_));
 sky130_fd_sc_hd__a21oi_1 _12358_ (.A1(_04894_),
    .A2(_02249_),
    .B1(_02245_),
    .Y(_05528_));
 sky130_fd_sc_hd__o221a_1 _12359_ (.A1(_04894_),
    .A2(net206),
    .B1(_05528_),
    .B2(_04916_),
    .C1(net215),
    .X(_05529_));
 sky130_fd_sc_hd__o221a_1 _12360_ (.A1(_02244_),
    .A2(_02586_),
    .B1(_02601_),
    .B2(net189),
    .C1(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__o211a_1 _12361_ (.A1(_05526_),
    .A2(_05527_),
    .B1(_05530_),
    .C1(_05523_),
    .X(_05531_));
 sky130_fd_sc_hd__or4b_1 _12362_ (.A(_05514_),
    .B(_05516_),
    .C(_05520_),
    .D_N(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__o221a_4 _12363_ (.A1(_04883_),
    .A2(net215),
    .B1(_05507_),
    .B2(_05532_),
    .C1(net266),
    .X(dest_val[29]));
 sky130_fd_sc_hd__a21o_1 _12364_ (.A1(net76),
    .A2(_05482_),
    .B1(_05484_),
    .X(_05533_));
 sky130_fd_sc_hd__o31a_1 _12365_ (.A1(net77),
    .A2(_00456_),
    .A3(net6),
    .B1(net32),
    .X(_05535_));
 sky130_fd_sc_hd__nor2_1 _12366_ (.A(net6),
    .B(_00600_),
    .Y(_05536_));
 sky130_fd_sc_hd__a21o_1 _12367_ (.A1(net13),
    .A2(_05536_),
    .B1(_05535_),
    .X(_05537_));
 sky130_fd_sc_hd__inv_2 _12368_ (.A(_05537_),
    .Y(_05538_));
 sky130_fd_sc_hd__o31a_1 _12369_ (.A1(net13),
    .A2(net32),
    .A3(_05536_),
    .B1(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__inv_2 _12370_ (.A(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2_1 _12371_ (.A(_05533_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__xnor2_1 _12372_ (.A(_05533_),
    .B(_05539_),
    .Y(_05542_));
 sky130_fd_sc_hd__or3_1 _12373_ (.A(_05487_),
    .B(_05490_),
    .C(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__inv_2 _12374_ (.A(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__o21a_1 _12375_ (.A1(_05487_),
    .A2(_05490_),
    .B1(_05542_),
    .X(_05546_));
 sky130_fd_sc_hd__nor2_1 _12376_ (.A(_05544_),
    .B(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__o21ai_1 _12377_ (.A1(_05317_),
    .A2(_05443_),
    .B1(_05446_),
    .Y(_05548_));
 sky130_fd_sc_hd__a21o_1 _12378_ (.A1(_05439_),
    .A2(_05494_),
    .B1(_05496_),
    .X(_05549_));
 sky130_fd_sc_hd__a31o_1 _12379_ (.A1(_05442_),
    .A2(_05497_),
    .A3(_05548_),
    .B1(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__nand4_1 _12380_ (.A(_05163_),
    .B(_05442_),
    .C(_05444_),
    .D(_05497_),
    .Y(_05551_));
 sky130_fd_sc_hd__o21ba_1 _12381_ (.A1(_04997_),
    .A2(_05551_),
    .B1_N(_05550_),
    .X(_05552_));
 sky130_fd_sc_hd__xnor2_2 _12382_ (.A(_05547_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__or2_1 _12383_ (.A(_05449_),
    .B(_05504_),
    .X(_05554_));
 sky130_fd_sc_hd__o31a_1 _12384_ (.A1(_05323_),
    .A2(_05450_),
    .A3(_05554_),
    .B1(net160),
    .X(_05555_));
 sky130_fd_sc_hd__a21oi_1 _12385_ (.A1(_05553_),
    .A2(_05555_),
    .B1(net209),
    .Y(_05557_));
 sky130_fd_sc_hd__o21a_1 _12386_ (.A1(_05553_),
    .A2(_05555_),
    .B1(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__a21bo_1 _12387_ (.A1(_04905_),
    .A2(_05508_),
    .B1_N(_04894_),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(_06403_),
    .A1(_05559_),
    .S(net304),
    .X(_05560_));
 sky130_fd_sc_hd__nand2_1 _12389_ (.A(_04851_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21a_1 _12390_ (.A1(_04851_),
    .A2(_05560_),
    .B1(_02247_),
    .X(_05562_));
 sky130_fd_sc_hd__a21o_1 _12391_ (.A1(_02152_),
    .A2(_02158_),
    .B1(net158),
    .X(_05563_));
 sky130_fd_sc_hd__xor2_1 _12392_ (.A(_02160_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__xor2_1 _12393_ (.A(reg1_val[30]),
    .B(_05517_),
    .X(_05565_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(net244),
    .B(_02459_),
    .Y(_05566_));
 sky130_fd_sc_hd__o211a_1 _12395_ (.A1(net244),
    .A2(_05565_),
    .B1(_05566_),
    .C1(_06446_),
    .X(_05568_));
 sky130_fd_sc_hd__or2_1 _12396_ (.A(\div_shifter[61] ),
    .B(_05521_),
    .X(_05569_));
 sky130_fd_sc_hd__a21oi_1 _12397_ (.A1(net248),
    .A2(_05569_),
    .B1(\div_shifter[62] ),
    .Y(_05570_));
 sky130_fd_sc_hd__a31o_1 _12398_ (.A1(\div_shifter[62] ),
    .A2(net248),
    .A3(_05569_),
    .B1(net250),
    .X(_05571_));
 sky130_fd_sc_hd__or2_1 _12399_ (.A(\div_res[29] ),
    .B(_05525_),
    .X(_05572_));
 sky130_fd_sc_hd__a21oi_1 _12400_ (.A1(_02070_),
    .A2(_05572_),
    .B1(\div_res[30] ),
    .Y(_05573_));
 sky130_fd_sc_hd__a31o_1 _12401_ (.A1(\div_res[30] ),
    .A2(net164),
    .A3(_05572_),
    .B1(net205),
    .X(_05574_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(net254),
    .A1(_02256_),
    .S(_04829_),
    .X(_05575_));
 sky130_fd_sc_hd__a21oi_1 _12403_ (.A1(net208),
    .A2(_05575_),
    .B1(_04840_),
    .Y(_05576_));
 sky130_fd_sc_hd__nor2_1 _12404_ (.A(_06459_),
    .B(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__o221a_1 _12405_ (.A1(_02175_),
    .A2(_02431_),
    .B1(_02459_),
    .B2(_02244_),
    .C1(_05577_),
    .X(_05579_));
 sky130_fd_sc_hd__o21a_1 _12406_ (.A1(_05573_),
    .A2(_05574_),
    .B1(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__o21ai_2 _12407_ (.A1(_05570_),
    .A2(_05571_),
    .B1(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__a211o_1 _12408_ (.A1(net252),
    .A2(_05564_),
    .B1(_05568_),
    .C1(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__a21o_1 _12409_ (.A1(_05561_),
    .A2(_05562_),
    .B1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__o221a_4 _12410_ (.A1(_04807_),
    .A2(_06460_),
    .B1(_05558_),
    .B2(_05583_),
    .C1(net266),
    .X(dest_val[30]));
 sky130_fd_sc_hd__o41a_1 _12411_ (.A1(_05323_),
    .A2(_05450_),
    .A3(_05553_),
    .A4(_05554_),
    .B1(net160),
    .X(_05584_));
 sky130_fd_sc_hd__nor2_1 _12412_ (.A(_00510_),
    .B(_00596_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_05497_),
    .B(_05547_),
    .Y(_05586_));
 sky130_fd_sc_hd__or3_1 _12414_ (.A(_05382_),
    .B(_05441_),
    .C(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__a21oi_1 _12415_ (.A1(_05496_),
    .A2(_05543_),
    .B1(_05546_),
    .Y(_05589_));
 sky130_fd_sc_hd__o221a_1 _12416_ (.A1(_05500_),
    .A2(_05586_),
    .B1(_05587_),
    .B2(_05388_),
    .C1(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__xnor2_1 _12417_ (.A(_05585_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(_05533_),
    .A1(_05541_),
    .S(_05538_),
    .X(_05592_));
 sky130_fd_sc_hd__xnor2_1 _12419_ (.A(_05591_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__a21oi_1 _12420_ (.A1(_05584_),
    .A2(_05593_),
    .B1(net209),
    .Y(_05594_));
 sky130_fd_sc_hd__o21a_1 _12421_ (.A1(_05584_),
    .A2(_05593_),
    .B1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a211o_1 _12422_ (.A1(_04851_),
    .A2(_05559_),
    .B1(net309),
    .C1(_04829_),
    .X(_05596_));
 sky130_fd_sc_hd__nand2_1 _12423_ (.A(net309),
    .B(_06404_),
    .Y(_05597_));
 sky130_fd_sc_hd__a21oi_1 _12424_ (.A1(_05596_),
    .A2(_05597_),
    .B1(_04698_),
    .Y(_05598_));
 sky130_fd_sc_hd__a31o_1 _12425_ (.A1(_04698_),
    .A2(_05596_),
    .A3(_05597_),
    .B1(_02248_),
    .X(_05600_));
 sky130_fd_sc_hd__or3_1 _12426_ (.A(net158),
    .B(_02161_),
    .C(_02166_),
    .X(_05601_));
 sky130_fd_sc_hd__o21ai_1 _12427_ (.A1(net158),
    .A2(_02161_),
    .B1(_02166_),
    .Y(_05602_));
 sky130_fd_sc_hd__and3_1 _12428_ (.A(_02253_),
    .B(_05601_),
    .C(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__and3_1 _12429_ (.A(reg1_val[30]),
    .B(net269),
    .C(_05517_),
    .X(_05604_));
 sky130_fd_sc_hd__xor2_1 _12430_ (.A(_02273_),
    .B(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__o21a_1 _12431_ (.A1(\div_shifter[62] ),
    .A2(_05569_),
    .B1(net247),
    .X(_05606_));
 sky130_fd_sc_hd__o21ai_1 _12432_ (.A1(\div_shifter[63] ),
    .A2(_05606_),
    .B1(_02258_),
    .Y(_05607_));
 sky130_fd_sc_hd__a21oi_1 _12433_ (.A1(\div_shifter[63] ),
    .A2(_05606_),
    .B1(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__o21ai_1 _12434_ (.A1(\div_res[30] ),
    .A2(_05572_),
    .B1(net164),
    .Y(_05609_));
 sky130_fd_sc_hd__xnor2_1 _12435_ (.A(\div_res[31] ),
    .B(_05609_),
    .Y(_05611_));
 sky130_fd_sc_hd__o21a_1 _12436_ (.A1(reg1_val[31]),
    .A2(_04687_),
    .B1(_02245_),
    .X(_05612_));
 sky130_fd_sc_hd__a311o_1 _12437_ (.A1(reg1_val[31]),
    .A2(_04687_),
    .A3(_02255_),
    .B1(_05612_),
    .C1(_06459_),
    .X(_05613_));
 sky130_fd_sc_hd__a221o_1 _12438_ (.A1(_04698_),
    .A2(_02249_),
    .B1(_02273_),
    .B2(_02243_),
    .C1(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__a211o_1 _12439_ (.A1(net191),
    .A2(_02238_),
    .B1(_05608_),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__a21o_1 _12440_ (.A1(_02260_),
    .A2(_05611_),
    .B1(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__a211o_1 _12441_ (.A1(_06446_),
    .A2(_05605_),
    .B1(_05616_),
    .C1(_05603_),
    .X(_05617_));
 sky130_fd_sc_hd__o21bai_1 _12442_ (.A1(_05598_),
    .A2(_05600_),
    .B1_N(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__o221a_4 _12443_ (.A1(_04687_),
    .A2(_06460_),
    .B1(_05595_),
    .B2(_05618_),
    .C1(net266),
    .X(dest_val[31]));
 sky130_fd_sc_hd__mux2_1 _12444_ (.A0(net308),
    .A1(curr_PC[0]),
    .S(net263),
    .X(_05619_));
 sky130_fd_sc_hd__nand2_1 _12445_ (.A(_04600_),
    .B(_05619_),
    .Y(_05621_));
 sky130_fd_sc_hd__or2_1 _12446_ (.A(_04600_),
    .B(_05619_),
    .X(_05622_));
 sky130_fd_sc_hd__and2_4 _12447_ (.A(_05621_),
    .B(_05622_),
    .X(new_PC[0]));
 sky130_fd_sc_hd__mux2_1 _12448_ (.A0(net307),
    .A1(curr_PC[1]),
    .S(net263),
    .X(_05623_));
 sky130_fd_sc_hd__nand2_1 _12449_ (.A(_05781_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__or2_1 _12450_ (.A(_05781_),
    .B(_05623_),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _12451_ (.A(_05624_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__or2_1 _12452_ (.A(_05621_),
    .B(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _12453_ (.A(_05621_),
    .B(_05626_),
    .Y(_05628_));
 sky130_fd_sc_hd__and2_4 _12454_ (.A(_05627_),
    .B(_05628_),
    .X(new_PC[1]));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(reg1_val[2]),
    .A1(curr_PC[2]),
    .S(net266),
    .X(_05630_));
 sky130_fd_sc_hd__nand2_1 _12456_ (.A(_05716_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__or2_1 _12457_ (.A(_05716_),
    .B(_05630_),
    .X(_05632_));
 sky130_fd_sc_hd__nand2_1 _12458_ (.A(_05631_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__a21o_1 _12459_ (.A1(_05624_),
    .A2(_05627_),
    .B1(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__nand3_1 _12460_ (.A(_05624_),
    .B(_05627_),
    .C(_05633_),
    .Y(_05635_));
 sky130_fd_sc_hd__and2_4 _12461_ (.A(_05634_),
    .B(_05635_),
    .X(new_PC[2]));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(reg1_val[3]),
    .A1(curr_PC[3]),
    .S(net264),
    .X(_05636_));
 sky130_fd_sc_hd__nand2_1 _12463_ (.A(_05629_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__or2_1 _12464_ (.A(_05629_),
    .B(_05636_),
    .X(_05638_));
 sky130_fd_sc_hd__nand2_1 _12465_ (.A(_05637_),
    .B(_05638_),
    .Y(_05640_));
 sky130_fd_sc_hd__a21o_1 _12466_ (.A1(_05631_),
    .A2(_05634_),
    .B1(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__nand3_1 _12467_ (.A(_05631_),
    .B(_05634_),
    .C(_05640_),
    .Y(_05642_));
 sky130_fd_sc_hd__and2_4 _12468_ (.A(_05641_),
    .B(_05642_),
    .X(new_PC[3]));
 sky130_fd_sc_hd__mux2_1 _12469_ (.A0(reg1_val[4]),
    .A1(curr_PC[4]),
    .S(net264),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_1 _12470_ (.A(_05545_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__or2_1 _12471_ (.A(_05545_),
    .B(_05643_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _12472_ (.A(_05644_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__a21o_1 _12473_ (.A1(_05637_),
    .A2(_05641_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand3_1 _12474_ (.A(_05637_),
    .B(_05641_),
    .C(_05646_),
    .Y(_05648_));
 sky130_fd_sc_hd__and2_4 _12475_ (.A(_05647_),
    .B(_05648_),
    .X(new_PC[4]));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(reg1_val[5]),
    .A1(curr_PC[5]),
    .S(net264),
    .X(_05650_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(_05394_),
    .B(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__or2_1 _12478_ (.A(_05394_),
    .B(_05650_),
    .X(_05652_));
 sky130_fd_sc_hd__nand2_1 _12479_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21o_1 _12480_ (.A1(_05644_),
    .A2(_05647_),
    .B1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__nand3_1 _12481_ (.A(_05644_),
    .B(_05647_),
    .C(_05653_),
    .Y(_05655_));
 sky130_fd_sc_hd__and2_4 _12482_ (.A(_05654_),
    .B(_05655_),
    .X(new_PC[5]));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(reg1_val[6]),
    .A1(curr_PC[6]),
    .S(net264),
    .X(_05656_));
 sky130_fd_sc_hd__nand2_1 _12484_ (.A(_05470_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__or2_1 _12485_ (.A(_05470_),
    .B(_05656_),
    .X(_05659_));
 sky130_fd_sc_hd__nand2_1 _12486_ (.A(_05657_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__a21o_1 _12487_ (.A1(_05651_),
    .A2(_05654_),
    .B1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__nand3_1 _12488_ (.A(_05651_),
    .B(_05654_),
    .C(_05660_),
    .Y(_05662_));
 sky130_fd_sc_hd__and2_4 _12489_ (.A(_05661_),
    .B(_05662_),
    .X(new_PC[6]));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(reg1_val[7]),
    .A1(curr_PC[7]),
    .S(net264),
    .X(_05663_));
 sky130_fd_sc_hd__nand2_1 _12491_ (.A(_05318_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__or2_1 _12492_ (.A(_05318_),
    .B(_05663_),
    .X(_05665_));
 sky130_fd_sc_hd__nand2_1 _12493_ (.A(_05664_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__a21o_1 _12494_ (.A1(_05657_),
    .A2(_05661_),
    .B1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__nand3_1 _12495_ (.A(_05657_),
    .B(_05661_),
    .C(_05666_),
    .Y(_05669_));
 sky130_fd_sc_hd__and2_4 _12496_ (.A(_05667_),
    .B(_05669_),
    .X(new_PC[7]));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(reg1_val[8]),
    .A1(curr_PC[8]),
    .S(net264),
    .X(_05670_));
 sky130_fd_sc_hd__nand2_1 _12498_ (.A(_05253_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__or2_1 _12499_ (.A(_05253_),
    .B(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_05671_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21o_1 _12501_ (.A1(_05664_),
    .A2(_05667_),
    .B1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__nand3_1 _12502_ (.A(_05664_),
    .B(_05667_),
    .C(_05673_),
    .Y(_05675_));
 sky130_fd_sc_hd__and2_4 _12503_ (.A(_05674_),
    .B(_05675_),
    .X(new_PC[8]));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(reg1_val[9]),
    .A1(curr_PC[9]),
    .S(net264),
    .X(_05676_));
 sky130_fd_sc_hd__nand2_1 _12505_ (.A(_05144_),
    .B(_05676_),
    .Y(_05678_));
 sky130_fd_sc_hd__or2_1 _12506_ (.A(_05144_),
    .B(_05676_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(_05678_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__a21o_1 _12508_ (.A1(_05671_),
    .A2(_05674_),
    .B1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__nand3_1 _12509_ (.A(_05671_),
    .B(_05674_),
    .C(_05680_),
    .Y(_05682_));
 sky130_fd_sc_hd__and2_4 _12510_ (.A(_05681_),
    .B(_05682_),
    .X(new_PC[9]));
 sky130_fd_sc_hd__mux2_1 _12511_ (.A0(reg1_val[10]),
    .A1(curr_PC[10]),
    .S(net265),
    .X(_05683_));
 sky130_fd_sc_hd__nand2_1 _12512_ (.A(_05014_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__or2_1 _12513_ (.A(_05014_),
    .B(_05683_),
    .X(_05685_));
 sky130_fd_sc_hd__nand2_1 _12514_ (.A(_05684_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__a21o_1 _12515_ (.A1(_05678_),
    .A2(_05681_),
    .B1(_05686_),
    .X(_05688_));
 sky130_fd_sc_hd__nand3_1 _12516_ (.A(_05678_),
    .B(_05681_),
    .C(_05686_),
    .Y(_05689_));
 sky130_fd_sc_hd__and2_4 _12517_ (.A(_05688_),
    .B(_05689_),
    .X(new_PC[10]));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(reg1_val[11]),
    .A1(curr_PC[11]),
    .S(net264),
    .X(_05690_));
 sky130_fd_sc_hd__nand2_1 _12519_ (.A(_05079_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__or2_1 _12520_ (.A(_05079_),
    .B(_05690_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _12521_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__a21o_1 _12522_ (.A1(_05684_),
    .A2(_05688_),
    .B1(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__nand3_1 _12523_ (.A(_05684_),
    .B(_05688_),
    .C(_05693_),
    .Y(_05695_));
 sky130_fd_sc_hd__and2_4 _12524_ (.A(_05694_),
    .B(_05695_),
    .X(new_PC[11]));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(reg1_val[12]),
    .A1(curr_PC[12]),
    .S(net265),
    .X(_05697_));
 sky130_fd_sc_hd__nand2_1 _12526_ (.A(_04709_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__or2_1 _12527_ (.A(_04709_),
    .B(_05697_),
    .X(_05699_));
 sky130_fd_sc_hd__nand2_1 _12528_ (.A(_05698_),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a21o_1 _12529_ (.A1(_05691_),
    .A2(_05694_),
    .B1(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__nand3_1 _12530_ (.A(_05691_),
    .B(_05694_),
    .C(_05700_),
    .Y(_05702_));
 sky130_fd_sc_hd__and2_4 _12531_ (.A(_05701_),
    .B(_05702_),
    .X(new_PC[12]));
 sky130_fd_sc_hd__mux2_1 _12532_ (.A0(reg1_val[13]),
    .A1(curr_PC[13]),
    .S(net265),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_1 _12533_ (.A(_04948_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__or2_1 _12534_ (.A(_04948_),
    .B(_05703_),
    .X(_05705_));
 sky130_fd_sc_hd__nand2_1 _12535_ (.A(_05704_),
    .B(_05705_),
    .Y(_05707_));
 sky130_fd_sc_hd__a21o_1 _12536_ (.A1(_05698_),
    .A2(_05701_),
    .B1(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__nand3_1 _12537_ (.A(_05698_),
    .B(_05701_),
    .C(_05707_),
    .Y(_05709_));
 sky130_fd_sc_hd__and2_4 _12538_ (.A(_05708_),
    .B(_05709_),
    .X(new_PC[13]));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(reg1_val[14]),
    .A1(curr_PC[14]),
    .S(net264),
    .X(_05710_));
 sky130_fd_sc_hd__nand2_1 _12540_ (.A(_04861_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__or2_1 _12541_ (.A(_04861_),
    .B(_05710_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _12542_ (.A(_05711_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__a21o_1 _12543_ (.A1(_05704_),
    .A2(_05708_),
    .B1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__nand3_1 _12544_ (.A(_05704_),
    .B(_05708_),
    .C(_05713_),
    .Y(_05715_));
 sky130_fd_sc_hd__and2_4 _12545_ (.A(_05714_),
    .B(_05715_),
    .X(new_PC[14]));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(reg1_val[15]),
    .A1(curr_PC[15]),
    .S(net265),
    .X(_05717_));
 sky130_fd_sc_hd__nand2_1 _12547_ (.A(_04785_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__or2_1 _12548_ (.A(_04785_),
    .B(_05717_),
    .X(_05719_));
 sky130_fd_sc_hd__nand2_1 _12549_ (.A(_05718_),
    .B(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__a21o_1 _12550_ (.A1(_05711_),
    .A2(_05714_),
    .B1(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__nand3_1 _12551_ (.A(_05711_),
    .B(_05714_),
    .C(_05720_),
    .Y(_05722_));
 sky130_fd_sc_hd__and2_4 _12552_ (.A(_05721_),
    .B(_05722_),
    .X(new_PC[15]));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(reg1_val[16]),
    .A1(curr_PC[16]),
    .S(net264),
    .X(_05723_));
 sky130_fd_sc_hd__xnor2_1 _12554_ (.A(net283),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__a21o_1 _12555_ (.A1(_05718_),
    .A2(_05721_),
    .B1(_05724_),
    .X(_05726_));
 sky130_fd_sc_hd__nand3_1 _12556_ (.A(_05718_),
    .B(_05721_),
    .C(_05724_),
    .Y(_05727_));
 sky130_fd_sc_hd__and2_4 _12557_ (.A(_05726_),
    .B(_05727_),
    .X(new_PC[16]));
 sky130_fd_sc_hd__mux2_2 _12558_ (.A0(reg1_val[17]),
    .A1(curr_PC[17]),
    .S(net265),
    .X(_05728_));
 sky130_fd_sc_hd__xnor2_4 _12559_ (.A(net283),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__a21bo_1 _12560_ (.A1(net283),
    .A2(_05723_),
    .B1_N(_05726_),
    .X(_05730_));
 sky130_fd_sc_hd__xnor2_4 _12561_ (.A(_05729_),
    .B(_05730_),
    .Y(new_PC[17]));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(reg1_val[18]),
    .A1(curr_PC[18]),
    .S(net265),
    .X(_05731_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(net283),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__or2_1 _12564_ (.A(net283),
    .B(_05731_),
    .X(_05733_));
 sky130_fd_sc_hd__nand2_1 _12565_ (.A(_05732_),
    .B(_05733_),
    .Y(_05735_));
 sky130_fd_sc_hd__or2_1 _12566_ (.A(_05726_),
    .B(_05729_),
    .X(_05736_));
 sky130_fd_sc_hd__o21ai_1 _12567_ (.A1(_05723_),
    .A2(_05728_),
    .B1(net283),
    .Y(_05737_));
 sky130_fd_sc_hd__a21o_1 _12568_ (.A1(_05736_),
    .A2(_05737_),
    .B1(_05735_),
    .X(_05738_));
 sky130_fd_sc_hd__nand3_1 _12569_ (.A(_05735_),
    .B(_05736_),
    .C(_05737_),
    .Y(_05739_));
 sky130_fd_sc_hd__and2_4 _12570_ (.A(_05738_),
    .B(_05739_),
    .X(new_PC[18]));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(reg1_val[19]),
    .A1(curr_PC[19]),
    .S(net265),
    .X(_05740_));
 sky130_fd_sc_hd__nand2_1 _12572_ (.A(net283),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__or2_1 _12573_ (.A(net283),
    .B(_05740_),
    .X(_05742_));
 sky130_fd_sc_hd__nand2_2 _12574_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_2 _12575_ (.A(_05732_),
    .B(_05738_),
    .Y(_05745_));
 sky130_fd_sc_hd__xnor2_4 _12576_ (.A(_05743_),
    .B(_05745_),
    .Y(new_PC[19]));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(reg1_val[20]),
    .A1(curr_PC[20]),
    .S(net265),
    .X(_05746_));
 sky130_fd_sc_hd__nand2_1 _12578_ (.A(net284),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__or2_1 _12579_ (.A(net284),
    .B(_05746_),
    .X(_05748_));
 sky130_fd_sc_hd__nand2_2 _12580_ (.A(_05747_),
    .B(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__or3_1 _12581_ (.A(_05735_),
    .B(_05736_),
    .C(_05743_),
    .X(_05750_));
 sky130_fd_sc_hd__and3_1 _12582_ (.A(_05732_),
    .B(_05737_),
    .C(_05741_),
    .X(_05751_));
 sky130_fd_sc_hd__nand2_2 _12583_ (.A(_05750_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__inv_2 _12584_ (.A(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__xnor2_4 _12585_ (.A(_05749_),
    .B(_05752_),
    .Y(new_PC[20]));
 sky130_fd_sc_hd__mux2_2 _12586_ (.A0(reg1_val[21]),
    .A1(curr_PC[21]),
    .S(net265),
    .X(_05755_));
 sky130_fd_sc_hd__xnor2_4 _12587_ (.A(net284),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21ai_2 _12588_ (.A1(_05749_),
    .A2(_05753_),
    .B1(_05747_),
    .Y(_05757_));
 sky130_fd_sc_hd__xnor2_4 _12589_ (.A(_05756_),
    .B(_05757_),
    .Y(new_PC[21]));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(reg1_val[22]),
    .A1(curr_PC[22]),
    .S(net264),
    .X(_05758_));
 sky130_fd_sc_hd__and2_1 _12591_ (.A(net283),
    .B(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__or2_1 _12592_ (.A(net283),
    .B(_05758_),
    .X(_05760_));
 sky130_fd_sc_hd__nand2b_2 _12593_ (.A_N(_05759_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_2 _12594_ (.A1(_05746_),
    .A2(_05755_),
    .B1(net284),
    .Y(_05762_));
 sky130_fd_sc_hd__nor2_1 _12595_ (.A(_05749_),
    .B(_05756_),
    .Y(_05764_));
 sky130_fd_sc_hd__inv_2 _12596_ (.A(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__o21ai_4 _12597_ (.A1(_05753_),
    .A2(_05765_),
    .B1(_05762_),
    .Y(_05766_));
 sky130_fd_sc_hd__xnor2_4 _12598_ (.A(_05761_),
    .B(_05766_),
    .Y(new_PC[22]));
 sky130_fd_sc_hd__mux2_2 _12599_ (.A0(reg1_val[23]),
    .A1(curr_PC[23]),
    .S(net264),
    .X(_05767_));
 sky130_fd_sc_hd__xnor2_4 _12600_ (.A(net283),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__a21o_1 _12601_ (.A1(_05760_),
    .A2(_05766_),
    .B1(_05759_),
    .X(_05769_));
 sky130_fd_sc_hd__xnor2_4 _12602_ (.A(_05768_),
    .B(_05769_),
    .Y(new_PC[23]));
 sky130_fd_sc_hd__mux2_2 _12603_ (.A0(reg1_val[24]),
    .A1(curr_PC[24]),
    .S(net264),
    .X(_05770_));
 sky130_fd_sc_hd__xnor2_4 _12604_ (.A(net283),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__or4_1 _12605_ (.A(_05750_),
    .B(_05761_),
    .C(_05765_),
    .D(_05768_),
    .X(_05773_));
 sky130_fd_sc_hd__o21ai_1 _12606_ (.A1(_05758_),
    .A2(_05767_),
    .B1(net283),
    .Y(_05774_));
 sky130_fd_sc_hd__and4_2 _12607_ (.A(_05751_),
    .B(_05762_),
    .C(_05773_),
    .D(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__xor2_4 _12608_ (.A(_05771_),
    .B(_05775_),
    .X(new_PC[24]));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(reg1_val[25]),
    .A1(curr_PC[25]),
    .S(net264),
    .X(_05776_));
 sky130_fd_sc_hd__and2_1 _12610_ (.A(net284),
    .B(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__nor2_1 _12611_ (.A(net284),
    .B(_05776_),
    .Y(_05778_));
 sky130_fd_sc_hd__nor2_2 _12612_ (.A(_05777_),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__o2bb2a_2 _12613_ (.A1_N(net284),
    .A2_N(_05770_),
    .B1(_05771_),
    .B2(_05775_),
    .X(_05780_));
 sky130_fd_sc_hd__xnor2_4 _12614_ (.A(_05779_),
    .B(_05780_),
    .Y(new_PC[25]));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(reg1_val[26]),
    .A1(curr_PC[26]),
    .S(net264),
    .X(_05782_));
 sky130_fd_sc_hd__and2_1 _12616_ (.A(net283),
    .B(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__nor2_1 _12617_ (.A(net283),
    .B(_05782_),
    .Y(_05784_));
 sky130_fd_sc_hd__nor2_2 _12618_ (.A(_05783_),
    .B(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__o21ba_2 _12619_ (.A1(_05778_),
    .A2(_05780_),
    .B1_N(_05777_),
    .X(_05786_));
 sky130_fd_sc_hd__xnor2_4 _12620_ (.A(_05785_),
    .B(_05786_),
    .Y(new_PC[26]));
 sky130_fd_sc_hd__o21ba_2 _12621_ (.A1(_05784_),
    .A2(_05786_),
    .B1_N(_05783_),
    .X(_05787_));
 sky130_fd_sc_hd__mux2_1 _12622_ (.A0(reg1_val[27]),
    .A1(curr_PC[27]),
    .S(net264),
    .X(_05788_));
 sky130_fd_sc_hd__xor2_2 _12623_ (.A(net283),
    .B(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__xnor2_4 _12624_ (.A(_05787_),
    .B(_05789_),
    .Y(new_PC[27]));
 sky130_fd_sc_hd__nand2_2 _12625_ (.A(net308),
    .B(_04600_),
    .Y(_05791_));
 sky130_fd_sc_hd__or2_1 _12626_ (.A(net308),
    .B(_04600_),
    .X(_05792_));
 sky130_fd_sc_hd__and2_4 _12627_ (.A(_05791_),
    .B(_05792_),
    .X(loadstore_address[0]));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(reg1_val[1]),
    .B(_05781_),
    .Y(_05793_));
 sky130_fd_sc_hd__or2_1 _12629_ (.A(reg1_val[1]),
    .B(_05781_),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_2 _12630_ (.A(_05793_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__xor2_4 _12631_ (.A(_05791_),
    .B(_05795_),
    .X(loadstore_address[1]));
 sky130_fd_sc_hd__o21a_2 _12632_ (.A1(_05791_),
    .A2(_05795_),
    .B1(_05793_),
    .X(_05796_));
 sky130_fd_sc_hd__nor2_1 _12633_ (.A(reg1_val[2]),
    .B(_05716_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_1 _12634_ (.A(reg1_val[2]),
    .B(_05716_),
    .Y(_05798_));
 sky130_fd_sc_hd__and2b_2 _12635_ (.A_N(_05797_),
    .B(_05798_),
    .X(_05800_));
 sky130_fd_sc_hd__xnor2_4 _12636_ (.A(_05796_),
    .B(_05800_),
    .Y(loadstore_address[2]));
 sky130_fd_sc_hd__o21a_2 _12637_ (.A1(_05796_),
    .A2(_05797_),
    .B1(_05798_),
    .X(_05801_));
 sky130_fd_sc_hd__nor2_1 _12638_ (.A(reg1_val[3]),
    .B(_05629_),
    .Y(_05802_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(reg1_val[3]),
    .B(_05629_),
    .Y(_05803_));
 sky130_fd_sc_hd__and2b_2 _12640_ (.A_N(_05802_),
    .B(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__xnor2_4 _12641_ (.A(_05801_),
    .B(_05804_),
    .Y(loadstore_address[3]));
 sky130_fd_sc_hd__o21a_2 _12642_ (.A1(_05801_),
    .A2(_05802_),
    .B1(_05803_),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _12643_ (.A(reg1_val[4]),
    .B(_05545_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _12644_ (.A(reg1_val[4]),
    .B(_05545_),
    .Y(_05807_));
 sky130_fd_sc_hd__and2b_1 _12645_ (.A_N(_05806_),
    .B(_05807_),
    .X(_05809_));
 sky130_fd_sc_hd__xnor2_4 _12646_ (.A(_05805_),
    .B(_05809_),
    .Y(loadstore_address[4]));
 sky130_fd_sc_hd__o21a_2 _12647_ (.A1(_05805_),
    .A2(_05806_),
    .B1(_05807_),
    .X(_05810_));
 sky130_fd_sc_hd__nor2_1 _12648_ (.A(reg1_val[5]),
    .B(_05394_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand2_1 _12649_ (.A(reg1_val[5]),
    .B(_05394_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand2b_2 _12650_ (.A_N(_05811_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__xor2_4 _12651_ (.A(_05810_),
    .B(_05813_),
    .X(loadstore_address[5]));
 sky130_fd_sc_hd__o21a_2 _12652_ (.A1(_05810_),
    .A2(_05811_),
    .B1(_05812_),
    .X(_05814_));
 sky130_fd_sc_hd__nor2_1 _12653_ (.A(reg1_val[6]),
    .B(_05470_),
    .Y(_05815_));
 sky130_fd_sc_hd__and2_1 _12654_ (.A(reg1_val[6]),
    .B(_05470_),
    .X(_05816_));
 sky130_fd_sc_hd__or2_2 _12655_ (.A(_05815_),
    .B(_05816_),
    .X(_05818_));
 sky130_fd_sc_hd__xor2_4 _12656_ (.A(_05814_),
    .B(_05818_),
    .X(loadstore_address[6]));
 sky130_fd_sc_hd__o21ba_2 _12657_ (.A1(_05814_),
    .A2(_05815_),
    .B1_N(_05816_),
    .X(_05819_));
 sky130_fd_sc_hd__nor2_1 _12658_ (.A(reg1_val[7]),
    .B(_05318_),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_1 _12659_ (.A(reg1_val[7]),
    .B(_05318_),
    .Y(_05821_));
 sky130_fd_sc_hd__nand2b_2 _12660_ (.A_N(_05820_),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__xor2_4 _12661_ (.A(_05819_),
    .B(_05822_),
    .X(loadstore_address[7]));
 sky130_fd_sc_hd__o21a_2 _12662_ (.A1(_05819_),
    .A2(_05820_),
    .B1(_05821_),
    .X(_05823_));
 sky130_fd_sc_hd__nor2_1 _12663_ (.A(reg1_val[8]),
    .B(_05253_),
    .Y(_05824_));
 sky130_fd_sc_hd__nand2_1 _12664_ (.A(reg1_val[8]),
    .B(_05253_),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2b_2 _12665_ (.A_N(_05824_),
    .B(_05825_),
    .Y(_05827_));
 sky130_fd_sc_hd__xor2_4 _12666_ (.A(_05823_),
    .B(_05827_),
    .X(loadstore_address[8]));
 sky130_fd_sc_hd__o21a_2 _12667_ (.A1(_05823_),
    .A2(_05824_),
    .B1(_05825_),
    .X(_05828_));
 sky130_fd_sc_hd__or2_1 _12668_ (.A(reg1_val[9]),
    .B(_05144_),
    .X(_05829_));
 sky130_fd_sc_hd__nand2_1 _12669_ (.A(reg1_val[9]),
    .B(_05144_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_2 _12670_ (.A(_05829_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__xor2_4 _12671_ (.A(_05828_),
    .B(_05831_),
    .X(loadstore_address[9]));
 sky130_fd_sc_hd__or2_1 _12672_ (.A(reg1_val[10]),
    .B(_05014_),
    .X(_05832_));
 sky130_fd_sc_hd__nand2_1 _12673_ (.A(reg1_val[10]),
    .B(_05014_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _12674_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2b_1 _12675_ (.A_N(_05828_),
    .B(_05829_),
    .Y(_05836_));
 sky130_fd_sc_hd__a21o_1 _12676_ (.A1(_05830_),
    .A2(_05836_),
    .B1(_05834_),
    .X(_05837_));
 sky130_fd_sc_hd__nand3_1 _12677_ (.A(_05830_),
    .B(_05834_),
    .C(_05836_),
    .Y(_05838_));
 sky130_fd_sc_hd__and2_4 _12678_ (.A(_05837_),
    .B(_05838_),
    .X(loadstore_address[10]));
 sky130_fd_sc_hd__or2_1 _12679_ (.A(reg1_val[11]),
    .B(_05079_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_1 _12680_ (.A(reg1_val[11]),
    .B(_05079_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _12681_ (.A(_05839_),
    .B(_05840_),
    .Y(_05841_));
 sky130_fd_sc_hd__a21o_1 _12682_ (.A1(_05833_),
    .A2(_05837_),
    .B1(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__nand3_1 _12683_ (.A(_05833_),
    .B(_05837_),
    .C(_05841_),
    .Y(_05843_));
 sky130_fd_sc_hd__and2_4 _12684_ (.A(_05842_),
    .B(_05843_),
    .X(loadstore_address[11]));
 sky130_fd_sc_hd__or2_1 _12685_ (.A(reg1_val[12]),
    .B(_04709_),
    .X(_05845_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(reg1_val[12]),
    .B(_04709_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _12687_ (.A(_05845_),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__a21o_1 _12688_ (.A1(_05840_),
    .A2(_05842_),
    .B1(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__nand3_1 _12689_ (.A(_05840_),
    .B(_05842_),
    .C(_05847_),
    .Y(_05849_));
 sky130_fd_sc_hd__and2_4 _12690_ (.A(_05848_),
    .B(_05849_),
    .X(loadstore_address[12]));
 sky130_fd_sc_hd__or2_1 _12691_ (.A(reg1_val[13]),
    .B(_04948_),
    .X(_05850_));
 sky130_fd_sc_hd__nand2_1 _12692_ (.A(reg1_val[13]),
    .B(_04948_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_1 _12693_ (.A(_05850_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__a21o_1 _12694_ (.A1(_05846_),
    .A2(_05848_),
    .B1(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__nand3_1 _12695_ (.A(_05846_),
    .B(_05848_),
    .C(_05852_),
    .Y(_05855_));
 sky130_fd_sc_hd__and2_4 _12696_ (.A(_05853_),
    .B(_05855_),
    .X(loadstore_address[13]));
 sky130_fd_sc_hd__or2_1 _12697_ (.A(reg1_val[14]),
    .B(_04861_),
    .X(_05856_));
 sky130_fd_sc_hd__nand2_1 _12698_ (.A(reg1_val[14]),
    .B(_04861_),
    .Y(_05857_));
 sky130_fd_sc_hd__nand2_1 _12699_ (.A(_05856_),
    .B(_05857_),
    .Y(_05858_));
 sky130_fd_sc_hd__a21o_1 _12700_ (.A1(_05851_),
    .A2(_05853_),
    .B1(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__nand3_1 _12701_ (.A(_05851_),
    .B(_05853_),
    .C(_05858_),
    .Y(_05860_));
 sky130_fd_sc_hd__and2_4 _12702_ (.A(_05859_),
    .B(_05860_),
    .X(loadstore_address[14]));
 sky130_fd_sc_hd__xnor2_2 _12703_ (.A(reg1_val[15]),
    .B(_04785_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21oi_4 _12704_ (.A1(_05857_),
    .A2(_05859_),
    .B1(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__and3_2 _12705_ (.A(_05857_),
    .B(_05859_),
    .C(_05861_),
    .X(_05864_));
 sky130_fd_sc_hd__nor2_8 _12706_ (.A(_05862_),
    .B(_05864_),
    .Y(loadstore_address[15]));
 sky130_fd_sc_hd__nor2_1 _12707_ (.A(reg1_val[16]),
    .B(net285),
    .Y(_05865_));
 sky130_fd_sc_hd__and2_1 _12708_ (.A(reg1_val[16]),
    .B(net285),
    .X(_05866_));
 sky130_fd_sc_hd__or2_2 _12709_ (.A(_05865_),
    .B(_05866_),
    .X(_05867_));
 sky130_fd_sc_hd__a21oi_4 _12710_ (.A1(reg1_val[15]),
    .A2(_04785_),
    .B1(_05862_),
    .Y(_05868_));
 sky130_fd_sc_hd__or2_1 _12711_ (.A(_05867_),
    .B(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__xor2_4 _12712_ (.A(_05867_),
    .B(_05868_),
    .X(loadstore_address[16]));
 sky130_fd_sc_hd__nand2b_2 _12713_ (.A_N(_05866_),
    .B(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__xnor2_4 _12714_ (.A(reg1_val[17]),
    .B(net285),
    .Y(_05871_));
 sky130_fd_sc_hd__xnor2_4 _12715_ (.A(_05870_),
    .B(_05871_),
    .Y(loadstore_address[17]));
 sky130_fd_sc_hd__or2_1 _12716_ (.A(reg1_val[18]),
    .B(net285),
    .X(_05873_));
 sky130_fd_sc_hd__nand2_1 _12717_ (.A(reg1_val[18]),
    .B(net285),
    .Y(_05874_));
 sky130_fd_sc_hd__nand2_2 _12718_ (.A(_05873_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__a2bb2o_2 _12719_ (.A1_N(_05869_),
    .A2_N(_05871_),
    .B1(net285),
    .B2(_06517_),
    .X(_05876_));
 sky130_fd_sc_hd__xnor2_4 _12720_ (.A(_05875_),
    .B(_05876_),
    .Y(loadstore_address[18]));
 sky130_fd_sc_hd__a21bo_1 _12721_ (.A1(_05873_),
    .A2(_05876_),
    .B1_N(_05874_),
    .X(_05877_));
 sky130_fd_sc_hd__xnor2_4 _12722_ (.A(reg1_val[19]),
    .B(net285),
    .Y(_05878_));
 sky130_fd_sc_hd__xnor2_4 _12723_ (.A(_05877_),
    .B(_05878_),
    .Y(loadstore_address[19]));
 sky130_fd_sc_hd__xnor2_2 _12724_ (.A(reg1_val[20]),
    .B(net285),
    .Y(_05879_));
 sky130_fd_sc_hd__or4_2 _12725_ (.A(_05869_),
    .B(_05871_),
    .C(_05875_),
    .D(_05878_),
    .X(_05881_));
 sky130_fd_sc_hd__nand2_1 _12726_ (.A(net285),
    .B(_06518_),
    .Y(_05882_));
 sky130_fd_sc_hd__a21oi_4 _12727_ (.A1(_05881_),
    .A2(_05882_),
    .B1(_05879_),
    .Y(_05883_));
 sky130_fd_sc_hd__and3_2 _12728_ (.A(_05879_),
    .B(_05881_),
    .C(_05882_),
    .X(_05884_));
 sky130_fd_sc_hd__nor2_8 _12729_ (.A(_05883_),
    .B(_05884_),
    .Y(loadstore_address[20]));
 sky130_fd_sc_hd__nor2_1 _12730_ (.A(reg1_val[21]),
    .B(net285),
    .Y(_05885_));
 sky130_fd_sc_hd__nand2_2 _12731_ (.A(reg1_val[21]),
    .B(net285),
    .Y(_05886_));
 sky130_fd_sc_hd__nand2b_2 _12732_ (.A_N(_05885_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__a21oi_4 _12733_ (.A1(reg1_val[20]),
    .A2(net285),
    .B1(_05883_),
    .Y(_05888_));
 sky130_fd_sc_hd__xor2_4 _12734_ (.A(_05887_),
    .B(_05888_),
    .X(loadstore_address[21]));
 sky130_fd_sc_hd__or2_1 _12735_ (.A(reg1_val[22]),
    .B(net285),
    .X(_05890_));
 sky130_fd_sc_hd__nand2_1 _12736_ (.A(reg1_val[22]),
    .B(net285),
    .Y(_05891_));
 sky130_fd_sc_hd__nand2_2 _12737_ (.A(_05890_),
    .B(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__o21ai_4 _12738_ (.A1(_05885_),
    .A2(_05888_),
    .B1(_05886_),
    .Y(_05893_));
 sky130_fd_sc_hd__xnor2_4 _12739_ (.A(_05892_),
    .B(_05893_),
    .Y(loadstore_address[22]));
 sky130_fd_sc_hd__a21bo_1 _12740_ (.A1(_05890_),
    .A2(_05893_),
    .B1_N(_05891_),
    .X(_05894_));
 sky130_fd_sc_hd__xnor2_4 _12741_ (.A(reg1_val[23]),
    .B(net285),
    .Y(_05895_));
 sky130_fd_sc_hd__xnor2_4 _12742_ (.A(_05894_),
    .B(_05895_),
    .Y(loadstore_address[23]));
 sky130_fd_sc_hd__or2_1 _12743_ (.A(reg1_val[24]),
    .B(net286),
    .X(_05896_));
 sky130_fd_sc_hd__nand2_1 _12744_ (.A(reg1_val[24]),
    .B(net286),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_2 _12745_ (.A(_05896_),
    .B(_05897_),
    .Y(_05899_));
 sky130_fd_sc_hd__or4_1 _12746_ (.A(_05879_),
    .B(_05887_),
    .C(_05892_),
    .D(_05895_),
    .X(_05900_));
 sky130_fd_sc_hd__a2bb2o_2 _12747_ (.A1_N(_05881_),
    .A2_N(_05900_),
    .B1(net285),
    .B2(_06519_),
    .X(_05901_));
 sky130_fd_sc_hd__nand2b_1 _12748_ (.A_N(_05899_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__xnor2_4 _12749_ (.A(_05899_),
    .B(_05901_),
    .Y(loadstore_address[24]));
 sky130_fd_sc_hd__nand2_2 _12750_ (.A(_05897_),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__xnor2_4 _12751_ (.A(reg1_val[25]),
    .B(net286),
    .Y(_05904_));
 sky130_fd_sc_hd__xnor2_4 _12752_ (.A(_05903_),
    .B(_05904_),
    .Y(loadstore_address[25]));
 sky130_fd_sc_hd__xnor2_2 _12753_ (.A(reg1_val[26]),
    .B(net286),
    .Y(_05905_));
 sky130_fd_sc_hd__or2_1 _12754_ (.A(_05902_),
    .B(_05904_),
    .X(_05906_));
 sky130_fd_sc_hd__o21ai_2 _12755_ (.A1(reg1_val[24]),
    .A2(reg1_val[25]),
    .B1(net286),
    .Y(_05908_));
 sky130_fd_sc_hd__a21oi_4 _12756_ (.A1(_05906_),
    .A2(_05908_),
    .B1(_05905_),
    .Y(_05909_));
 sky130_fd_sc_hd__and3_2 _12757_ (.A(_05905_),
    .B(_05906_),
    .C(_05908_),
    .X(_05910_));
 sky130_fd_sc_hd__nor2_8 _12758_ (.A(_05909_),
    .B(_05910_),
    .Y(loadstore_address[26]));
 sky130_fd_sc_hd__a21o_1 _12759_ (.A1(reg1_val[26]),
    .A2(net286),
    .B1(_05909_),
    .X(_05911_));
 sky130_fd_sc_hd__xnor2_4 _12760_ (.A(reg1_val[27]),
    .B(net286),
    .Y(_05912_));
 sky130_fd_sc_hd__xnor2_4 _12761_ (.A(_05911_),
    .B(_05912_),
    .Y(loadstore_address[27]));
 sky130_fd_sc_hd__nor2_1 _12762_ (.A(reg1_val[28]),
    .B(net286),
    .Y(_05913_));
 sky130_fd_sc_hd__and2_1 _12763_ (.A(reg1_val[28]),
    .B(net286),
    .X(_05914_));
 sky130_fd_sc_hd__or2_1 _12764_ (.A(_05913_),
    .B(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__nand2_1 _12765_ (.A(net286),
    .B(_00344_),
    .Y(_05917_));
 sky130_fd_sc_hd__or3_1 _12766_ (.A(_05905_),
    .B(_05906_),
    .C(_05912_),
    .X(_05918_));
 sky130_fd_sc_hd__a21oi_2 _12767_ (.A1(_05917_),
    .A2(_05918_),
    .B1(_05915_),
    .Y(_05919_));
 sky130_fd_sc_hd__and3_2 _12768_ (.A(_05915_),
    .B(_05917_),
    .C(_05918_),
    .X(_05920_));
 sky130_fd_sc_hd__nor2_8 _12769_ (.A(_05919_),
    .B(_05920_),
    .Y(loadstore_address[28]));
 sky130_fd_sc_hd__nand2_1 _12770_ (.A(reg1_val[29]),
    .B(net286),
    .Y(_05921_));
 sky130_fd_sc_hd__or2_1 _12771_ (.A(reg1_val[29]),
    .B(net286),
    .X(_05922_));
 sky130_fd_sc_hd__nand2_2 _12772_ (.A(_05921_),
    .B(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__or2_2 _12773_ (.A(_05914_),
    .B(_05919_),
    .X(_05924_));
 sky130_fd_sc_hd__xnor2_4 _12774_ (.A(_05923_),
    .B(_05924_),
    .Y(loadstore_address[29]));
 sky130_fd_sc_hd__or2_1 _12775_ (.A(reg1_val[30]),
    .B(net286),
    .X(_05926_));
 sky130_fd_sc_hd__nand2_1 _12776_ (.A(reg1_val[30]),
    .B(net286),
    .Y(_05927_));
 sky130_fd_sc_hd__nand2_2 _12777_ (.A(_05926_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__a21bo_2 _12778_ (.A1(_05922_),
    .A2(_05924_),
    .B1_N(_05921_),
    .X(_05929_));
 sky130_fd_sc_hd__xnor2_4 _12779_ (.A(_05928_),
    .B(_05929_),
    .Y(loadstore_address[30]));
 sky130_fd_sc_hd__a21bo_1 _12780_ (.A1(_05926_),
    .A2(_05929_),
    .B1_N(_05927_),
    .X(_05930_));
 sky130_fd_sc_hd__xnor2_2 _12781_ (.A(reg1_val[31]),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__xnor2_4 _12782_ (.A(net286),
    .B(_05931_),
    .Y(loadstore_address[31]));
 sky130_fd_sc_hd__nand2_1 _12783_ (.A(net482),
    .B(net373),
    .Y(_05932_));
 sky130_fd_sc_hd__nand3_1 _12784_ (.A(net476),
    .B(net482),
    .C(net373),
    .Y(_05933_));
 sky130_fd_sc_hd__and4_1 _12785_ (.A(net411),
    .B(net476),
    .C(\div_counter[1] ),
    .D(net373),
    .X(_05935_));
 sky130_fd_sc_hd__inv_2 _12786_ (.A(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand2_1 _12787_ (.A(net363),
    .B(net477),
    .Y(_05937_));
 sky130_fd_sc_hd__nor2_1 _12788_ (.A(net274),
    .B(net478),
    .Y(_05938_));
 sky130_fd_sc_hd__nor3_1 _12789_ (.A(rst),
    .B(net223),
    .C(_05938_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _12790_ (.A(net280),
    .B(_06431_),
    .Y(_05939_));
 sky130_fd_sc_hd__nand2_1 _12791_ (.A(net273),
    .B(_06430_),
    .Y(_05940_));
 sky130_fd_sc_hd__or2_1 _12792_ (.A(net371),
    .B(net200),
    .X(_05941_));
 sky130_fd_sc_hd__o211a_1 _12793_ (.A1(net35),
    .A2(net197),
    .B1(net372),
    .C1(net297),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _12794_ (.A(net229),
    .B(net202),
    .Y(_05942_));
 sky130_fd_sc_hd__o211a_1 _12795_ (.A1(net369),
    .A2(net202),
    .B1(_05942_),
    .C1(net300),
    .X(_00002_));
 sky130_fd_sc_hd__or2_1 _12796_ (.A(net442),
    .B(net202),
    .X(_05944_));
 sky130_fd_sc_hd__o211a_1 _12797_ (.A1(_06526_),
    .A2(net198),
    .B1(net443),
    .C1(net300),
    .X(_00003_));
 sky130_fd_sc_hd__nand2_1 _12798_ (.A(net183),
    .B(net202),
    .Y(_05945_));
 sky130_fd_sc_hd__o211a_1 _12799_ (.A1(net337),
    .A2(net202),
    .B1(_05945_),
    .C1(net299),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _12800_ (.A(net398),
    .B(net201),
    .X(_05946_));
 sky130_fd_sc_hd__o211a_1 _12801_ (.A1(_06565_),
    .A2(net198),
    .B1(net399),
    .C1(net299),
    .X(_00005_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(net144),
    .B(net201),
    .Y(_05947_));
 sky130_fd_sc_hd__o211a_1 _12803_ (.A1(net359),
    .A2(net201),
    .B1(_05947_),
    .C1(net299),
    .X(_00006_));
 sky130_fd_sc_hd__nand2_1 _12804_ (.A(net148),
    .B(net201),
    .Y(_05948_));
 sky130_fd_sc_hd__o211a_1 _12805_ (.A1(net345),
    .A2(net201),
    .B1(_05948_),
    .C1(net299),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _12806_ (.A(net400),
    .B(net201),
    .X(_05950_));
 sky130_fd_sc_hd__o211a_1 _12807_ (.A1(_06556_),
    .A2(net197),
    .B1(net401),
    .C1(net297),
    .X(_00008_));
 sky130_fd_sc_hd__nand2_1 _12808_ (.A(net142),
    .B(net200),
    .Y(_05951_));
 sky130_fd_sc_hd__o211a_1 _12809_ (.A1(net361),
    .A2(net200),
    .B1(_05951_),
    .C1(net297),
    .X(_00009_));
 sky130_fd_sc_hd__nand2_1 _12810_ (.A(net140),
    .B(net200),
    .Y(_05952_));
 sky130_fd_sc_hd__o211a_1 _12811_ (.A1(net365),
    .A2(net200),
    .B1(_05952_),
    .C1(net297),
    .X(_00010_));
 sky130_fd_sc_hd__nand2_1 _12812_ (.A(_00186_),
    .B(net200),
    .Y(_05953_));
 sky130_fd_sc_hd__o211a_1 _12813_ (.A1(net317),
    .A2(net200),
    .B1(_05953_),
    .C1(net297),
    .X(_00011_));
 sky130_fd_sc_hd__nand2_1 _12814_ (.A(_00191_),
    .B(net201),
    .Y(_05954_));
 sky130_fd_sc_hd__o211a_1 _12815_ (.A1(net343),
    .A2(net201),
    .B1(_05954_),
    .C1(net297),
    .X(_00012_));
 sky130_fd_sc_hd__nand2_1 _12816_ (.A(_00158_),
    .B(net201),
    .Y(_05956_));
 sky130_fd_sc_hd__o211a_1 _12817_ (.A1(net347),
    .A2(net201),
    .B1(_05956_),
    .C1(net301),
    .X(_00013_));
 sky130_fd_sc_hd__nand2_1 _12818_ (.A(net97),
    .B(net201),
    .Y(_05957_));
 sky130_fd_sc_hd__o211a_1 _12819_ (.A1(net355),
    .A2(net201),
    .B1(_05957_),
    .C1(net301),
    .X(_00014_));
 sky130_fd_sc_hd__nand2_1 _12820_ (.A(net90),
    .B(net203),
    .Y(_05958_));
 sky130_fd_sc_hd__o211a_1 _12821_ (.A1(net353),
    .A2(net201),
    .B1(_05958_),
    .C1(net301),
    .X(_00015_));
 sky130_fd_sc_hd__nand2_1 _12822_ (.A(_06502_),
    .B(net203),
    .Y(_05959_));
 sky130_fd_sc_hd__o211a_1 _12823_ (.A1(net333),
    .A2(net203),
    .B1(_05959_),
    .C1(net301),
    .X(_00016_));
 sky130_fd_sc_hd__nand2_1 _12824_ (.A(_06509_),
    .B(net203),
    .Y(_05960_));
 sky130_fd_sc_hd__o211a_1 _12825_ (.A1(net323),
    .A2(net201),
    .B1(_05960_),
    .C1(net301),
    .X(_00017_));
 sky130_fd_sc_hd__nand2_1 _12826_ (.A(_06491_),
    .B(net203),
    .Y(_05962_));
 sky130_fd_sc_hd__o211a_1 _12827_ (.A1(net327),
    .A2(net203),
    .B1(_05962_),
    .C1(net301),
    .X(_00018_));
 sky130_fd_sc_hd__nand2_1 _12828_ (.A(_06494_),
    .B(net203),
    .Y(_05963_));
 sky130_fd_sc_hd__o211a_1 _12829_ (.A1(net335),
    .A2(net203),
    .B1(_05963_),
    .C1(net301),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_1 _12830_ (.A(net86),
    .B(net203),
    .Y(_05964_));
 sky130_fd_sc_hd__o211a_1 _12831_ (.A1(net357),
    .A2(net201),
    .B1(_05964_),
    .C1(net298),
    .X(_00020_));
 sky130_fd_sc_hd__nand2_1 _12832_ (.A(net81),
    .B(net200),
    .Y(_05965_));
 sky130_fd_sc_hd__o211a_1 _12833_ (.A1(net331),
    .A2(net200),
    .B1(_05965_),
    .C1(net298),
    .X(_00021_));
 sky130_fd_sc_hd__nand2_1 _12834_ (.A(net43),
    .B(net199),
    .Y(_05966_));
 sky130_fd_sc_hd__o211a_1 _12835_ (.A1(net325),
    .A2(net199),
    .B1(_05966_),
    .C1(net295),
    .X(_00022_));
 sky130_fd_sc_hd__nand2_1 _12836_ (.A(net40),
    .B(net199),
    .Y(_05968_));
 sky130_fd_sc_hd__o211a_1 _12837_ (.A1(net319),
    .A2(net199),
    .B1(_05968_),
    .C1(net296),
    .X(_00023_));
 sky130_fd_sc_hd__nand2_1 _12838_ (.A(net49),
    .B(net199),
    .Y(_05969_));
 sky130_fd_sc_hd__o211a_1 _12839_ (.A1(net313),
    .A2(net199),
    .B1(_05969_),
    .C1(net295),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _12840_ (.A(net46),
    .B(net199),
    .Y(_05970_));
 sky130_fd_sc_hd__o211a_1 _12841_ (.A1(net311),
    .A2(net199),
    .B1(_05970_),
    .C1(net296),
    .X(_00025_));
 sky130_fd_sc_hd__nand2_1 _12842_ (.A(net55),
    .B(net199),
    .Y(_05971_));
 sky130_fd_sc_hd__o211a_1 _12843_ (.A1(net329),
    .A2(net199),
    .B1(_05971_),
    .C1(net295),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _12844_ (.A(net52),
    .B(net199),
    .Y(_05972_));
 sky130_fd_sc_hd__o211a_1 _12845_ (.A1(net351),
    .A2(net199),
    .B1(_05972_),
    .C1(net296),
    .X(_00027_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(net63),
    .B(net199),
    .Y(_05974_));
 sky130_fd_sc_hd__o211a_1 _12847_ (.A1(net339),
    .A2(net199),
    .B1(_05974_),
    .C1(net296),
    .X(_00028_));
 sky130_fd_sc_hd__nand2_1 _12848_ (.A(net60),
    .B(net199),
    .Y(_05975_));
 sky130_fd_sc_hd__o211a_1 _12849_ (.A1(net349),
    .A2(net199),
    .B1(_05975_),
    .C1(net298),
    .X(_00029_));
 sky130_fd_sc_hd__or2_1 _12850_ (.A(net450),
    .B(net200),
    .X(_05976_));
 sky130_fd_sc_hd__o211a_1 _12851_ (.A1(_00242_),
    .A2(net197),
    .B1(net451),
    .C1(net297),
    .X(_00030_));
 sky130_fd_sc_hd__nand2_1 _12852_ (.A(net19),
    .B(net200),
    .Y(_05977_));
 sky130_fd_sc_hd__o211a_1 _12853_ (.A1(net341),
    .A2(net200),
    .B1(_05977_),
    .C1(net297),
    .X(_00031_));
 sky130_fd_sc_hd__nand2_1 _12854_ (.A(net14),
    .B(net200),
    .Y(_05978_));
 sky130_fd_sc_hd__o211a_1 _12855_ (.A1(net321),
    .A2(net200),
    .B1(_05978_),
    .C1(net298),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _12856_ (.A(net396),
    .B(net200),
    .X(_05980_));
 sky130_fd_sc_hd__o211a_1 _12857_ (.A1(_00510_),
    .A2(net197),
    .B1(net397),
    .C1(net298),
    .X(_00033_));
 sky130_fd_sc_hd__and2b_1 _12858_ (.A_N(net321),
    .B(\div_shifter[61] ),
    .X(_05981_));
 sky130_fd_sc_hd__and2b_1 _12859_ (.A_N(\div_shifter[61] ),
    .B(net321),
    .X(_05982_));
 sky130_fd_sc_hd__nor2_1 _12860_ (.A(_05981_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__and2b_1 _12861_ (.A_N(net341),
    .B(net576),
    .X(_05984_));
 sky130_fd_sc_hd__nand2b_1 _12862_ (.A_N(net576),
    .B(net341),
    .Y(_05985_));
 sky130_fd_sc_hd__and2b_1 _12863_ (.A_N(net450),
    .B(net566),
    .X(_05986_));
 sky130_fd_sc_hd__and2b_1 _12864_ (.A_N(net349),
    .B(\div_shifter[58] ),
    .X(_05987_));
 sky130_fd_sc_hd__nand2b_1 _12865_ (.A_N(\div_shifter[58] ),
    .B(net349),
    .Y(_05989_));
 sky130_fd_sc_hd__and2b_1 _12866_ (.A_N(net339),
    .B(net571),
    .X(_05990_));
 sky130_fd_sc_hd__nand2b_1 _12867_ (.A_N(net571),
    .B(net339),
    .Y(_05991_));
 sky130_fd_sc_hd__nand2b_1 _12868_ (.A_N(_05990_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__and2b_1 _12869_ (.A_N(net351),
    .B(net564),
    .X(_05993_));
 sky130_fd_sc_hd__nand2b_1 _12870_ (.A_N(net564),
    .B(net351),
    .Y(_05994_));
 sky130_fd_sc_hd__and2b_1 _12871_ (.A_N(net329),
    .B(\div_shifter[55] ),
    .X(_05995_));
 sky130_fd_sc_hd__and2b_1 _12872_ (.A_N(net311),
    .B(net556),
    .X(_05996_));
 sky130_fd_sc_hd__nand2b_1 _12873_ (.A_N(net556),
    .B(net311),
    .Y(_05997_));
 sky130_fd_sc_hd__and2b_1 _12874_ (.A_N(net313),
    .B(net562),
    .X(_05998_));
 sky130_fd_sc_hd__and2b_1 _12875_ (.A_N(net319),
    .B(\div_shifter[52] ),
    .X(_06000_));
 sky130_fd_sc_hd__nand2b_1 _12876_ (.A_N(\div_shifter[52] ),
    .B(net319),
    .Y(_06001_));
 sky130_fd_sc_hd__and2b_1 _12877_ (.A_N(net325),
    .B(\div_shifter[51] ),
    .X(_06002_));
 sky130_fd_sc_hd__and2b_1 _12878_ (.A_N(net331),
    .B(net573),
    .X(_06003_));
 sky130_fd_sc_hd__nand2b_1 _12879_ (.A_N(net573),
    .B(net331),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2b_1 _12880_ (.A_N(net587),
    .B(net357),
    .Y(_06005_));
 sky130_fd_sc_hd__and2b_1 _12881_ (.A_N(net335),
    .B(\div_shifter[48] ),
    .X(_06006_));
 sky130_fd_sc_hd__nand2b_1 _12882_ (.A_N(\div_shifter[48] ),
    .B(net335),
    .Y(_06007_));
 sky130_fd_sc_hd__and2b_1 _12883_ (.A_N(net327),
    .B(net581),
    .X(_06008_));
 sky130_fd_sc_hd__nand2b_1 _12884_ (.A_N(net581),
    .B(net327),
    .Y(_06009_));
 sky130_fd_sc_hd__and2b_1 _12885_ (.A_N(net323),
    .B(net589),
    .X(_06011_));
 sky130_fd_sc_hd__nand2b_1 _12886_ (.A_N(net589),
    .B(net323),
    .Y(_06012_));
 sky130_fd_sc_hd__and2b_1 _12887_ (.A_N(net333),
    .B(\div_shifter[45] ),
    .X(_06013_));
 sky130_fd_sc_hd__nand2b_1 _12888_ (.A_N(\div_shifter[45] ),
    .B(net333),
    .Y(_06014_));
 sky130_fd_sc_hd__and2b_1 _12889_ (.A_N(net353),
    .B(\div_shifter[44] ),
    .X(_06015_));
 sky130_fd_sc_hd__nand2b_1 _12890_ (.A_N(\div_shifter[44] ),
    .B(net353),
    .Y(_06016_));
 sky130_fd_sc_hd__and2b_1 _12891_ (.A_N(net355),
    .B(net595),
    .X(_06017_));
 sky130_fd_sc_hd__nand2b_1 _12892_ (.A_N(net595),
    .B(net355),
    .Y(_06018_));
 sky130_fd_sc_hd__and2b_1 _12893_ (.A_N(net347),
    .B(net579),
    .X(_06019_));
 sky130_fd_sc_hd__nand2b_1 _12894_ (.A_N(net579),
    .B(net347),
    .Y(_06020_));
 sky130_fd_sc_hd__and2b_1 _12895_ (.A_N(net343),
    .B(\div_shifter[41] ),
    .X(_06022_));
 sky130_fd_sc_hd__nand2b_1 _12896_ (.A_N(\div_shifter[41] ),
    .B(net343),
    .Y(_06023_));
 sky130_fd_sc_hd__and2b_1 _12897_ (.A_N(net317),
    .B(net583),
    .X(_06024_));
 sky130_fd_sc_hd__nand2b_1 _12898_ (.A_N(net583),
    .B(net317),
    .Y(_06025_));
 sky130_fd_sc_hd__and2b_1 _12899_ (.A_N(net365),
    .B(\div_shifter[39] ),
    .X(_06026_));
 sky130_fd_sc_hd__nand2b_1 _12900_ (.A_N(\div_shifter[39] ),
    .B(net365),
    .Y(_06027_));
 sky130_fd_sc_hd__and2b_1 _12901_ (.A_N(net361),
    .B(net552),
    .X(_06028_));
 sky130_fd_sc_hd__nand2b_1 _12902_ (.A_N(net552),
    .B(net361),
    .Y(_06029_));
 sky130_fd_sc_hd__and2b_1 _12903_ (.A_N(net400),
    .B(net568),
    .X(_06030_));
 sky130_fd_sc_hd__nand2b_1 _12904_ (.A_N(net568),
    .B(net400),
    .Y(_06031_));
 sky130_fd_sc_hd__and2b_1 _12905_ (.A_N(net345),
    .B(\div_shifter[36] ),
    .X(_06033_));
 sky130_fd_sc_hd__nand2b_1 _12906_ (.A_N(\div_shifter[36] ),
    .B(net345),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2b_1 _12907_ (.A_N(_06033_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__and2b_1 _12908_ (.A_N(net359),
    .B(net594),
    .X(_06036_));
 sky130_fd_sc_hd__nand2b_1 _12909_ (.A_N(net594),
    .B(net359),
    .Y(_06037_));
 sky130_fd_sc_hd__nand2b_1 _12910_ (.A_N(_06036_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__and2b_1 _12911_ (.A_N(net398),
    .B(net550),
    .X(_06039_));
 sky130_fd_sc_hd__nand2b_1 _12912_ (.A_N(net550),
    .B(net398),
    .Y(_06040_));
 sky130_fd_sc_hd__and2b_1 _12913_ (.A_N(net337),
    .B(net554),
    .X(_06041_));
 sky130_fd_sc_hd__nand2b_1 _12914_ (.A_N(net554),
    .B(net337),
    .Y(_06042_));
 sky130_fd_sc_hd__and2b_1 _12915_ (.A_N(net442),
    .B(\div_shifter[32] ),
    .X(_06044_));
 sky130_fd_sc_hd__xnor2_1 _12916_ (.A(\div_shifter[32] ),
    .B(net442),
    .Y(_06045_));
 sky130_fd_sc_hd__nand2b_1 _12917_ (.A_N(net380),
    .B(net369),
    .Y(_06046_));
 sky130_fd_sc_hd__a21o_1 _12918_ (.A1(_06045_),
    .A2(_06046_),
    .B1(_06044_),
    .X(_06047_));
 sky130_fd_sc_hd__a21o_1 _12919_ (.A1(_06042_),
    .A2(_06047_),
    .B1(_06041_),
    .X(_06048_));
 sky130_fd_sc_hd__a21o_1 _12920_ (.A1(_06040_),
    .A2(_06048_),
    .B1(_06039_),
    .X(_06049_));
 sky130_fd_sc_hd__a21o_1 _12921_ (.A1(_06037_),
    .A2(_06049_),
    .B1(_06036_),
    .X(_06050_));
 sky130_fd_sc_hd__a21o_1 _12922_ (.A1(_06034_),
    .A2(_06050_),
    .B1(_06033_),
    .X(_06051_));
 sky130_fd_sc_hd__a21o_1 _12923_ (.A1(_06031_),
    .A2(_06051_),
    .B1(_06030_),
    .X(_06052_));
 sky130_fd_sc_hd__a21o_1 _12924_ (.A1(_06029_),
    .A2(_06052_),
    .B1(_06028_),
    .X(_06053_));
 sky130_fd_sc_hd__a21o_1 _12925_ (.A1(_06027_),
    .A2(_06053_),
    .B1(_06026_),
    .X(_06055_));
 sky130_fd_sc_hd__a21o_1 _12926_ (.A1(_06025_),
    .A2(_06055_),
    .B1(_06024_),
    .X(_06056_));
 sky130_fd_sc_hd__a21o_1 _12927_ (.A1(_06023_),
    .A2(_06056_),
    .B1(_06022_),
    .X(_06057_));
 sky130_fd_sc_hd__a21o_1 _12928_ (.A1(_06020_),
    .A2(_06057_),
    .B1(_06019_),
    .X(_06058_));
 sky130_fd_sc_hd__a21o_1 _12929_ (.A1(_06018_),
    .A2(_06058_),
    .B1(_06017_),
    .X(_06059_));
 sky130_fd_sc_hd__a21o_1 _12930_ (.A1(_06016_),
    .A2(_06059_),
    .B1(_06015_),
    .X(_06060_));
 sky130_fd_sc_hd__a21o_1 _12931_ (.A1(_06014_),
    .A2(_06060_),
    .B1(_06013_),
    .X(_06061_));
 sky130_fd_sc_hd__a21o_1 _12932_ (.A1(_06012_),
    .A2(_06061_),
    .B1(_06011_),
    .X(_06062_));
 sky130_fd_sc_hd__a21o_1 _12933_ (.A1(_06009_),
    .A2(_06062_),
    .B1(_06008_),
    .X(_06063_));
 sky130_fd_sc_hd__a21o_1 _12934_ (.A1(_06007_),
    .A2(_06063_),
    .B1(_06006_),
    .X(_06064_));
 sky130_fd_sc_hd__nand2b_1 _12935_ (.A_N(net357),
    .B(net587),
    .Y(_06066_));
 sky130_fd_sc_hd__a21bo_1 _12936_ (.A1(_06005_),
    .A2(_06064_),
    .B1_N(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__a21o_1 _12937_ (.A1(_06004_),
    .A2(_06067_),
    .B1(_06003_),
    .X(_06068_));
 sky130_fd_sc_hd__nand2b_1 _12938_ (.A_N(\div_shifter[51] ),
    .B(net325),
    .Y(_06069_));
 sky130_fd_sc_hd__nand2b_1 _12939_ (.A_N(_06002_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__a21o_1 _12940_ (.A1(_06068_),
    .A2(_06069_),
    .B1(_06002_),
    .X(_06071_));
 sky130_fd_sc_hd__a21o_1 _12941_ (.A1(_06001_),
    .A2(_06071_),
    .B1(_06000_),
    .X(_06072_));
 sky130_fd_sc_hd__nand2b_1 _12942_ (.A_N(net562),
    .B(net313),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2b_1 _12943_ (.A_N(_05998_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__a21o_1 _12944_ (.A1(_06072_),
    .A2(_06073_),
    .B1(_05998_),
    .X(_06075_));
 sky130_fd_sc_hd__a21o_1 _12945_ (.A1(_05997_),
    .A2(_06075_),
    .B1(_05996_),
    .X(_06077_));
 sky130_fd_sc_hd__nand2b_1 _12946_ (.A_N(\div_shifter[55] ),
    .B(net329),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2b_1 _12947_ (.A_N(_05995_),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__a21o_1 _12948_ (.A1(_06077_),
    .A2(_06078_),
    .B1(_05995_),
    .X(_06080_));
 sky130_fd_sc_hd__a21o_1 _12949_ (.A1(_05994_),
    .A2(_06080_),
    .B1(_05993_),
    .X(_06081_));
 sky130_fd_sc_hd__a21o_1 _12950_ (.A1(_05991_),
    .A2(_06081_),
    .B1(_05990_),
    .X(_06082_));
 sky130_fd_sc_hd__a21o_1 _12951_ (.A1(_05989_),
    .A2(_06082_),
    .B1(_05987_),
    .X(_06083_));
 sky130_fd_sc_hd__nand2b_1 _12952_ (.A_N(net566),
    .B(net450),
    .Y(_06084_));
 sky130_fd_sc_hd__nand2b_1 _12953_ (.A_N(_05986_),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__a21o_1 _12954_ (.A1(_06083_),
    .A2(_06084_),
    .B1(_05986_),
    .X(_06086_));
 sky130_fd_sc_hd__a21oi_1 _12955_ (.A1(_05985_),
    .A2(_06086_),
    .B1(_05984_),
    .Y(_06088_));
 sky130_fd_sc_hd__o21ba_1 _12956_ (.A1(_05982_),
    .A2(_06088_),
    .B1_N(_05981_),
    .X(_06089_));
 sky130_fd_sc_hd__a21boi_1 _12957_ (.A1(net396),
    .A2(_06089_),
    .B1_N(net560),
    .Y(_06090_));
 sky130_fd_sc_hd__nor2_1 _12958_ (.A(net396),
    .B(_06089_),
    .Y(_06091_));
 sky130_fd_sc_hd__or2_2 _12959_ (.A(_06090_),
    .B(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__a22o_1 _12960_ (.A1(net600),
    .A2(net221),
    .B1(net2),
    .B2(net277),
    .X(_06093_));
 sky130_fd_sc_hd__and2_1 _12961_ (.A(net295),
    .B(_06093_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _12962_ (.A1(\div_res[0] ),
    .A2(net277),
    .B1(net221),
    .B2(net558),
    .X(_06094_));
 sky130_fd_sc_hd__and2_1 _12963_ (.A(net295),
    .B(net559),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _12964_ (.A1(\div_res[1] ),
    .A2(net277),
    .B1(net221),
    .B2(net548),
    .X(_06095_));
 sky130_fd_sc_hd__and2_1 _12965_ (.A(net295),
    .B(net549),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _12966_ (.A1(\div_res[2] ),
    .A2(net277),
    .B1(net221),
    .B2(net507),
    .X(_06097_));
 sky130_fd_sc_hd__and2_1 _12967_ (.A(net295),
    .B(net508),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _12968_ (.A1(net507),
    .A2(net275),
    .B1(net220),
    .B2(net497),
    .X(_06098_));
 sky130_fd_sc_hd__and2_1 _12969_ (.A(net294),
    .B(net545),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _12970_ (.A1(net497),
    .A2(net275),
    .B1(net220),
    .B2(net495),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _12971_ (.A(net294),
    .B(net498),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _12972_ (.A1(net495),
    .A2(net276),
    .B1(net220),
    .B2(net467),
    .X(_06100_));
 sky130_fd_sc_hd__and2_1 _12973_ (.A(net294),
    .B(net496),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _12974_ (.A1(net467),
    .A2(net276),
    .B1(net220),
    .B2(\div_res[7] ),
    .X(_06101_));
 sky130_fd_sc_hd__and2_1 _12975_ (.A(net294),
    .B(net468),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _12976_ (.A1(\div_res[7] ),
    .A2(net276),
    .B1(net219),
    .B2(net530),
    .X(_06103_));
 sky130_fd_sc_hd__and2_1 _12977_ (.A(net293),
    .B(net531),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _12978_ (.A1(net530),
    .A2(net275),
    .B1(net219),
    .B2(net540),
    .X(_06104_));
 sky130_fd_sc_hd__and2_1 _12979_ (.A(net293),
    .B(net543),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _12980_ (.A1(net540),
    .A2(net275),
    .B1(net219),
    .B2(net513),
    .X(_06105_));
 sky130_fd_sc_hd__and2_1 _12981_ (.A(net293),
    .B(net541),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _12982_ (.A1(net513),
    .A2(net275),
    .B1(net219),
    .B2(net499),
    .X(_06106_));
 sky130_fd_sc_hd__and2_1 _12983_ (.A(net293),
    .B(net514),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _12984_ (.A1(net499),
    .A2(net275),
    .B1(net219),
    .B2(\div_res[12] ),
    .X(_06107_));
 sky130_fd_sc_hd__and2_1 _12985_ (.A(net293),
    .B(net500),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _12986_ (.A1(\div_res[12] ),
    .A2(net275),
    .B1(net219),
    .B2(net522),
    .X(_06109_));
 sky130_fd_sc_hd__and2_1 _12987_ (.A(net293),
    .B(net523),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _12988_ (.A1(net522),
    .A2(net275),
    .B1(net219),
    .B2(net515),
    .X(_06110_));
 sky130_fd_sc_hd__and2_1 _12989_ (.A(net293),
    .B(net539),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _12990_ (.A1(net515),
    .A2(net275),
    .B1(net219),
    .B2(net493),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _12991_ (.A(net293),
    .B(net516),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _12992_ (.A1(net493),
    .A2(net275),
    .B1(net219),
    .B2(net484),
    .X(_06112_));
 sky130_fd_sc_hd__and2_1 _12993_ (.A(net293),
    .B(net494),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _12994_ (.A1(net484),
    .A2(net275),
    .B1(net219),
    .B2(\div_res[17] ),
    .X(_06113_));
 sky130_fd_sc_hd__and2_1 _12995_ (.A(net293),
    .B(net485),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _12996_ (.A1(\div_res[17] ),
    .A2(net275),
    .B1(net219),
    .B2(net510),
    .X(_06115_));
 sky130_fd_sc_hd__and2_1 _12997_ (.A(net293),
    .B(net511),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _12998_ (.A1(\div_res[18] ),
    .A2(net275),
    .B1(net219),
    .B2(net487),
    .X(_06116_));
 sky130_fd_sc_hd__and2_1 _12999_ (.A(net293),
    .B(net488),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _13000_ (.A1(net487),
    .A2(net275),
    .B1(net219),
    .B2(net520),
    .X(_06117_));
 sky130_fd_sc_hd__and2_1 _13001_ (.A(net293),
    .B(net521),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _13002_ (.A1(net520),
    .A2(net275),
    .B1(net219),
    .B2(net546),
    .X(_06118_));
 sky130_fd_sc_hd__and2_1 _13003_ (.A(net294),
    .B(net547),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _13004_ (.A1(\div_res[21] ),
    .A2(net275),
    .B1(net219),
    .B2(net535),
    .X(_06119_));
 sky130_fd_sc_hd__and2_1 _13005_ (.A(net294),
    .B(net536),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _13006_ (.A1(\div_res[22] ),
    .A2(net276),
    .B1(net219),
    .B2(net502),
    .X(_06121_));
 sky130_fd_sc_hd__and2_1 _13007_ (.A(net293),
    .B(net503),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _13008_ (.A1(net502),
    .A2(net276),
    .B1(net220),
    .B2(net528),
    .X(_06122_));
 sky130_fd_sc_hd__and2_1 _13009_ (.A(net294),
    .B(net529),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _13010_ (.A1(\div_res[24] ),
    .A2(net276),
    .B1(net220),
    .B2(net517),
    .X(_06123_));
 sky130_fd_sc_hd__and2_1 _13011_ (.A(net293),
    .B(net518),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _13012_ (.A1(\div_res[25] ),
    .A2(net276),
    .B1(net220),
    .B2(net490),
    .X(_06124_));
 sky130_fd_sc_hd__and2_1 _13013_ (.A(net293),
    .B(net491),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _13014_ (.A1(net490),
    .A2(net276),
    .B1(net220),
    .B2(net505),
    .X(_06125_));
 sky130_fd_sc_hd__and2_1 _13015_ (.A(net295),
    .B(net534),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _13016_ (.A1(net505),
    .A2(net276),
    .B1(net220),
    .B2(net479),
    .X(_06127_));
 sky130_fd_sc_hd__and2_1 _13017_ (.A(net295),
    .B(net506),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _13018_ (.A1(net479),
    .A2(net277),
    .B1(net221),
    .B2(\div_res[29] ),
    .X(_06128_));
 sky130_fd_sc_hd__and2_1 _13019_ (.A(net295),
    .B(net480),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _13020_ (.A1(\div_res[29] ),
    .A2(net277),
    .B1(net221),
    .B2(net525),
    .X(_06129_));
 sky130_fd_sc_hd__and2_1 _13021_ (.A(net295),
    .B(net526),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _13022_ (.A1(\div_res[30] ),
    .A2(net277),
    .B1(net221),
    .B2(net428),
    .X(_06130_));
 sky130_fd_sc_hd__and2_1 _13023_ (.A(net295),
    .B(net429),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _13024_ (.A1(net405),
    .A2(net222),
    .B1(net202),
    .B2(reg1_val[0]),
    .X(_06131_));
 sky130_fd_sc_hd__and2_1 _13025_ (.A(net302),
    .B(net406),
    .X(_00066_));
 sky130_fd_sc_hd__o221a_1 _13026_ (.A1(net405),
    .A2(net274),
    .B1(net218),
    .B2(net414),
    .C1(net300),
    .X(_06133_));
 sky130_fd_sc_hd__o21a_1 _13027_ (.A1(_00213_),
    .A2(net198),
    .B1(net422),
    .X(_00067_));
 sky130_fd_sc_hd__o221a_1 _13028_ (.A1(net414),
    .A2(net274),
    .B1(net218),
    .B2(\div_shifter[2] ),
    .C1(net300),
    .X(_06134_));
 sky130_fd_sc_hd__a21boi_1 _13029_ (.A1(_00216_),
    .A2(net202),
    .B1_N(net415),
    .Y(_00068_));
 sky130_fd_sc_hd__a21oi_1 _13030_ (.A1(_04395_),
    .A2(net278),
    .B1(rst),
    .Y(_06135_));
 sky130_fd_sc_hd__o221a_1 _13031_ (.A1(net367),
    .A2(net218),
    .B1(_00210_),
    .B2(net198),
    .C1(_06135_),
    .X(_00069_));
 sky130_fd_sc_hd__a221o_1 _13032_ (.A1(_04384_),
    .A2(net278),
    .B1(net222),
    .B2(net390),
    .C1(rst),
    .X(_06136_));
 sky130_fd_sc_hd__a21oi_1 _13033_ (.A1(_00252_),
    .A2(net202),
    .B1(net391),
    .Y(_00070_));
 sky130_fd_sc_hd__a21oi_1 _13034_ (.A1(_04373_),
    .A2(net278),
    .B1(rst),
    .Y(_06137_));
 sky130_fd_sc_hd__o221a_1 _13035_ (.A1(net315),
    .A2(net218),
    .B1(_00249_),
    .B2(net197),
    .C1(_06137_),
    .X(_00071_));
 sky130_fd_sc_hd__o221a_1 _13036_ (.A1(net315),
    .A2(net274),
    .B1(net218),
    .B2(net458),
    .C1(net300),
    .X(_06139_));
 sky130_fd_sc_hd__a21boi_1 _13037_ (.A1(_00276_),
    .A2(net202),
    .B1_N(net459),
    .Y(_00072_));
 sky130_fd_sc_hd__o221a_1 _13038_ (.A1(net458),
    .A2(net274),
    .B1(net218),
    .B2(net465),
    .C1(net300),
    .X(_06140_));
 sky130_fd_sc_hd__a21boi_1 _13039_ (.A1(net194),
    .A2(net202),
    .B1_N(net466),
    .Y(_00073_));
 sky130_fd_sc_hd__o221a_1 _13040_ (.A1(\div_shifter[7] ),
    .A2(net274),
    .B1(net218),
    .B2(net455),
    .C1(net300),
    .X(_06141_));
 sky130_fd_sc_hd__a21boi_1 _13041_ (.A1(_00306_),
    .A2(net202),
    .B1_N(net456),
    .Y(_00074_));
 sky130_fd_sc_hd__o221a_1 _13042_ (.A1(\div_shifter[8] ),
    .A2(net274),
    .B1(net218),
    .B2(net452),
    .C1(net300),
    .X(_06142_));
 sky130_fd_sc_hd__a21boi_1 _13043_ (.A1(net168),
    .A2(net202),
    .B1_N(net453),
    .Y(_00075_));
 sky130_fd_sc_hd__o221a_1 _13044_ (.A1(net452),
    .A2(net274),
    .B1(net217),
    .B2(net460),
    .C1(net300),
    .X(_06143_));
 sky130_fd_sc_hd__a21boi_1 _13045_ (.A1(_00292_),
    .A2(net203),
    .B1_N(net461),
    .Y(_00076_));
 sky130_fd_sc_hd__o221a_1 _13046_ (.A1(\div_shifter[10] ),
    .A2(net274),
    .B1(net218),
    .B2(net444),
    .C1(net300),
    .X(_06145_));
 sky130_fd_sc_hd__o21a_1 _13047_ (.A1(_06470_),
    .A2(net197),
    .B1(net445),
    .X(_00077_));
 sky130_fd_sc_hd__o221a_1 _13048_ (.A1(net444),
    .A2(net274),
    .B1(net218),
    .B2(net474),
    .C1(net300),
    .X(_06146_));
 sky130_fd_sc_hd__a21boi_1 _13049_ (.A1(_06472_),
    .A2(net202),
    .B1_N(net475),
    .Y(_00078_));
 sky130_fd_sc_hd__o221a_1 _13050_ (.A1(\div_shifter[12] ),
    .A2(net274),
    .B1(net218),
    .B2(net462),
    .C1(net299),
    .X(_06147_));
 sky130_fd_sc_hd__a21boi_1 _13051_ (.A1(net153),
    .A2(net202),
    .B1_N(net463),
    .Y(_00079_));
 sky130_fd_sc_hd__o221a_1 _13052_ (.A1(net462),
    .A2(net273),
    .B1(net217),
    .B2(net431),
    .C1(net299),
    .X(_06148_));
 sky130_fd_sc_hd__a21boi_1 _13053_ (.A1(_06503_),
    .A2(net201),
    .B1_N(net473),
    .Y(_00080_));
 sky130_fd_sc_hd__o221a_1 _13054_ (.A1(net431),
    .A2(net273),
    .B1(net217),
    .B2(net386),
    .C1(net299),
    .X(_06149_));
 sky130_fd_sc_hd__o21a_1 _13055_ (.A1(_06499_),
    .A2(net197),
    .B1(net432),
    .X(_00081_));
 sky130_fd_sc_hd__o221a_1 _13056_ (.A1(net386),
    .A2(net273),
    .B1(net217),
    .B2(\div_shifter[16] ),
    .C1(net297),
    .X(_06151_));
 sky130_fd_sc_hd__o21a_1 _13057_ (.A1(_00159_),
    .A2(net197),
    .B1(net387),
    .X(_00082_));
 sky130_fd_sc_hd__o221a_1 _13058_ (.A1(\div_shifter[16] ),
    .A2(net273),
    .B1(net217),
    .B2(net447),
    .C1(net297),
    .X(_06152_));
 sky130_fd_sc_hd__o21a_1 _13059_ (.A1(net101),
    .A2(net197),
    .B1(net448),
    .X(_00083_));
 sky130_fd_sc_hd__o221a_1 _13060_ (.A1(\div_shifter[17] ),
    .A2(net273),
    .B1(net217),
    .B2(net402),
    .C1(net297),
    .X(_06153_));
 sky130_fd_sc_hd__o21a_1 _13061_ (.A1(_00187_),
    .A2(net197),
    .B1(net403),
    .X(_00084_));
 sky130_fd_sc_hd__o221a_1 _13062_ (.A1(net402),
    .A2(net273),
    .B1(net217),
    .B2(net409),
    .C1(net297),
    .X(_06154_));
 sky130_fd_sc_hd__o21a_1 _13063_ (.A1(_00174_),
    .A2(net197),
    .B1(net410),
    .X(_00085_));
 sky130_fd_sc_hd__o221a_1 _13064_ (.A1(net409),
    .A2(net273),
    .B1(net217),
    .B2(net440),
    .C1(net297),
    .X(_06155_));
 sky130_fd_sc_hd__o21a_1 _13065_ (.A1(_00175_),
    .A2(net197),
    .B1(net441),
    .X(_00086_));
 sky130_fd_sc_hd__o221a_1 _13066_ (.A1(\div_shifter[20] ),
    .A2(net273),
    .B1(net217),
    .B2(net433),
    .C1(net299),
    .X(_06157_));
 sky130_fd_sc_hd__o21a_1 _13067_ (.A1(net103),
    .A2(net197),
    .B1(net434),
    .X(_00087_));
 sky130_fd_sc_hd__o221a_1 _13068_ (.A1(net433),
    .A2(net273),
    .B1(net217),
    .B2(net426),
    .C1(net299),
    .X(_06158_));
 sky130_fd_sc_hd__o21a_1 _13069_ (.A1(_06551_),
    .A2(net198),
    .B1(net437),
    .X(_00088_));
 sky130_fd_sc_hd__o221a_1 _13070_ (.A1(net426),
    .A2(net273),
    .B1(net217),
    .B2(net417),
    .C1(net299),
    .X(_06159_));
 sky130_fd_sc_hd__o21a_1 _13071_ (.A1(net107),
    .A2(net198),
    .B1(net427),
    .X(_00089_));
 sky130_fd_sc_hd__o221a_1 _13072_ (.A1(net417),
    .A2(net273),
    .B1(net217),
    .B2(net407),
    .C1(net299),
    .X(_06160_));
 sky130_fd_sc_hd__o21a_1 _13073_ (.A1(_00136_),
    .A2(net198),
    .B1(net418),
    .X(_00090_));
 sky130_fd_sc_hd__o221a_1 _13074_ (.A1(net407),
    .A2(net273),
    .B1(net217),
    .B2(net377),
    .C1(net299),
    .X(_06161_));
 sky130_fd_sc_hd__o21a_1 _13075_ (.A1(net110),
    .A2(net198),
    .B1(net408),
    .X(_00091_));
 sky130_fd_sc_hd__o221a_1 _13076_ (.A1(net377),
    .A2(net273),
    .B1(net217),
    .B2(\div_shifter[26] ),
    .C1(net299),
    .X(_06163_));
 sky130_fd_sc_hd__o21a_1 _13077_ (.A1(_06531_),
    .A2(net198),
    .B1(net378),
    .X(_00092_));
 sky130_fd_sc_hd__o221a_1 _13078_ (.A1(\div_shifter[26] ),
    .A2(net273),
    .B1(net217),
    .B2(net423),
    .C1(net299),
    .X(_06164_));
 sky130_fd_sc_hd__o21a_1 _13079_ (.A1(_06523_),
    .A2(net197),
    .B1(net424),
    .X(_00093_));
 sky130_fd_sc_hd__o221a_1 _13080_ (.A1(net423),
    .A2(net273),
    .B1(net217),
    .B2(net382),
    .C1(net299),
    .X(_06165_));
 sky130_fd_sc_hd__o21a_1 _13081_ (.A1(_00350_),
    .A2(net197),
    .B1(net439),
    .X(_00094_));
 sky130_fd_sc_hd__a221o_1 _13082_ (.A1(net383),
    .A2(net278),
    .B1(net222),
    .B2(_04351_),
    .C1(rst),
    .X(_06166_));
 sky130_fd_sc_hd__a21oi_1 _13083_ (.A1(net78),
    .A2(net202),
    .B1(net384),
    .Y(_00095_));
 sky130_fd_sc_hd__a221o_1 _13084_ (.A1(net393),
    .A2(net278),
    .B1(net222),
    .B2(_04340_),
    .C1(rst),
    .X(_06167_));
 sky130_fd_sc_hd__a21oi_1 _13085_ (.A1(_00456_),
    .A2(net202),
    .B1(net394),
    .Y(_00096_));
 sky130_fd_sc_hd__a21oi_1 _13086_ (.A1(_04340_),
    .A2(net278),
    .B1(rst),
    .Y(_06169_));
 sky130_fd_sc_hd__o221a_1 _13087_ (.A1(net380),
    .A2(net218),
    .B1(_00595_),
    .B2(net197),
    .C1(_06169_),
    .X(_00097_));
 sky130_fd_sc_hd__nand3_1 _13088_ (.A(net380),
    .B(net369),
    .C(net1),
    .Y(_06170_));
 sky130_fd_sc_hd__a21o_1 _13089_ (.A1(net369),
    .A2(net1),
    .B1(net380),
    .X(_06171_));
 sky130_fd_sc_hd__a32o_1 _13090_ (.A1(net278),
    .A2(net612),
    .A3(_06171_),
    .B1(net222),
    .B2(net570),
    .X(_06172_));
 sky130_fd_sc_hd__and2_1 _13091_ (.A(net300),
    .B(net613),
    .X(_00098_));
 sky130_fd_sc_hd__xor2_1 _13092_ (.A(_06045_),
    .B(_06046_),
    .X(_06173_));
 sky130_fd_sc_hd__mux2_1 _13093_ (.A0(\div_shifter[32] ),
    .A1(_06173_),
    .S(net1),
    .X(_06174_));
 sky130_fd_sc_hd__a22o_1 _13094_ (.A1(net554),
    .A2(net222),
    .B1(_06174_),
    .B2(net278),
    .X(_06175_));
 sky130_fd_sc_hd__and2_1 _13095_ (.A(net301),
    .B(net555),
    .X(_00099_));
 sky130_fd_sc_hd__nand2b_1 _13096_ (.A_N(_06041_),
    .B(_06042_),
    .Y(_06177_));
 sky130_fd_sc_hd__xnor2_1 _13097_ (.A(_06047_),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__mux2_1 _13098_ (.A0(\div_shifter[33] ),
    .A1(_06178_),
    .S(net1),
    .X(_06179_));
 sky130_fd_sc_hd__a22o_1 _13099_ (.A1(net550),
    .A2(net222),
    .B1(_06179_),
    .B2(net278),
    .X(_06180_));
 sky130_fd_sc_hd__and2_1 _13100_ (.A(net301),
    .B(net551),
    .X(_00100_));
 sky130_fd_sc_hd__nand2b_1 _13101_ (.A_N(_06039_),
    .B(_06040_),
    .Y(_06181_));
 sky130_fd_sc_hd__xnor2_1 _13102_ (.A(_06048_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__mux2_1 _13103_ (.A0(net550),
    .A1(_06182_),
    .S(net1),
    .X(_06183_));
 sky130_fd_sc_hd__a22o_1 _13104_ (.A1(net594),
    .A2(net222),
    .B1(_06183_),
    .B2(net278),
    .X(_06184_));
 sky130_fd_sc_hd__and2_1 _13105_ (.A(net301),
    .B(_06184_),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _13106_ (.A(_06038_),
    .B(_06049_),
    .Y(_06186_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(net594),
    .A1(_06186_),
    .S(net1),
    .X(_06187_));
 sky130_fd_sc_hd__a22o_1 _13108_ (.A1(net601),
    .A2(net222),
    .B1(_06187_),
    .B2(net278),
    .X(_06188_));
 sky130_fd_sc_hd__and2_1 _13109_ (.A(net300),
    .B(_06188_),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _13110_ (.A(_06035_),
    .B(_06050_),
    .Y(_06189_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(\div_shifter[36] ),
    .A1(_06189_),
    .S(net2),
    .X(_06190_));
 sky130_fd_sc_hd__a22o_1 _13112_ (.A1(net568),
    .A2(net222),
    .B1(_06190_),
    .B2(net278),
    .X(_06191_));
 sky130_fd_sc_hd__and2_1 _13113_ (.A(net299),
    .B(net569),
    .X(_00103_));
 sky130_fd_sc_hd__nand2b_1 _13114_ (.A_N(_06030_),
    .B(_06031_),
    .Y(_06192_));
 sky130_fd_sc_hd__xnor2_1 _13115_ (.A(_06051_),
    .B(_06192_),
    .Y(_06194_));
 sky130_fd_sc_hd__mux2_1 _13116_ (.A0(\div_shifter[37] ),
    .A1(_06194_),
    .S(net1),
    .X(_06195_));
 sky130_fd_sc_hd__a22o_1 _13117_ (.A1(net552),
    .A2(net223),
    .B1(_06195_),
    .B2(net280),
    .X(_06196_));
 sky130_fd_sc_hd__and2_1 _13118_ (.A(net297),
    .B(net553),
    .X(_00104_));
 sky130_fd_sc_hd__nand2b_1 _13119_ (.A_N(_06028_),
    .B(_06029_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_1 _13120_ (.A(_06052_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(net552),
    .A1(_06198_),
    .S(net1),
    .X(_06199_));
 sky130_fd_sc_hd__a22o_1 _13122_ (.A1(net604),
    .A2(net223),
    .B1(_06199_),
    .B2(net280),
    .X(_06200_));
 sky130_fd_sc_hd__and2_1 _13123_ (.A(net297),
    .B(_06200_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2b_1 _13124_ (.A_N(_06026_),
    .B(_06027_),
    .Y(_06201_));
 sky130_fd_sc_hd__xnor2_1 _13125_ (.A(_06053_),
    .B(_06201_),
    .Y(_06203_));
 sky130_fd_sc_hd__mux2_1 _13126_ (.A0(\div_shifter[39] ),
    .A1(_06203_),
    .S(net1),
    .X(_06204_));
 sky130_fd_sc_hd__a22o_1 _13127_ (.A1(net583),
    .A2(net223),
    .B1(_06204_),
    .B2(net280),
    .X(_06205_));
 sky130_fd_sc_hd__and2_1 _13128_ (.A(net297),
    .B(net584),
    .X(_00106_));
 sky130_fd_sc_hd__nand2b_1 _13129_ (.A_N(_06024_),
    .B(_06025_),
    .Y(_06206_));
 sky130_fd_sc_hd__xnor2_1 _13130_ (.A(_06055_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__mux2_1 _13131_ (.A0(net583),
    .A1(_06207_),
    .S(net1),
    .X(_06208_));
 sky130_fd_sc_hd__a22o_1 _13132_ (.A1(net598),
    .A2(net223),
    .B1(_06208_),
    .B2(net280),
    .X(_06209_));
 sky130_fd_sc_hd__and2_1 _13133_ (.A(net298),
    .B(net599),
    .X(_00107_));
 sky130_fd_sc_hd__nand2b_1 _13134_ (.A_N(_06022_),
    .B(_06023_),
    .Y(_06210_));
 sky130_fd_sc_hd__xnor2_1 _13135_ (.A(_06056_),
    .B(_06210_),
    .Y(_06212_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(\div_shifter[41] ),
    .A1(_06212_),
    .S(net1),
    .X(_06213_));
 sky130_fd_sc_hd__a22o_1 _13137_ (.A1(net579),
    .A2(net223),
    .B1(_06213_),
    .B2(net280),
    .X(_06214_));
 sky130_fd_sc_hd__and2_1 _13138_ (.A(net298),
    .B(net580),
    .X(_00108_));
 sky130_fd_sc_hd__nand2b_1 _13139_ (.A_N(_06019_),
    .B(_06020_),
    .Y(_06215_));
 sky130_fd_sc_hd__xnor2_1 _13140_ (.A(_06057_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__mux2_1 _13141_ (.A0(net579),
    .A1(_06216_),
    .S(net1),
    .X(_06217_));
 sky130_fd_sc_hd__a22o_1 _13142_ (.A1(net595),
    .A2(net223),
    .B1(_06217_),
    .B2(net280),
    .X(_06218_));
 sky130_fd_sc_hd__and2_1 _13143_ (.A(net298),
    .B(net596),
    .X(_00109_));
 sky130_fd_sc_hd__nand2b_1 _13144_ (.A_N(_06017_),
    .B(_06018_),
    .Y(_06219_));
 sky130_fd_sc_hd__xnor2_1 _13145_ (.A(_06058_),
    .B(_06219_),
    .Y(_06221_));
 sky130_fd_sc_hd__mux2_1 _13146_ (.A0(net595),
    .A1(_06221_),
    .S(net1),
    .X(_06222_));
 sky130_fd_sc_hd__a22o_1 _13147_ (.A1(net597),
    .A2(_06432_),
    .B1(_06222_),
    .B2(net279),
    .X(_06223_));
 sky130_fd_sc_hd__and2_1 _13148_ (.A(net301),
    .B(_06223_),
    .X(_00110_));
 sky130_fd_sc_hd__nand2b_1 _13149_ (.A_N(_06015_),
    .B(_06016_),
    .Y(_06224_));
 sky130_fd_sc_hd__xnor2_1 _13150_ (.A(_06059_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(\div_shifter[44] ),
    .A1(_06225_),
    .S(net1),
    .X(_06226_));
 sky130_fd_sc_hd__a22o_1 _13152_ (.A1(net592),
    .A2(_06432_),
    .B1(_06226_),
    .B2(net279),
    .X(_06227_));
 sky130_fd_sc_hd__and2_1 _13153_ (.A(net301),
    .B(net593),
    .X(_00111_));
 sky130_fd_sc_hd__nand2b_1 _13154_ (.A_N(_06013_),
    .B(_06014_),
    .Y(_06228_));
 sky130_fd_sc_hd__xnor2_1 _13155_ (.A(_06060_),
    .B(_06228_),
    .Y(_06230_));
 sky130_fd_sc_hd__mux2_1 _13156_ (.A0(\div_shifter[45] ),
    .A1(_06230_),
    .S(net2),
    .X(_06231_));
 sky130_fd_sc_hd__a22o_1 _13157_ (.A1(net589),
    .A2(net222),
    .B1(_06231_),
    .B2(net279),
    .X(_06232_));
 sky130_fd_sc_hd__and2_1 _13158_ (.A(net302),
    .B(net590),
    .X(_00112_));
 sky130_fd_sc_hd__nand2b_1 _13159_ (.A_N(_06011_),
    .B(_06012_),
    .Y(_06233_));
 sky130_fd_sc_hd__xnor2_1 _13160_ (.A(_06061_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__mux2_1 _13161_ (.A0(\div_shifter[46] ),
    .A1(_06234_),
    .S(_06092_),
    .X(_06235_));
 sky130_fd_sc_hd__a22o_1 _13162_ (.A1(net581),
    .A2(_06432_),
    .B1(_06235_),
    .B2(net279),
    .X(_06236_));
 sky130_fd_sc_hd__and2_1 _13163_ (.A(net301),
    .B(net582),
    .X(_00113_));
 sky130_fd_sc_hd__nand2b_1 _13164_ (.A_N(_06008_),
    .B(_06009_),
    .Y(_06237_));
 sky130_fd_sc_hd__xnor2_1 _13165_ (.A(_06062_),
    .B(_06237_),
    .Y(_06239_));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(net581),
    .A1(_06239_),
    .S(_06092_),
    .X(_06240_));
 sky130_fd_sc_hd__a22o_1 _13167_ (.A1(net602),
    .A2(net223),
    .B1(_06240_),
    .B2(net279),
    .X(_06241_));
 sky130_fd_sc_hd__and2_1 _13168_ (.A(net301),
    .B(_06241_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2b_1 _13169_ (.A_N(_06006_),
    .B(_06007_),
    .Y(_06242_));
 sky130_fd_sc_hd__xnor2_1 _13170_ (.A(_06063_),
    .B(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__mux2_1 _13171_ (.A0(\div_shifter[48] ),
    .A1(_06243_),
    .S(net2),
    .X(_06244_));
 sky130_fd_sc_hd__a22o_1 _13172_ (.A1(net587),
    .A2(_06432_),
    .B1(_06244_),
    .B2(net279),
    .X(_06245_));
 sky130_fd_sc_hd__and2_1 _13173_ (.A(net301),
    .B(net588),
    .X(_00115_));
 sky130_fd_sc_hd__nand2_1 _13174_ (.A(_06005_),
    .B(_06066_),
    .Y(_06246_));
 sky130_fd_sc_hd__xnor2_1 _13175_ (.A(_06064_),
    .B(_06246_),
    .Y(_06248_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(\div_shifter[49] ),
    .A1(_06248_),
    .S(net1),
    .X(_06249_));
 sky130_fd_sc_hd__a22o_1 _13177_ (.A1(net573),
    .A2(net223),
    .B1(_06249_),
    .B2(net280),
    .X(_06250_));
 sky130_fd_sc_hd__and2_1 _13178_ (.A(net298),
    .B(net574),
    .X(_00116_));
 sky130_fd_sc_hd__nand2b_1 _13179_ (.A_N(_06003_),
    .B(_06004_),
    .Y(_06251_));
 sky130_fd_sc_hd__xnor2_1 _13180_ (.A(_06067_),
    .B(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(net573),
    .A1(_06252_),
    .S(net1),
    .X(_06253_));
 sky130_fd_sc_hd__a22o_1 _13182_ (.A1(net603),
    .A2(net223),
    .B1(_06253_),
    .B2(net280),
    .X(_06254_));
 sky130_fd_sc_hd__and2_1 _13183_ (.A(net298),
    .B(_06254_),
    .X(_00117_));
 sky130_fd_sc_hd__xnor2_1 _13184_ (.A(_06068_),
    .B(_06070_),
    .Y(_06255_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(\div_shifter[51] ),
    .A1(_06255_),
    .S(net2),
    .X(_06257_));
 sky130_fd_sc_hd__a22o_1 _13186_ (.A1(net585),
    .A2(net221),
    .B1(_06257_),
    .B2(net277),
    .X(_06258_));
 sky130_fd_sc_hd__and2_1 _13187_ (.A(net296),
    .B(net586),
    .X(_00118_));
 sky130_fd_sc_hd__nand2b_1 _13188_ (.A_N(_06000_),
    .B(_06001_),
    .Y(_06259_));
 sky130_fd_sc_hd__xnor2_1 _13189_ (.A(_06071_),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(\div_shifter[52] ),
    .A1(_06260_),
    .S(net2),
    .X(_06261_));
 sky130_fd_sc_hd__a22o_1 _13191_ (.A1(net562),
    .A2(net221),
    .B1(_06261_),
    .B2(net277),
    .X(_06262_));
 sky130_fd_sc_hd__and2_1 _13192_ (.A(net295),
    .B(net563),
    .X(_00119_));
 sky130_fd_sc_hd__xnor2_1 _13193_ (.A(_06072_),
    .B(_06074_),
    .Y(_06263_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(\div_shifter[53] ),
    .A1(_06263_),
    .S(net2),
    .X(_06264_));
 sky130_fd_sc_hd__a22o_1 _13195_ (.A1(net556),
    .A2(net221),
    .B1(_06264_),
    .B2(net277),
    .X(_06266_));
 sky130_fd_sc_hd__and2_1 _13196_ (.A(net295),
    .B(net557),
    .X(_00120_));
 sky130_fd_sc_hd__nand2b_1 _13197_ (.A_N(_05996_),
    .B(_05997_),
    .Y(_06267_));
 sky130_fd_sc_hd__xnor2_1 _13198_ (.A(_06075_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__mux2_1 _13199_ (.A0(net556),
    .A1(_06268_),
    .S(net2),
    .X(_06269_));
 sky130_fd_sc_hd__a22o_1 _13200_ (.A1(net575),
    .A2(net221),
    .B1(_06269_),
    .B2(net277),
    .X(_06270_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(net295),
    .B(_06270_),
    .X(_00121_));
 sky130_fd_sc_hd__xnor2_1 _13202_ (.A(_06077_),
    .B(_06079_),
    .Y(_06271_));
 sky130_fd_sc_hd__mux2_1 _13203_ (.A0(\div_shifter[55] ),
    .A1(_06271_),
    .S(net2),
    .X(_06272_));
 sky130_fd_sc_hd__a22o_1 _13204_ (.A1(net564),
    .A2(net221),
    .B1(_06272_),
    .B2(net277),
    .X(_06273_));
 sky130_fd_sc_hd__and2_1 _13205_ (.A(net296),
    .B(net565),
    .X(_00122_));
 sky130_fd_sc_hd__nand2b_1 _13206_ (.A_N(_05993_),
    .B(_05994_),
    .Y(_06275_));
 sky130_fd_sc_hd__xnor2_1 _13207_ (.A(_06080_),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(net564),
    .A1(_06276_),
    .S(net2),
    .X(_06277_));
 sky130_fd_sc_hd__a22o_1 _13209_ (.A1(net571),
    .A2(net221),
    .B1(_06277_),
    .B2(net277),
    .X(_06278_));
 sky130_fd_sc_hd__and2_1 _13210_ (.A(net296),
    .B(net572),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_1 _13211_ (.A(_05992_),
    .B(_06081_),
    .Y(_06279_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(net571),
    .A1(_06279_),
    .S(net2),
    .X(_06280_));
 sky130_fd_sc_hd__a22o_1 _13213_ (.A1(net591),
    .A2(net221),
    .B1(_06280_),
    .B2(net277),
    .X(_06281_));
 sky130_fd_sc_hd__and2_1 _13214_ (.A(net295),
    .B(_06281_),
    .X(_00124_));
 sky130_fd_sc_hd__nand2b_1 _13215_ (.A_N(_05987_),
    .B(_05989_),
    .Y(_06283_));
 sky130_fd_sc_hd__xnor2_1 _13216_ (.A(_06082_),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(\div_shifter[58] ),
    .A1(_06284_),
    .S(net2),
    .X(_06285_));
 sky130_fd_sc_hd__a22o_1 _13218_ (.A1(net566),
    .A2(net223),
    .B1(_06285_),
    .B2(net280),
    .X(_06286_));
 sky130_fd_sc_hd__and2_1 _13219_ (.A(net298),
    .B(net567),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_1 _13220_ (.A(_06083_),
    .B(_06085_),
    .Y(_06287_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(net566),
    .A1(_06287_),
    .S(net2),
    .X(_06288_));
 sky130_fd_sc_hd__a22o_1 _13222_ (.A1(net576),
    .A2(net223),
    .B1(_06288_),
    .B2(net280),
    .X(_06289_));
 sky130_fd_sc_hd__and2_1 _13223_ (.A(net298),
    .B(net577),
    .X(_00126_));
 sky130_fd_sc_hd__nand2b_1 _13224_ (.A_N(_05984_),
    .B(_05985_),
    .Y(_06290_));
 sky130_fd_sc_hd__xnor2_1 _13225_ (.A(_06086_),
    .B(_06290_),
    .Y(_06292_));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(net576),
    .A1(_06292_),
    .S(net2),
    .X(_06293_));
 sky130_fd_sc_hd__a22o_1 _13227_ (.A1(net578),
    .A2(net223),
    .B1(_06293_),
    .B2(net280),
    .X(_06294_));
 sky130_fd_sc_hd__and2_1 _13228_ (.A(net298),
    .B(_06294_),
    .X(_00127_));
 sky130_fd_sc_hd__xnor2_1 _13229_ (.A(_05983_),
    .B(_06088_),
    .Y(_06295_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(\div_shifter[61] ),
    .A1(_06295_),
    .S(net2),
    .X(_06296_));
 sky130_fd_sc_hd__a22o_1 _13231_ (.A1(net560),
    .A2(net223),
    .B1(_06296_),
    .B2(net280),
    .X(_06297_));
 sky130_fd_sc_hd__and2_1 _13232_ (.A(net298),
    .B(net561),
    .X(_00128_));
 sky130_fd_sc_hd__nand2b_1 _13233_ (.A_N(_06091_),
    .B(_06090_),
    .Y(_06298_));
 sky130_fd_sc_hd__a32o_1 _13234_ (.A1(net608),
    .A2(net280),
    .A3(_06298_),
    .B1(net223),
    .B2(net419),
    .X(_06299_));
 sky130_fd_sc_hd__and2_1 _13235_ (.A(net298),
    .B(net420),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _13236_ (.A(net373),
    .B(net218),
    .Y(_06301_));
 sky130_fd_sc_hd__o211a_1 _13237_ (.A1(net373),
    .A2(net279),
    .B1(net300),
    .C1(_06301_),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _13238_ (.A1(net607),
    .A2(net222),
    .B1(_05932_),
    .B2(net278),
    .X(_06302_));
 sky130_fd_sc_hd__o211a_1 _13239_ (.A1(net482),
    .A2(net373),
    .B1(net300),
    .C1(_06302_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _13240_ (.A1(net476),
    .A2(net222),
    .B1(_05933_),
    .B2(net278),
    .X(_06303_));
 sky130_fd_sc_hd__a21o_1 _13241_ (.A1(net482),
    .A2(net373),
    .B1(net476),
    .X(_06304_));
 sky130_fd_sc_hd__and3_1 _13242_ (.A(net302),
    .B(net610),
    .C(net483),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _13243_ (.A1(net411),
    .A2(net222),
    .B1(_05936_),
    .B2(net278),
    .X(_06305_));
 sky130_fd_sc_hd__a31o_1 _13244_ (.A1(\div_counter[2] ),
    .A2(\div_counter[1] ),
    .A3(net373),
    .B1(net411),
    .X(_06306_));
 sky130_fd_sc_hd__and3_1 _13245_ (.A(net301),
    .B(_06305_),
    .C(net412),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13246_ (.A1(net363),
    .A2(net222),
    .B1(_05937_),
    .B2(net279),
    .X(_06308_));
 sky130_fd_sc_hd__o211a_1 _13247_ (.A1(net363),
    .A2(_05935_),
    .B1(_06308_),
    .C1(net302),
    .X(_00134_));
 sky130_fd_sc_hd__o21a_1 _13248_ (.A1(net470),
    .A2(_05938_),
    .B1(net302),
    .X(_00135_));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00000_),
    .Q(busy_l));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00001_),
    .Q(divi1_sign));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net370),
    .Q(\divi2_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00003_),
    .Q(\divi2_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net338),
    .Q(\divi2_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00005_),
    .Q(\divi2_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net360),
    .Q(\divi2_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net346),
    .Q(\divi2_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00008_),
    .Q(\divi2_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net362),
    .Q(\divi2_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net366),
    .Q(\divi2_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net318),
    .Q(\divi2_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net344),
    .Q(\divi2_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net348),
    .Q(\divi2_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net356),
    .Q(\divi2_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net354),
    .Q(\divi2_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net334),
    .Q(\divi2_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net324),
    .Q(\divi2_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net328),
    .Q(\divi2_l[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net336),
    .Q(\divi2_l[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net358),
    .Q(\divi2_l[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net332),
    .Q(\divi2_l[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net326),
    .Q(\divi2_l[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net320),
    .Q(\divi2_l[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net314),
    .Q(\divi2_l[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13274_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net312),
    .Q(\divi2_l[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net330),
    .Q(\divi2_l[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net352),
    .Q(\divi2_l[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net340),
    .Q(\divi2_l[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net350),
    .Q(\divi2_l[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00030_),
    .Q(\divi2_l[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net342),
    .Q(\divi2_l[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net322),
    .Q(\divi2_l[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00033_),
    .Q(\divi2_l[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00034_),
    .Q(\div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00035_),
    .Q(\div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00036_),
    .Q(\div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net509),
    .Q(\div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00038_),
    .Q(\div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00039_),
    .Q(\div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00040_),
    .Q(\div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net469),
    .Q(\div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net532),
    .Q(\div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00043_),
    .Q(\div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00044_),
    .Q(\div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00045_),
    .Q(\div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net501),
    .Q(\div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net524),
    .Q(\div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00048_),
    .Q(\div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00049_),
    .Q(\div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00050_),
    .Q(\div_res[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net486),
    .Q(\div_res[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net512),
    .Q(\div_res[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net489),
    .Q(\div_res[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00054_),
    .Q(\div_res[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00055_),
    .Q(\div_res[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net537),
    .Q(\div_res[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net504),
    .Q(\div_res[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00058_),
    .Q(\div_res[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net519),
    .Q(\div_res[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net492),
    .Q(\div_res[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00061_),
    .Q(\div_res[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00062_),
    .Q(\div_res[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net481),
    .Q(\div_res[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net527),
    .Q(\div_res[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net430),
    .Q(\div_res[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00066_),
    .Q(\div_shifter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00067_),
    .Q(\div_shifter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net416),
    .Q(\div_shifter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net368),
    .Q(\div_shifter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00070_),
    .Q(\div_shifter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13320_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net316),
    .Q(\div_shifter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00072_),
    .Q(\div_shifter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00073_),
    .Q(\div_shifter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net457),
    .Q(\div_shifter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net454),
    .Q(\div_shifter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13325_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00076_),
    .Q(\div_shifter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13326_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net446),
    .Q(\div_shifter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13327_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00078_),
    .Q(\div_shifter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13328_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net464),
    .Q(\div_shifter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13329_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00080_),
    .Q(\div_shifter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00081_),
    .Q(\div_shifter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net388),
    .Q(\div_shifter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net449),
    .Q(\div_shifter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net404),
    .Q(\div_shifter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13334_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00085_),
    .Q(\div_shifter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00086_),
    .Q(\div_shifter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net435),
    .Q(\div_shifter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13337_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00088_),
    .Q(\div_shifter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13338_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00089_),
    .Q(\div_shifter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00090_),
    .Q(\div_shifter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13340_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00091_),
    .Q(\div_shifter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net379),
    .Q(\div_shifter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net425),
    .Q(\div_shifter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00094_),
    .Q(\div_shifter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net385),
    .Q(\div_shifter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net395),
    .Q(\div_shifter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net381),
    .Q(\div_shifter[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13347_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00098_),
    .Q(\div_shifter[32] ));
 sky130_fd_sc_hd__dfxtp_2 _13348_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00099_),
    .Q(\div_shifter[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00100_),
    .Q(\div_shifter[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00101_),
    .Q(\div_shifter[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00102_),
    .Q(\div_shifter[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00103_),
    .Q(\div_shifter[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00104_),
    .Q(\div_shifter[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00105_),
    .Q(\div_shifter[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00106_),
    .Q(\div_shifter[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00107_),
    .Q(\div_shifter[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00108_),
    .Q(\div_shifter[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00109_),
    .Q(\div_shifter[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00110_),
    .Q(\div_shifter[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00111_),
    .Q(\div_shifter[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13361_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00112_),
    .Q(\div_shifter[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00113_),
    .Q(\div_shifter[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00114_),
    .Q(\div_shifter[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00115_),
    .Q(\div_shifter[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00116_),
    .Q(\div_shifter[50] ));
 sky130_fd_sc_hd__dfxtp_2 _13366_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00117_),
    .Q(\div_shifter[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00118_),
    .Q(\div_shifter[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00119_),
    .Q(\div_shifter[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13369_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00120_),
    .Q(\div_shifter[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00121_),
    .Q(\div_shifter[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00122_),
    .Q(\div_shifter[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00123_),
    .Q(\div_shifter[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13373_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00124_),
    .Q(\div_shifter[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00125_),
    .Q(\div_shifter[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00126_),
    .Q(\div_shifter[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13376_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00127_),
    .Q(\div_shifter[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13377_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00128_),
    .Q(\div_shifter[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13378_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00129_),
    .Q(\div_shifter[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13379_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net376),
    .Q(\div_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13380_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net374),
    .Q(\div_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13381_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00132_),
    .Q(\div_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13382_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net413),
    .Q(\div_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net364),
    .Q(\div_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net471),
    .Q(div_complete));
 sky130_fd_sc_hd__buf_12 _13385_ (.A(instruction[11]),
    .X(loadstore_dest[0]));
 sky130_fd_sc_hd__buf_12 _13386_ (.A(instruction[12]),
    .X(loadstore_dest[1]));
 sky130_fd_sc_hd__buf_12 _13387_ (.A(instruction[13]),
    .X(loadstore_dest[2]));
 sky130_fd_sc_hd__buf_12 _13388_ (.A(instruction[14]),
    .X(loadstore_dest[3]));
 sky130_fd_sc_hd__buf_12 _13389_ (.A(instruction[15]),
    .X(loadstore_dest[4]));
 sky130_fd_sc_hd__buf_12 _13390_ (.A(instruction[5]),
    .X(loadstore_size[0]));
 sky130_fd_sc_hd__buf_12 _13391_ (.A(instruction[6]),
    .X(loadstore_size[1]));
 sky130_fd_sc_hd__buf_12 _13392_ (.A(instruction[8]),
    .X(pred_idx[0]));
 sky130_fd_sc_hd__buf_12 _13393_ (.A(instruction[9]),
    .X(pred_idx[1]));
 sky130_fd_sc_hd__buf_12 _13394_ (.A(instruction[10]),
    .X(pred_idx[2]));
 sky130_fd_sc_hd__buf_12 _13395_ (.A(instruction[4]),
    .X(sign_extend));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_16 fanout101 (.A(_00152_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_16 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_12 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_16 fanout104 (.A(_06549_),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(net107),
    .X(net105));
 sky130_fd_sc_hd__buf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_06543_),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_8 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_4 fanout11 (.A(_00457_),
    .X(net11));
 sky130_fd_sc_hd__buf_8 fanout110 (.A(_06530_),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_16 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_16 fanout112 (.A(_06523_),
    .X(net112));
 sky130_fd_sc_hd__buf_6 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 fanout114 (.A(_06509_),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(_06507_),
    .X(net116));
 sky130_fd_sc_hd__buf_6 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_6 fanout118 (.A(_06502_),
    .X(net118));
 sky130_fd_sc_hd__buf_6 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_8 fanout12 (.A(net14),
    .X(net12));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(_06494_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_8 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_6 fanout122 (.A(_06492_),
    .X(net122));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_8 fanout124 (.A(_06491_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_8 fanout126 (.A(_06476_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_8 fanout128 (.A(_00313_),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_4 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__buf_8 fanout130 (.A(_00309_),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_8 fanout132 (.A(_00280_),
    .X(net132));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_8 fanout134 (.A(_00256_),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_8 fanout135 (.A(_00191_),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(_00191_),
    .X(net136));
 sky130_fd_sc_hd__buf_6 fanout137 (.A(_00186_),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(_00186_),
    .X(net138));
 sky130_fd_sc_hd__buf_6 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout14 (.A(_00436_),
    .X(net14));
 sky130_fd_sc_hd__buf_8 fanout140 (.A(_00180_),
    .X(net140));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_8 fanout142 (.A(_00171_),
    .X(net142));
 sky130_fd_sc_hd__buf_6 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(_00142_),
    .X(net144));
 sky130_fd_sc_hd__buf_6 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_8 fanout146 (.A(_06557_),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(_06547_),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_16 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_6 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__buf_12 fanout150 (.A(_06500_),
    .X(net150));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_8 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_12 fanout154 (.A(_06467_),
    .X(net154));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_2 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(_02071_),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_8 fanout16 (.A(_00353_),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(_02070_),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(_02070_),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(_02070_),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_16 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_16 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_8 fanout168 (.A(_00290_),
    .X(net168));
 sky130_fd_sc_hd__buf_8 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout17 (.A(net19),
    .X(net17));
 sky130_fd_sc_hd__buf_8 fanout170 (.A(_00283_),
    .X(net170));
 sky130_fd_sc_hd__buf_6 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_8 fanout172 (.A(_00258_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_8 fanout173 (.A(net175),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(_00230_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_00219_),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(_06564_),
    .X(net180));
 sky130_fd_sc_hd__buf_8 fanout181 (.A(net183),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(_06537_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_8 fanout185 (.A(_06527_),
    .X(net185));
 sky130_fd_sc_hd__buf_12 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_12 fanout187 (.A(_06469_),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(_02244_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(_02175_),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(_00245_),
    .X(net19));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(_02175_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(_02174_),
    .X(net192));
 sky130_fd_sc_hd__buf_12 fanout193 (.A(net195),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_16 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_8 fanout195 (.A(_00274_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(_06477_),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(_05940_),
    .X(net197));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(_05940_),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(_05939_),
    .X(net199));
 sky130_fd_sc_hd__buf_6 fanout2 (.A(_06092_),
    .X(net2));
 sky130_fd_sc_hd__buf_6 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(_05939_),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net203),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(_05939_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_02261_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(_02261_),
    .X(net205));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(_02256_),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(_02246_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(_02246_),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(_02172_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 fanout21 (.A(_00190_),
    .X(net21));
 sky130_fd_sc_hd__buf_12 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(_00250_),
    .X(net211));
 sky130_fd_sc_hd__buf_12 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_12 fanout213 (.A(_00211_),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout215 (.A(_06460_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_8 fanout216 (.A(_06446_),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(_06433_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(_06433_),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__buf_8 fanout22 (.A(_00178_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(_06432_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_8 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(_06432_),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_8 fanout224 (.A(_06351_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(net229),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net229),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(_06350_),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_8 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_6 fanout230 (.A(_06345_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_8 fanout232 (.A(_06344_),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 fanout233 (.A(_06338_),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(_06338_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_8 fanout235 (.A(_06337_),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(_06331_),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(_06324_),
    .X(net239));
 sky130_fd_sc_hd__buf_6 fanout24 (.A(_00139_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_2 fanout242 (.A(_06323_),
    .X(net242));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(_06315_),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(_04665_),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(_02445_),
    .X(net246));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(net249),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(_02445_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_8 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(_02259_),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(_02253_),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(_02250_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 fanout254 (.A(_02250_),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(_02248_),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_8 fanout257 (.A(_00240_),
    .X(net257));
 sky130_fd_sc_hd__buf_12 fanout258 (.A(net260),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 fanout26 (.A(_06554_),
    .X(net26));
 sky130_fd_sc_hd__buf_12 fanout260 (.A(_00214_),
    .X(net260));
 sky130_fd_sc_hd__buf_6 fanout262 (.A(net266),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(net266),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 fanout264 (.A(net266),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_16 fanout266 (.A(_06425_),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_16 fanout267 (.A(_06424_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_8 fanout268 (.A(_06314_),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(_06314_),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(net272),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(_04644_),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(_04406_),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net277),
    .X(net275));
 sky130_fd_sc_hd__buf_2 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(net375),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_6 fanout28 (.A(_06538_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_8 fanout280 (.A(net375),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_8 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_8 fanout282 (.A(_06461_),
    .X(net282));
 sky130_fd_sc_hd__buf_8 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_4 fanout284 (.A(_04567_),
    .X(net284));
 sky130_fd_sc_hd__buf_8 fanout285 (.A(_04567_),
    .X(net285));
 sky130_fd_sc_hd__buf_8 fanout286 (.A(_04567_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_8 fanout287 (.A(_04556_),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(_04556_),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_8 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_4 fanout291 (.A(_04535_),
    .X(net291));
 sky130_fd_sc_hd__buf_6 fanout292 (.A(_04524_),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 fanout294 (.A(_04471_),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_2 fanout296 (.A(_04471_),
    .X(net296));
 sky130_fd_sc_hd__buf_4 fanout297 (.A(net302),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(net302),
    .X(net298));
 sky130_fd_sc_hd__buf_4 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(_06535_),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(net302),
    .X(net300));
 sky130_fd_sc_hd__buf_4 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__buf_2 fanout302 (.A(_04471_),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_8 fanout303 (.A(_04460_),
    .X(net303));
 sky130_fd_sc_hd__buf_4 fanout304 (.A(_04460_),
    .X(net304));
 sky130_fd_sc_hd__buf_6 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_8 fanout306 (.A(_04428_),
    .X(net306));
 sky130_fd_sc_hd__buf_8 fanout307 (.A(reg1_val[1]),
    .X(net307));
 sky130_fd_sc_hd__buf_8 fanout308 (.A(reg1_val[0]),
    .X(net308));
 sky130_fd_sc_hd__buf_6 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(_00596_),
    .X(net31));
 sky130_fd_sc_hd__buf_8 fanout310 (.A(instruction[7]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_8 fanout32 (.A(_00596_),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_8 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__buf_8 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_8 fanout35 (.A(_00595_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_8 fanout37 (.A(_00354_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_8 fanout4 (.A(net5),
    .X(net4));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(_00317_),
    .X(net40));
 sky130_fd_sc_hd__buf_6 fanout41 (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_8 fanout43 (.A(_00312_),
    .X(net43));
 sky130_fd_sc_hd__buf_6 fanout44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__buf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_8 fanout46 (.A(_00285_),
    .X(net46));
 sky130_fd_sc_hd__buf_6 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_8 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 fanout49 (.A(_00282_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout5 (.A(_00601_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout52 (.A(_00260_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 fanout53 (.A(net55),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(_00257_),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__buf_6 fanout57 (.A(_00241_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_8 fanout6 (.A(net8),
    .X(net6));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(_00236_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 fanout63 (.A(_00229_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_6 fanout65 (.A(_00192_),
    .X(net65));
 sky130_fd_sc_hd__buf_6 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_6 fanout67 (.A(_00181_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(_00163_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_8 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_8 fanout71 (.A(_00143_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 fanout73 (.A(_06558_),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(_06506_),
    .X(net75));
 sky130_fd_sc_hd__buf_8 fanout76 (.A(net78),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(_00347_),
    .X(net78));
 sky130_fd_sc_hd__buf_6 fanout79 (.A(net81),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout8 (.A(_00511_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_8 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(_00301_),
    .X(net81));
 sky130_fd_sc_hd__buf_6 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_8 fanout83 (.A(_00299_),
    .X(net83));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(net86),
    .X(net84));
 sky130_fd_sc_hd__buf_4 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(_00298_),
    .X(net86));
 sky130_fd_sc_hd__buf_6 fanout87 (.A(_00295_),
    .X(net87));
 sky130_fd_sc_hd__buf_6 fanout88 (.A(_00295_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_8 fanout89 (.A(_00269_),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout9 (.A(net11),
    .X(net9));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(_00269_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_16 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(_00174_),
    .X(net92));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(_00174_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(_00167_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_8 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_8 fanout97 (.A(_00166_),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_8 fanout99 (.A(_00158_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\divi2_l[23] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00023_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_06154_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\div_counter[3] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_06306_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_00133_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net421),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_06134_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_00068_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\div_shifter[23] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_06160_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\div_shifter[63] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\divi2_l[30] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_06299_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\div_shifter[1] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_06133_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net438),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_06164_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00093_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net436),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_06159_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\div_res[31] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_06130_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00032_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_00065_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\div_shifter[14] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_06149_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\div_shifter[21] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_06157_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_00087_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\div_shifter[22] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_06158_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\div_shifter[27] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_06165_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\divi2_l[15] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\div_shifter[20] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_06155_),
    .X(net441));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold132 (.A(\divi2_l[1] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_05944_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\div_shifter[11] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_06145_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_00077_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\div_shifter[17] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_06152_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_00083_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00017_),
    .X(net324));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold140 (.A(\divi2_l[28] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_05976_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\div_shifter[9] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_06142_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_00075_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\div_shifter[8] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_06141_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_00074_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\div_shifter[6] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_06139_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\divi2_l[20] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\div_shifter[10] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_06143_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(net472),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_06147_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_00079_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\div_shifter[7] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_06140_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\div_res[6] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_06101_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_00041_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00022_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(div_complete),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_00135_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\div_shifter[13] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_06148_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\div_shifter[12] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_06146_),
    .X(net475));
 sky130_fd_sc_hd__buf_1 hold166 (.A(net609),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_05935_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_05937_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\div_res[28] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\divi2_l[16] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_06128_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_00063_),
    .X(net481));
 sky130_fd_sc_hd__buf_1 hold172 (.A(\div_counter[1] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_06304_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\div_res[16] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_06113_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_00051_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\div_res[19] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_06116_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_00053_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_00018_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net533),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_06124_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_00060_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\div_res[15] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_06112_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\div_res[5] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_06100_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\div_res[4] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_06099_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\div_res[11] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\divi2_l[24] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_06107_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_00046_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\div_res[23] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_06121_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_00057_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\div_res[27] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_06127_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(net544),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_06097_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_00037_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00025_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00026_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\div_res[18] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_06115_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00052_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\div_res[10] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_06106_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net538),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_06111_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\div_res[25] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_06123_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_00059_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\divi2_l[19] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\div_res[20] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_06117_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\div_res[13] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_06109_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_00047_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\div_res[30] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_06129_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_00064_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\div_res[24] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_06122_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_00021_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\div_res[8] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_06103_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_00042_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\div_res[26] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_06125_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\div_res[22] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_06119_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_00056_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\div_res[14] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_06110_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\divi2_l[14] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(net542),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_06105_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\div_res[9] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_06104_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\div_res[3] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_06098_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\div_res[21] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_06118_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\div_res[2] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_06095_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_00016_),
    .X(net334));
 sky130_fd_sc_hd__buf_1 hold240 (.A(\div_shifter[34] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_06180_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\div_shifter[38] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_06196_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\div_shifter[33] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_06175_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\div_shifter[54] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_06266_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\div_res[1] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_06094_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\divi2_l[17] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\div_shifter[62] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_06297_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\div_shifter[53] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_06262_),
    .X(net563));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold254 (.A(\div_shifter[56] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_06273_),
    .X(net565));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold256 (.A(\div_shifter[59] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_06286_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\div_shifter[37] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_06191_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_00019_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\div_shifter[32] ),
    .X(net570));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold261 (.A(\div_shifter[57] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_06278_),
    .X(net572));
 sky130_fd_sc_hd__buf_1 hold263 (.A(\div_shifter[50] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_06250_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\div_shifter[55] ),
    .X(net575));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold266 (.A(\div_shifter[60] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_06289_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\div_shifter[61] ),
    .X(net578));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold269 (.A(\div_shifter[42] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\divi2_l[2] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_06214_),
    .X(net580));
 sky130_fd_sc_hd__buf_1 hold271 (.A(\div_shifter[47] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_06236_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\div_shifter[40] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_06205_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\div_shifter[52] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_06258_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\div_shifter[49] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_06245_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\div_shifter[46] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_00004_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_06232_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\div_shifter[58] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\div_shifter[45] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_06227_),
    .X(net593));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold284 (.A(\div_shifter[35] ),
    .X(net594));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold285 (.A(\div_shifter[43] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_06218_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\div_shifter[44] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\div_shifter[41] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_06209_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\divi2_l[26] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\div_res[0] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\div_shifter[36] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\div_shifter[48] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\div_shifter[51] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\div_shifter[39] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\div_shifter[30] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\div_shifter[2] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\div_counter[1] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\div_shifter[62] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\div_counter[2] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\divi2_l[22] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00028_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_06303_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\div_shifter[31] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_06170_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_06172_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\divi2_l[29] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_00031_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\divi2_l[10] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_00012_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\divi2_l[5] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_00007_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\divi2_l[11] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_00013_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\divi2_l[27] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00024_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_00029_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\divi2_l[25] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_00027_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\divi2_l[13] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_00015_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\divi2_l[12] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_00014_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\divi2_l[18] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_00020_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\divi2_l[4] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\div_shifter[5] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_00006_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\divi2_l[7] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_00009_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\div_counter[4] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_00134_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\divi2_l[8] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_00010_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\div_shifter[3] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_00069_),
    .X(net368));
 sky130_fd_sc_hd__buf_1 hold59 (.A(\divi2_l[0] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00071_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_00002_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(divi1_sign),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_05941_),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 hold63 (.A(\div_counter[0] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_00131_),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 hold65 (.A(busy_l),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_00130_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\div_shifter[25] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_06163_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_00092_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\divi2_l[9] ),
    .X(net317));
 sky130_fd_sc_hd__buf_1 hold70 (.A(net611),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_00097_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\div_shifter[28] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_04362_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_06166_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00095_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\div_shifter[15] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_06151_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_00082_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\div_shifter[4] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00011_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_04373_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_06136_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\div_shifter[29] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_04351_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_06167_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_00096_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\divi2_l[31] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_05980_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\divi2_l[3] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_05946_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\divi2_l[21] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\divi2_l[6] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_05950_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\div_shifter[18] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_06153_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00084_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\div_shifter[0] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_06131_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\div_shifter[24] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_06161_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\div_shifter[19] ),
    .X(net409));
 sky130_fd_sc_hd__buf_6 load_slew214 (.A(_00210_),
    .X(net214));
 sky130_fd_sc_hd__buf_6 max_cap151 (.A(_06499_),
    .X(net151));
 sky130_fd_sc_hd__buf_4 max_cap238 (.A(_06330_),
    .X(net238));
 sky130_fd_sc_hd__buf_6 max_cap261 (.A(_00213_),
    .X(net261));
 sky130_fd_sc_hd__buf_1 wire3 (.A(_02737_),
    .X(net3));
endmodule

