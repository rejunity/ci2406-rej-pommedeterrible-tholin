VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 1100.000 ;
  PIN cap_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END cap_addr[0]
  PIN cap_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END cap_addr[1]
  PIN cap_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END cap_addr[2]
  PIN cap_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END cap_addr[3]
  PIN cap_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END cap_addr[4]
  PIN cap_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END cap_addr[5]
  PIN cap_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END cap_addr[6]
  PIN cap_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END cap_addr[7]
  PIN cap_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END cap_addr[8]
  PIN cap_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 15.270 1096.000 15.550 1100.000 ;
    END
  END cap_io_in[0]
  PIN cap_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 1096.000 19.230 1100.000 ;
    END
  END cap_io_in[1]
  PIN cap_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 1096.000 22.910 1100.000 ;
    END
  END cap_io_in[2]
  PIN cap_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 26.310 1096.000 26.590 1100.000 ;
    END
  END cap_io_in[3]
  PIN cap_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 29.990 1096.000 30.270 1100.000 ;
    END
  END cap_io_in[4]
  PIN cap_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 1096.000 33.950 1100.000 ;
    END
  END cap_io_in[5]
  PIN cap_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 37.350 1096.000 37.630 1100.000 ;
    END
  END cap_io_in[6]
  PIN cap_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 41.030 1096.000 41.310 1100.000 ;
    END
  END cap_io_in[7]
  PIN cap_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 44.710 1096.000 44.990 1100.000 ;
    END
  END cap_io_in[8]
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END custom_settings[9]
  PIN io_in_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 11.590 1096.000 11.870 1100.000 ;
    END
  END io_in_0
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END io_oeb[9]
  PIN io_oeb_6502
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 353.640 200.000 354.240 ;
    END
  END io_oeb_6502
  PIN io_oeb_8x305[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END io_oeb_8x305[0]
  PIN io_oeb_8x305[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END io_oeb_8x305[1]
  PIN io_oeb_8x305[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END io_oeb_8x305[2]
  PIN io_oeb_8x305[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END io_oeb_8x305[3]
  PIN io_oeb_8x305[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 995.560 4.000 996.160 ;
    END
  END io_oeb_8x305[4]
  PIN io_oeb_as1802
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 946.600 200.000 947.200 ;
    END
  END io_oeb_as1802
  PIN io_oeb_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END io_oeb_scrapcpu[0]
  PIN io_oeb_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END io_oeb_scrapcpu[10]
  PIN io_oeb_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END io_oeb_scrapcpu[11]
  PIN io_oeb_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END io_oeb_scrapcpu[12]
  PIN io_oeb_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END io_oeb_scrapcpu[13]
  PIN io_oeb_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END io_oeb_scrapcpu[14]
  PIN io_oeb_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END io_oeb_scrapcpu[15]
  PIN io_oeb_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END io_oeb_scrapcpu[16]
  PIN io_oeb_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END io_oeb_scrapcpu[17]
  PIN io_oeb_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END io_oeb_scrapcpu[18]
  PIN io_oeb_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END io_oeb_scrapcpu[19]
  PIN io_oeb_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END io_oeb_scrapcpu[1]
  PIN io_oeb_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END io_oeb_scrapcpu[20]
  PIN io_oeb_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END io_oeb_scrapcpu[21]
  PIN io_oeb_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END io_oeb_scrapcpu[22]
  PIN io_oeb_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END io_oeb_scrapcpu[23]
  PIN io_oeb_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END io_oeb_scrapcpu[24]
  PIN io_oeb_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END io_oeb_scrapcpu[25]
  PIN io_oeb_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END io_oeb_scrapcpu[26]
  PIN io_oeb_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_oeb_scrapcpu[27]
  PIN io_oeb_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END io_oeb_scrapcpu[28]
  PIN io_oeb_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END io_oeb_scrapcpu[29]
  PIN io_oeb_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io_oeb_scrapcpu[2]
  PIN io_oeb_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END io_oeb_scrapcpu[30]
  PIN io_oeb_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END io_oeb_scrapcpu[31]
  PIN io_oeb_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END io_oeb_scrapcpu[32]
  PIN io_oeb_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END io_oeb_scrapcpu[33]
  PIN io_oeb_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END io_oeb_scrapcpu[34]
  PIN io_oeb_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END io_oeb_scrapcpu[35]
  PIN io_oeb_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END io_oeb_scrapcpu[3]
  PIN io_oeb_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END io_oeb_scrapcpu[4]
  PIN io_oeb_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END io_oeb_scrapcpu[5]
  PIN io_oeb_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END io_oeb_scrapcpu[6]
  PIN io_oeb_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io_oeb_scrapcpu[7]
  PIN io_oeb_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END io_oeb_scrapcpu[8]
  PIN io_oeb_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END io_oeb_scrapcpu[9]
  PIN io_oeb_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END io_oeb_vliw[0]
  PIN io_oeb_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END io_oeb_vliw[10]
  PIN io_oeb_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END io_oeb_vliw[11]
  PIN io_oeb_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END io_oeb_vliw[12]
  PIN io_oeb_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END io_oeb_vliw[13]
  PIN io_oeb_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END io_oeb_vliw[14]
  PIN io_oeb_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END io_oeb_vliw[15]
  PIN io_oeb_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END io_oeb_vliw[16]
  PIN io_oeb_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END io_oeb_vliw[17]
  PIN io_oeb_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END io_oeb_vliw[18]
  PIN io_oeb_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END io_oeb_vliw[19]
  PIN io_oeb_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END io_oeb_vliw[1]
  PIN io_oeb_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END io_oeb_vliw[20]
  PIN io_oeb_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END io_oeb_vliw[21]
  PIN io_oeb_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END io_oeb_vliw[22]
  PIN io_oeb_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io_oeb_vliw[23]
  PIN io_oeb_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END io_oeb_vliw[24]
  PIN io_oeb_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END io_oeb_vliw[25]
  PIN io_oeb_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END io_oeb_vliw[26]
  PIN io_oeb_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END io_oeb_vliw[27]
  PIN io_oeb_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io_oeb_vliw[28]
  PIN io_oeb_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END io_oeb_vliw[29]
  PIN io_oeb_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END io_oeb_vliw[2]
  PIN io_oeb_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END io_oeb_vliw[30]
  PIN io_oeb_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END io_oeb_vliw[31]
  PIN io_oeb_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END io_oeb_vliw[32]
  PIN io_oeb_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END io_oeb_vliw[33]
  PIN io_oeb_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END io_oeb_vliw[34]
  PIN io_oeb_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END io_oeb_vliw[35]
  PIN io_oeb_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_oeb_vliw[3]
  PIN io_oeb_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END io_oeb_vliw[4]
  PIN io_oeb_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END io_oeb_vliw[5]
  PIN io_oeb_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END io_oeb_vliw[6]
  PIN io_oeb_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END io_oeb_vliw[7]
  PIN io_oeb_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END io_oeb_vliw[8]
  PIN io_oeb_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END io_oeb_vliw[9]
  PIN io_oeb_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 652.840 200.000 653.440 ;
    END
  END io_oeb_z80[0]
  PIN io_oeb_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 680.040 200.000 680.640 ;
    END
  END io_oeb_z80[10]
  PIN io_oeb_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 682.760 200.000 683.360 ;
    END
  END io_oeb_z80[11]
  PIN io_oeb_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 685.480 200.000 686.080 ;
    END
  END io_oeb_z80[12]
  PIN io_oeb_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 688.200 200.000 688.800 ;
    END
  END io_oeb_z80[13]
  PIN io_oeb_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 690.920 200.000 691.520 ;
    END
  END io_oeb_z80[14]
  PIN io_oeb_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 693.640 200.000 694.240 ;
    END
  END io_oeb_z80[15]
  PIN io_oeb_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 696.360 200.000 696.960 ;
    END
  END io_oeb_z80[16]
  PIN io_oeb_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 699.080 200.000 699.680 ;
    END
  END io_oeb_z80[17]
  PIN io_oeb_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 701.800 200.000 702.400 ;
    END
  END io_oeb_z80[18]
  PIN io_oeb_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 704.520 200.000 705.120 ;
    END
  END io_oeb_z80[19]
  PIN io_oeb_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 655.560 200.000 656.160 ;
    END
  END io_oeb_z80[1]
  PIN io_oeb_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 707.240 200.000 707.840 ;
    END
  END io_oeb_z80[20]
  PIN io_oeb_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 709.960 200.000 710.560 ;
    END
  END io_oeb_z80[21]
  PIN io_oeb_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 712.680 200.000 713.280 ;
    END
  END io_oeb_z80[22]
  PIN io_oeb_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 715.400 200.000 716.000 ;
    END
  END io_oeb_z80[23]
  PIN io_oeb_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 718.120 200.000 718.720 ;
    END
  END io_oeb_z80[24]
  PIN io_oeb_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 720.840 200.000 721.440 ;
    END
  END io_oeb_z80[25]
  PIN io_oeb_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 723.560 200.000 724.160 ;
    END
  END io_oeb_z80[26]
  PIN io_oeb_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 726.280 200.000 726.880 ;
    END
  END io_oeb_z80[27]
  PIN io_oeb_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 729.000 200.000 729.600 ;
    END
  END io_oeb_z80[28]
  PIN io_oeb_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 731.720 200.000 732.320 ;
    END
  END io_oeb_z80[29]
  PIN io_oeb_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 658.280 200.000 658.880 ;
    END
  END io_oeb_z80[2]
  PIN io_oeb_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 734.440 200.000 735.040 ;
    END
  END io_oeb_z80[30]
  PIN io_oeb_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 737.160 200.000 737.760 ;
    END
  END io_oeb_z80[31]
  PIN io_oeb_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 739.880 200.000 740.480 ;
    END
  END io_oeb_z80[32]
  PIN io_oeb_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 742.600 200.000 743.200 ;
    END
  END io_oeb_z80[33]
  PIN io_oeb_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 745.320 200.000 745.920 ;
    END
  END io_oeb_z80[34]
  PIN io_oeb_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 748.040 200.000 748.640 ;
    END
  END io_oeb_z80[35]
  PIN io_oeb_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 661.000 200.000 661.600 ;
    END
  END io_oeb_z80[3]
  PIN io_oeb_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 663.720 200.000 664.320 ;
    END
  END io_oeb_z80[4]
  PIN io_oeb_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 666.440 200.000 667.040 ;
    END
  END io_oeb_z80[5]
  PIN io_oeb_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 669.160 200.000 669.760 ;
    END
  END io_oeb_z80[6]
  PIN io_oeb_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 671.880 200.000 672.480 ;
    END
  END io_oeb_z80[7]
  PIN io_oeb_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 674.600 200.000 675.200 ;
    END
  END io_oeb_z80[8]
  PIN io_oeb_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 677.320 200.000 677.920 ;
    END
  END io_oeb_z80[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 200.000 152.960 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 200.000 180.160 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 182.280 200.000 182.880 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.000 200.000 185.600 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.720 200.000 188.320 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 200.000 191.040 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.160 200.000 193.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 195.880 200.000 196.480 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 198.600 200.000 199.200 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 201.320 200.000 201.920 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 204.040 200.000 204.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.080 200.000 155.680 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 206.760 200.000 207.360 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 209.480 200.000 210.080 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 212.200 200.000 212.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 214.920 200.000 215.520 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 217.640 200.000 218.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 220.360 200.000 220.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 223.080 200.000 223.680 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 225.800 200.000 226.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 228.520 200.000 229.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 231.240 200.000 231.840 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.800 200.000 158.400 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 233.960 200.000 234.560 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 236.680 200.000 237.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 239.400 200.000 240.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 242.120 200.000 242.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 244.840 200.000 245.440 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 247.560 200.000 248.160 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 250.280 200.000 250.880 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 253.000 200.000 253.600 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 160.520 200.000 161.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 200.000 163.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.960 200.000 166.560 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 171.400 200.000 172.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 174.120 200.000 174.720 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END io_out[9]
  PIN io_out_6502[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 255.720 200.000 256.320 ;
    END
  END io_out_6502[0]
  PIN io_out_6502[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.920 200.000 283.520 ;
    END
  END io_out_6502[10]
  PIN io_out_6502[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 285.640 200.000 286.240 ;
    END
  END io_out_6502[11]
  PIN io_out_6502[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 288.360 200.000 288.960 ;
    END
  END io_out_6502[12]
  PIN io_out_6502[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 291.080 200.000 291.680 ;
    END
  END io_out_6502[13]
  PIN io_out_6502[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 293.800 200.000 294.400 ;
    END
  END io_out_6502[14]
  PIN io_out_6502[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 296.520 200.000 297.120 ;
    END
  END io_out_6502[15]
  PIN io_out_6502[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 299.240 200.000 299.840 ;
    END
  END io_out_6502[16]
  PIN io_out_6502[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 301.960 200.000 302.560 ;
    END
  END io_out_6502[17]
  PIN io_out_6502[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 304.680 200.000 305.280 ;
    END
  END io_out_6502[18]
  PIN io_out_6502[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 307.400 200.000 308.000 ;
    END
  END io_out_6502[19]
  PIN io_out_6502[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 258.440 200.000 259.040 ;
    END
  END io_out_6502[1]
  PIN io_out_6502[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 310.120 200.000 310.720 ;
    END
  END io_out_6502[20]
  PIN io_out_6502[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 312.840 200.000 313.440 ;
    END
  END io_out_6502[21]
  PIN io_out_6502[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 315.560 200.000 316.160 ;
    END
  END io_out_6502[22]
  PIN io_out_6502[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 318.280 200.000 318.880 ;
    END
  END io_out_6502[23]
  PIN io_out_6502[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 321.000 200.000 321.600 ;
    END
  END io_out_6502[24]
  PIN io_out_6502[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 323.720 200.000 324.320 ;
    END
  END io_out_6502[25]
  PIN io_out_6502[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 326.440 200.000 327.040 ;
    END
  END io_out_6502[26]
  PIN io_out_6502[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 329.160 200.000 329.760 ;
    END
  END io_out_6502[27]
  PIN io_out_6502[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 331.880 200.000 332.480 ;
    END
  END io_out_6502[28]
  PIN io_out_6502[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 334.600 200.000 335.200 ;
    END
  END io_out_6502[29]
  PIN io_out_6502[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 261.160 200.000 261.760 ;
    END
  END io_out_6502[2]
  PIN io_out_6502[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 337.320 200.000 337.920 ;
    END
  END io_out_6502[30]
  PIN io_out_6502[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 340.040 200.000 340.640 ;
    END
  END io_out_6502[31]
  PIN io_out_6502[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 342.760 200.000 343.360 ;
    END
  END io_out_6502[32]
  PIN io_out_6502[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 345.480 200.000 346.080 ;
    END
  END io_out_6502[33]
  PIN io_out_6502[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 348.200 200.000 348.800 ;
    END
  END io_out_6502[34]
  PIN io_out_6502[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 350.920 200.000 351.520 ;
    END
  END io_out_6502[35]
  PIN io_out_6502[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 263.880 200.000 264.480 ;
    END
  END io_out_6502[3]
  PIN io_out_6502[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 266.600 200.000 267.200 ;
    END
  END io_out_6502[4]
  PIN io_out_6502[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 269.320 200.000 269.920 ;
    END
  END io_out_6502[5]
  PIN io_out_6502[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 272.040 200.000 272.640 ;
    END
  END io_out_6502[6]
  PIN io_out_6502[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 274.760 200.000 275.360 ;
    END
  END io_out_6502[7]
  PIN io_out_6502[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 277.480 200.000 278.080 ;
    END
  END io_out_6502[8]
  PIN io_out_6502[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 280.200 200.000 280.800 ;
    END
  END io_out_6502[9]
  PIN io_out_8x305[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END io_out_8x305[0]
  PIN io_out_8x305[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END io_out_8x305[10]
  PIN io_out_8x305[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END io_out_8x305[11]
  PIN io_out_8x305[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END io_out_8x305[12]
  PIN io_out_8x305[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 4.000 886.000 ;
    END
  END io_out_8x305[13]
  PIN io_out_8x305[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END io_out_8x305[14]
  PIN io_out_8x305[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END io_out_8x305[15]
  PIN io_out_8x305[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END io_out_8x305[16]
  PIN io_out_8x305[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 4.000 902.320 ;
    END
  END io_out_8x305[17]
  PIN io_out_8x305[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END io_out_8x305[18]
  PIN io_out_8x305[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END io_out_8x305[19]
  PIN io_out_8x305[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END io_out_8x305[1]
  PIN io_out_8x305[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.960 4.000 914.560 ;
    END
  END io_out_8x305[20]
  PIN io_out_8x305[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END io_out_8x305[21]
  PIN io_out_8x305[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.120 4.000 922.720 ;
    END
  END io_out_8x305[22]
  PIN io_out_8x305[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 4.000 926.800 ;
    END
  END io_out_8x305[23]
  PIN io_out_8x305[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.280 4.000 930.880 ;
    END
  END io_out_8x305[24]
  PIN io_out_8x305[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END io_out_8x305[25]
  PIN io_out_8x305[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END io_out_8x305[26]
  PIN io_out_8x305[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 942.520 4.000 943.120 ;
    END
  END io_out_8x305[27]
  PIN io_out_8x305[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 946.600 4.000 947.200 ;
    END
  END io_out_8x305[28]
  PIN io_out_8x305[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END io_out_8x305[29]
  PIN io_out_8x305[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END io_out_8x305[2]
  PIN io_out_8x305[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END io_out_8x305[30]
  PIN io_out_8x305[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END io_out_8x305[31]
  PIN io_out_8x305[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.920 4.000 963.520 ;
    END
  END io_out_8x305[32]
  PIN io_out_8x305[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.000 4.000 967.600 ;
    END
  END io_out_8x305[33]
  PIN io_out_8x305[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END io_out_8x305[34]
  PIN io_out_8x305[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END io_out_8x305[35]
  PIN io_out_8x305[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END io_out_8x305[3]
  PIN io_out_8x305[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END io_out_8x305[4]
  PIN io_out_8x305[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END io_out_8x305[5]
  PIN io_out_8x305[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END io_out_8x305[6]
  PIN io_out_8x305[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END io_out_8x305[7]
  PIN io_out_8x305[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END io_out_8x305[8]
  PIN io_out_8x305[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.080 4.000 869.680 ;
    END
  END io_out_8x305[9]
  PIN io_out_as1802[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 848.680 200.000 849.280 ;
    END
  END io_out_as1802[0]
  PIN io_out_as1802[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 875.880 200.000 876.480 ;
    END
  END io_out_as1802[10]
  PIN io_out_as1802[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 878.600 200.000 879.200 ;
    END
  END io_out_as1802[11]
  PIN io_out_as1802[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 881.320 200.000 881.920 ;
    END
  END io_out_as1802[12]
  PIN io_out_as1802[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 884.040 200.000 884.640 ;
    END
  END io_out_as1802[13]
  PIN io_out_as1802[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 886.760 200.000 887.360 ;
    END
  END io_out_as1802[14]
  PIN io_out_as1802[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 889.480 200.000 890.080 ;
    END
  END io_out_as1802[15]
  PIN io_out_as1802[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 892.200 200.000 892.800 ;
    END
  END io_out_as1802[16]
  PIN io_out_as1802[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 894.920 200.000 895.520 ;
    END
  END io_out_as1802[17]
  PIN io_out_as1802[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 897.640 200.000 898.240 ;
    END
  END io_out_as1802[18]
  PIN io_out_as1802[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 900.360 200.000 900.960 ;
    END
  END io_out_as1802[19]
  PIN io_out_as1802[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 851.400 200.000 852.000 ;
    END
  END io_out_as1802[1]
  PIN io_out_as1802[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 903.080 200.000 903.680 ;
    END
  END io_out_as1802[20]
  PIN io_out_as1802[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 905.800 200.000 906.400 ;
    END
  END io_out_as1802[21]
  PIN io_out_as1802[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 908.520 200.000 909.120 ;
    END
  END io_out_as1802[22]
  PIN io_out_as1802[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 911.240 200.000 911.840 ;
    END
  END io_out_as1802[23]
  PIN io_out_as1802[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 913.960 200.000 914.560 ;
    END
  END io_out_as1802[24]
  PIN io_out_as1802[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 916.680 200.000 917.280 ;
    END
  END io_out_as1802[25]
  PIN io_out_as1802[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 919.400 200.000 920.000 ;
    END
  END io_out_as1802[26]
  PIN io_out_as1802[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 922.120 200.000 922.720 ;
    END
  END io_out_as1802[27]
  PIN io_out_as1802[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 924.840 200.000 925.440 ;
    END
  END io_out_as1802[28]
  PIN io_out_as1802[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 927.560 200.000 928.160 ;
    END
  END io_out_as1802[29]
  PIN io_out_as1802[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 854.120 200.000 854.720 ;
    END
  END io_out_as1802[2]
  PIN io_out_as1802[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 930.280 200.000 930.880 ;
    END
  END io_out_as1802[30]
  PIN io_out_as1802[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 933.000 200.000 933.600 ;
    END
  END io_out_as1802[31]
  PIN io_out_as1802[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 935.720 200.000 936.320 ;
    END
  END io_out_as1802[32]
  PIN io_out_as1802[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 938.440 200.000 939.040 ;
    END
  END io_out_as1802[33]
  PIN io_out_as1802[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 941.160 200.000 941.760 ;
    END
  END io_out_as1802[34]
  PIN io_out_as1802[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 943.880 200.000 944.480 ;
    END
  END io_out_as1802[35]
  PIN io_out_as1802[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 856.840 200.000 857.440 ;
    END
  END io_out_as1802[3]
  PIN io_out_as1802[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 859.560 200.000 860.160 ;
    END
  END io_out_as1802[4]
  PIN io_out_as1802[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 862.280 200.000 862.880 ;
    END
  END io_out_as1802[5]
  PIN io_out_as1802[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 865.000 200.000 865.600 ;
    END
  END io_out_as1802[6]
  PIN io_out_as1802[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 867.720 200.000 868.320 ;
    END
  END io_out_as1802[7]
  PIN io_out_as1802[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 870.440 200.000 871.040 ;
    END
  END io_out_as1802[8]
  PIN io_out_as1802[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 873.160 200.000 873.760 ;
    END
  END io_out_as1802[9]
  PIN io_out_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 750.760 200.000 751.360 ;
    END
  END io_out_scrapcpu[0]
  PIN io_out_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 777.960 200.000 778.560 ;
    END
  END io_out_scrapcpu[10]
  PIN io_out_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 780.680 200.000 781.280 ;
    END
  END io_out_scrapcpu[11]
  PIN io_out_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 783.400 200.000 784.000 ;
    END
  END io_out_scrapcpu[12]
  PIN io_out_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 786.120 200.000 786.720 ;
    END
  END io_out_scrapcpu[13]
  PIN io_out_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 788.840 200.000 789.440 ;
    END
  END io_out_scrapcpu[14]
  PIN io_out_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 791.560 200.000 792.160 ;
    END
  END io_out_scrapcpu[15]
  PIN io_out_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 794.280 200.000 794.880 ;
    END
  END io_out_scrapcpu[16]
  PIN io_out_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 797.000 200.000 797.600 ;
    END
  END io_out_scrapcpu[17]
  PIN io_out_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 799.720 200.000 800.320 ;
    END
  END io_out_scrapcpu[18]
  PIN io_out_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 802.440 200.000 803.040 ;
    END
  END io_out_scrapcpu[19]
  PIN io_out_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 753.480 200.000 754.080 ;
    END
  END io_out_scrapcpu[1]
  PIN io_out_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 805.160 200.000 805.760 ;
    END
  END io_out_scrapcpu[20]
  PIN io_out_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 807.880 200.000 808.480 ;
    END
  END io_out_scrapcpu[21]
  PIN io_out_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 810.600 200.000 811.200 ;
    END
  END io_out_scrapcpu[22]
  PIN io_out_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 813.320 200.000 813.920 ;
    END
  END io_out_scrapcpu[23]
  PIN io_out_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 816.040 200.000 816.640 ;
    END
  END io_out_scrapcpu[24]
  PIN io_out_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 818.760 200.000 819.360 ;
    END
  END io_out_scrapcpu[25]
  PIN io_out_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 821.480 200.000 822.080 ;
    END
  END io_out_scrapcpu[26]
  PIN io_out_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 824.200 200.000 824.800 ;
    END
  END io_out_scrapcpu[27]
  PIN io_out_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 826.920 200.000 827.520 ;
    END
  END io_out_scrapcpu[28]
  PIN io_out_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 829.640 200.000 830.240 ;
    END
  END io_out_scrapcpu[29]
  PIN io_out_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 756.200 200.000 756.800 ;
    END
  END io_out_scrapcpu[2]
  PIN io_out_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 832.360 200.000 832.960 ;
    END
  END io_out_scrapcpu[30]
  PIN io_out_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 835.080 200.000 835.680 ;
    END
  END io_out_scrapcpu[31]
  PIN io_out_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 837.800 200.000 838.400 ;
    END
  END io_out_scrapcpu[32]
  PIN io_out_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 840.520 200.000 841.120 ;
    END
  END io_out_scrapcpu[33]
  PIN io_out_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 843.240 200.000 843.840 ;
    END
  END io_out_scrapcpu[34]
  PIN io_out_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 845.960 200.000 846.560 ;
    END
  END io_out_scrapcpu[35]
  PIN io_out_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 758.920 200.000 759.520 ;
    END
  END io_out_scrapcpu[3]
  PIN io_out_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 761.640 200.000 762.240 ;
    END
  END io_out_scrapcpu[4]
  PIN io_out_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 764.360 200.000 764.960 ;
    END
  END io_out_scrapcpu[5]
  PIN io_out_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 767.080 200.000 767.680 ;
    END
  END io_out_scrapcpu[6]
  PIN io_out_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 769.800 200.000 770.400 ;
    END
  END io_out_scrapcpu[7]
  PIN io_out_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 772.520 200.000 773.120 ;
    END
  END io_out_scrapcpu[8]
  PIN io_out_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 775.240 200.000 775.840 ;
    END
  END io_out_scrapcpu[9]
  PIN io_out_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 1096.000 52.350 1100.000 ;
    END
  END io_out_vliw[0]
  PIN io_out_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 1096.000 89.150 1100.000 ;
    END
  END io_out_vliw[10]
  PIN io_out_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 1096.000 92.830 1100.000 ;
    END
  END io_out_vliw[11]
  PIN io_out_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 96.230 1096.000 96.510 1100.000 ;
    END
  END io_out_vliw[12]
  PIN io_out_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 1096.000 100.190 1100.000 ;
    END
  END io_out_vliw[13]
  PIN io_out_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 103.590 1096.000 103.870 1100.000 ;
    END
  END io_out_vliw[14]
  PIN io_out_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 1096.000 107.550 1100.000 ;
    END
  END io_out_vliw[15]
  PIN io_out_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 1096.000 111.230 1100.000 ;
    END
  END io_out_vliw[16]
  PIN io_out_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 114.630 1096.000 114.910 1100.000 ;
    END
  END io_out_vliw[17]
  PIN io_out_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 118.310 1096.000 118.590 1100.000 ;
    END
  END io_out_vliw[18]
  PIN io_out_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 121.990 1096.000 122.270 1100.000 ;
    END
  END io_out_vliw[19]
  PIN io_out_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 1096.000 56.030 1100.000 ;
    END
  END io_out_vliw[1]
  PIN io_out_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 1096.000 125.950 1100.000 ;
    END
  END io_out_vliw[20]
  PIN io_out_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 1096.000 129.630 1100.000 ;
    END
  END io_out_vliw[21]
  PIN io_out_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 133.030 1096.000 133.310 1100.000 ;
    END
  END io_out_vliw[22]
  PIN io_out_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 1096.000 136.990 1100.000 ;
    END
  END io_out_vliw[23]
  PIN io_out_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 140.390 1096.000 140.670 1100.000 ;
    END
  END io_out_vliw[24]
  PIN io_out_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.070 1096.000 144.350 1100.000 ;
    END
  END io_out_vliw[25]
  PIN io_out_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 147.750 1096.000 148.030 1100.000 ;
    END
  END io_out_vliw[26]
  PIN io_out_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 1096.000 151.710 1100.000 ;
    END
  END io_out_vliw[27]
  PIN io_out_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 155.110 1096.000 155.390 1100.000 ;
    END
  END io_out_vliw[28]
  PIN io_out_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 158.790 1096.000 159.070 1100.000 ;
    END
  END io_out_vliw[29]
  PIN io_out_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 1096.000 59.710 1100.000 ;
    END
  END io_out_vliw[2]
  PIN io_out_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 162.470 1096.000 162.750 1100.000 ;
    END
  END io_out_vliw[30]
  PIN io_out_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 166.150 1096.000 166.430 1100.000 ;
    END
  END io_out_vliw[31]
  PIN io_out_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 169.830 1096.000 170.110 1100.000 ;
    END
  END io_out_vliw[32]
  PIN io_out_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.510 1096.000 173.790 1100.000 ;
    END
  END io_out_vliw[33]
  PIN io_out_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 1096.000 177.470 1100.000 ;
    END
  END io_out_vliw[34]
  PIN io_out_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 180.870 1096.000 181.150 1100.000 ;
    END
  END io_out_vliw[35]
  PIN io_out_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 63.110 1096.000 63.390 1100.000 ;
    END
  END io_out_vliw[3]
  PIN io_out_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 66.790 1096.000 67.070 1100.000 ;
    END
  END io_out_vliw[4]
  PIN io_out_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 70.470 1096.000 70.750 1100.000 ;
    END
  END io_out_vliw[5]
  PIN io_out_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 1096.000 74.430 1100.000 ;
    END
  END io_out_vliw[6]
  PIN io_out_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 77.830 1096.000 78.110 1100.000 ;
    END
  END io_out_vliw[7]
  PIN io_out_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 1096.000 81.790 1100.000 ;
    END
  END io_out_vliw[8]
  PIN io_out_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 85.190 1096.000 85.470 1100.000 ;
    END
  END io_out_vliw[9]
  PIN io_out_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 552.200 200.000 552.800 ;
    END
  END io_out_z80[0]
  PIN io_out_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 579.400 200.000 580.000 ;
    END
  END io_out_z80[10]
  PIN io_out_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 582.120 200.000 582.720 ;
    END
  END io_out_z80[11]
  PIN io_out_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 584.840 200.000 585.440 ;
    END
  END io_out_z80[12]
  PIN io_out_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 587.560 200.000 588.160 ;
    END
  END io_out_z80[13]
  PIN io_out_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 590.280 200.000 590.880 ;
    END
  END io_out_z80[14]
  PIN io_out_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 593.000 200.000 593.600 ;
    END
  END io_out_z80[15]
  PIN io_out_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 595.720 200.000 596.320 ;
    END
  END io_out_z80[16]
  PIN io_out_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 598.440 200.000 599.040 ;
    END
  END io_out_z80[17]
  PIN io_out_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 601.160 200.000 601.760 ;
    END
  END io_out_z80[18]
  PIN io_out_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 603.880 200.000 604.480 ;
    END
  END io_out_z80[19]
  PIN io_out_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 554.920 200.000 555.520 ;
    END
  END io_out_z80[1]
  PIN io_out_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 606.600 200.000 607.200 ;
    END
  END io_out_z80[20]
  PIN io_out_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 609.320 200.000 609.920 ;
    END
  END io_out_z80[21]
  PIN io_out_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 612.040 200.000 612.640 ;
    END
  END io_out_z80[22]
  PIN io_out_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 614.760 200.000 615.360 ;
    END
  END io_out_z80[23]
  PIN io_out_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 617.480 200.000 618.080 ;
    END
  END io_out_z80[24]
  PIN io_out_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 620.200 200.000 620.800 ;
    END
  END io_out_z80[25]
  PIN io_out_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 622.920 200.000 623.520 ;
    END
  END io_out_z80[26]
  PIN io_out_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 625.640 200.000 626.240 ;
    END
  END io_out_z80[27]
  PIN io_out_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 628.360 200.000 628.960 ;
    END
  END io_out_z80[28]
  PIN io_out_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 631.080 200.000 631.680 ;
    END
  END io_out_z80[29]
  PIN io_out_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 557.640 200.000 558.240 ;
    END
  END io_out_z80[2]
  PIN io_out_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 633.800 200.000 634.400 ;
    END
  END io_out_z80[30]
  PIN io_out_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 636.520 200.000 637.120 ;
    END
  END io_out_z80[31]
  PIN io_out_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 639.240 200.000 639.840 ;
    END
  END io_out_z80[32]
  PIN io_out_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 641.960 200.000 642.560 ;
    END
  END io_out_z80[33]
  PIN io_out_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 644.680 200.000 645.280 ;
    END
  END io_out_z80[34]
  PIN io_out_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 647.400 200.000 648.000 ;
    END
  END io_out_z80[35]
  PIN io_out_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 560.360 200.000 560.960 ;
    END
  END io_out_z80[3]
  PIN io_out_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 563.080 200.000 563.680 ;
    END
  END io_out_z80[4]
  PIN io_out_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 565.800 200.000 566.400 ;
    END
  END io_out_z80[5]
  PIN io_out_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 568.520 200.000 569.120 ;
    END
  END io_out_z80[6]
  PIN io_out_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 571.240 200.000 571.840 ;
    END
  END io_out_z80[7]
  PIN io_out_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 573.960 200.000 574.560 ;
    END
  END io_out_z80[8]
  PIN io_out_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 576.680 200.000 577.280 ;
    END
  END io_out_z80[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 443.400 200.000 444.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 470.600 200.000 471.200 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 473.320 200.000 473.920 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 476.040 200.000 476.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 478.760 200.000 479.360 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 481.480 200.000 482.080 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 484.200 200.000 484.800 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 486.920 200.000 487.520 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 489.640 200.000 490.240 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 492.360 200.000 492.960 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 495.080 200.000 495.680 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 446.120 200.000 446.720 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 497.800 200.000 498.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 500.520 200.000 501.120 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 503.240 200.000 503.840 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 505.960 200.000 506.560 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 508.680 200.000 509.280 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 511.400 200.000 512.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 514.120 200.000 514.720 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 516.840 200.000 517.440 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 519.560 200.000 520.160 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 522.280 200.000 522.880 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 448.840 200.000 449.440 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 525.000 200.000 525.600 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 527.720 200.000 528.320 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 530.440 200.000 531.040 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 533.160 200.000 533.760 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.880 200.000 536.480 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 538.600 200.000 539.200 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 541.320 200.000 541.920 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 544.040 200.000 544.640 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 546.760 200.000 547.360 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 549.480 200.000 550.080 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 451.560 200.000 452.160 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 454.280 200.000 454.880 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 457.000 200.000 457.600 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 459.720 200.000 460.320 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 462.440 200.000 463.040 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 465.160 200.000 465.760 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 467.880 200.000 468.480 ;
    END
  END la_data_out[9]
  PIN rst_6502
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END rst_6502
  PIN rst_8x305
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END rst_8x305
  PIN rst_as1802
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 188.230 1096.000 188.510 1100.000 ;
    END
  END rst_as1802
  PIN rst_scrapcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 184.550 1096.000 184.830 1100.000 ;
    END
  END rst_scrapcpu
  PIN rst_vliw
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 1096.000 48.670 1100.000 ;
    END
  END rst_vliw
  PIN rst_z80
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 650.120 200.000 650.720 ;
    END
  END rst_z80
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 356.360 200.000 356.960 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 383.560 200.000 384.160 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 386.280 200.000 386.880 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 389.000 200.000 389.600 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 391.720 200.000 392.320 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 394.440 200.000 395.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 397.160 200.000 397.760 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 399.880 200.000 400.480 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 402.600 200.000 403.200 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 405.320 200.000 405.920 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 408.040 200.000 408.640 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 359.080 200.000 359.680 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 410.760 200.000 411.360 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 413.480 200.000 414.080 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 416.200 200.000 416.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 418.920 200.000 419.520 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 421.640 200.000 422.240 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 424.360 200.000 424.960 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 427.080 200.000 427.680 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 429.800 200.000 430.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 432.520 200.000 433.120 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 435.240 200.000 435.840 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 361.800 200.000 362.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 437.960 200.000 438.560 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 440.680 200.000 441.280 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 364.520 200.000 365.120 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 367.240 200.000 367.840 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 369.960 200.000 370.560 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 372.680 200.000 373.280 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 375.400 200.000 376.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 378.120 200.000 378.720 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 380.840 200.000 381.440 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 1088.085 ;
      LAYER met1 ;
        RECT 0.070 10.640 199.940 1088.240 ;
      LAYER met2 ;
        RECT 0.100 1095.720 11.310 1096.570 ;
        RECT 12.150 1095.720 14.990 1096.570 ;
        RECT 15.830 1095.720 18.670 1096.570 ;
        RECT 19.510 1095.720 22.350 1096.570 ;
        RECT 23.190 1095.720 26.030 1096.570 ;
        RECT 26.870 1095.720 29.710 1096.570 ;
        RECT 30.550 1095.720 33.390 1096.570 ;
        RECT 34.230 1095.720 37.070 1096.570 ;
        RECT 37.910 1095.720 40.750 1096.570 ;
        RECT 41.590 1095.720 44.430 1096.570 ;
        RECT 45.270 1095.720 48.110 1096.570 ;
        RECT 48.950 1095.720 51.790 1096.570 ;
        RECT 52.630 1095.720 55.470 1096.570 ;
        RECT 56.310 1095.720 59.150 1096.570 ;
        RECT 59.990 1095.720 62.830 1096.570 ;
        RECT 63.670 1095.720 66.510 1096.570 ;
        RECT 67.350 1095.720 70.190 1096.570 ;
        RECT 71.030 1095.720 73.870 1096.570 ;
        RECT 74.710 1095.720 77.550 1096.570 ;
        RECT 78.390 1095.720 81.230 1096.570 ;
        RECT 82.070 1095.720 84.910 1096.570 ;
        RECT 85.750 1095.720 88.590 1096.570 ;
        RECT 89.430 1095.720 92.270 1096.570 ;
        RECT 93.110 1095.720 95.950 1096.570 ;
        RECT 96.790 1095.720 99.630 1096.570 ;
        RECT 100.470 1095.720 103.310 1096.570 ;
        RECT 104.150 1095.720 106.990 1096.570 ;
        RECT 107.830 1095.720 110.670 1096.570 ;
        RECT 111.510 1095.720 114.350 1096.570 ;
        RECT 115.190 1095.720 118.030 1096.570 ;
        RECT 118.870 1095.720 121.710 1096.570 ;
        RECT 122.550 1095.720 125.390 1096.570 ;
        RECT 126.230 1095.720 129.070 1096.570 ;
        RECT 129.910 1095.720 132.750 1096.570 ;
        RECT 133.590 1095.720 136.430 1096.570 ;
        RECT 137.270 1095.720 140.110 1096.570 ;
        RECT 140.950 1095.720 143.790 1096.570 ;
        RECT 144.630 1095.720 147.470 1096.570 ;
        RECT 148.310 1095.720 151.150 1096.570 ;
        RECT 151.990 1095.720 154.830 1096.570 ;
        RECT 155.670 1095.720 158.510 1096.570 ;
        RECT 159.350 1095.720 162.190 1096.570 ;
        RECT 163.030 1095.720 165.870 1096.570 ;
        RECT 166.710 1095.720 169.550 1096.570 ;
        RECT 170.390 1095.720 173.230 1096.570 ;
        RECT 174.070 1095.720 176.910 1096.570 ;
        RECT 177.750 1095.720 180.590 1096.570 ;
        RECT 181.430 1095.720 184.270 1096.570 ;
        RECT 185.110 1095.720 187.950 1096.570 ;
        RECT 188.790 1095.720 199.940 1096.570 ;
        RECT 0.100 4.280 199.940 1095.720 ;
        RECT 0.100 4.000 5.330 4.280 ;
        RECT 6.170 4.000 9.930 4.280 ;
        RECT 10.770 4.000 14.530 4.280 ;
        RECT 15.370 4.000 19.130 4.280 ;
        RECT 19.970 4.000 23.730 4.280 ;
        RECT 24.570 4.000 28.330 4.280 ;
        RECT 29.170 4.000 32.930 4.280 ;
        RECT 33.770 4.000 37.530 4.280 ;
        RECT 38.370 4.000 42.130 4.280 ;
        RECT 42.970 4.000 46.730 4.280 ;
        RECT 47.570 4.000 51.330 4.280 ;
        RECT 52.170 4.000 55.930 4.280 ;
        RECT 56.770 4.000 60.530 4.280 ;
        RECT 61.370 4.000 65.130 4.280 ;
        RECT 65.970 4.000 69.730 4.280 ;
        RECT 70.570 4.000 74.330 4.280 ;
        RECT 75.170 4.000 78.930 4.280 ;
        RECT 79.770 4.000 83.530 4.280 ;
        RECT 84.370 4.000 88.130 4.280 ;
        RECT 88.970 4.000 92.730 4.280 ;
        RECT 93.570 4.000 97.330 4.280 ;
        RECT 98.170 4.000 101.930 4.280 ;
        RECT 102.770 4.000 106.530 4.280 ;
        RECT 107.370 4.000 111.130 4.280 ;
        RECT 111.970 4.000 115.730 4.280 ;
        RECT 116.570 4.000 120.330 4.280 ;
        RECT 121.170 4.000 124.930 4.280 ;
        RECT 125.770 4.000 129.530 4.280 ;
        RECT 130.370 4.000 134.130 4.280 ;
        RECT 134.970 4.000 138.730 4.280 ;
        RECT 139.570 4.000 143.330 4.280 ;
        RECT 144.170 4.000 147.930 4.280 ;
        RECT 148.770 4.000 152.530 4.280 ;
        RECT 153.370 4.000 157.130 4.280 ;
        RECT 157.970 4.000 161.730 4.280 ;
        RECT 162.570 4.000 166.330 4.280 ;
        RECT 167.170 4.000 170.930 4.280 ;
        RECT 171.770 4.000 175.530 4.280 ;
        RECT 176.370 4.000 180.130 4.280 ;
        RECT 180.970 4.000 184.730 4.280 ;
        RECT 185.570 4.000 189.330 4.280 ;
        RECT 190.170 4.000 193.930 4.280 ;
        RECT 194.770 4.000 199.940 4.280 ;
      LAYER met3 ;
        RECT 0.525 1000.640 196.000 1088.165 ;
        RECT 4.400 999.240 196.000 1000.640 ;
        RECT 0.525 996.560 196.000 999.240 ;
        RECT 4.400 995.160 196.000 996.560 ;
        RECT 0.525 992.480 196.000 995.160 ;
        RECT 4.400 991.080 196.000 992.480 ;
        RECT 0.525 988.400 196.000 991.080 ;
        RECT 4.400 987.000 196.000 988.400 ;
        RECT 0.525 984.320 196.000 987.000 ;
        RECT 4.400 982.920 196.000 984.320 ;
        RECT 0.525 980.240 196.000 982.920 ;
        RECT 4.400 978.840 196.000 980.240 ;
        RECT 0.525 976.160 196.000 978.840 ;
        RECT 4.400 974.760 196.000 976.160 ;
        RECT 0.525 972.080 196.000 974.760 ;
        RECT 4.400 970.680 196.000 972.080 ;
        RECT 0.525 968.000 196.000 970.680 ;
        RECT 4.400 966.600 196.000 968.000 ;
        RECT 0.525 963.920 196.000 966.600 ;
        RECT 4.400 962.520 196.000 963.920 ;
        RECT 0.525 959.840 196.000 962.520 ;
        RECT 4.400 958.440 196.000 959.840 ;
        RECT 0.525 955.760 196.000 958.440 ;
        RECT 4.400 954.360 196.000 955.760 ;
        RECT 0.525 951.680 196.000 954.360 ;
        RECT 4.400 950.280 196.000 951.680 ;
        RECT 0.525 947.600 196.000 950.280 ;
        RECT 4.400 946.200 195.600 947.600 ;
        RECT 0.525 944.880 196.000 946.200 ;
        RECT 0.525 943.520 195.600 944.880 ;
        RECT 4.400 943.480 195.600 943.520 ;
        RECT 4.400 942.160 196.000 943.480 ;
        RECT 4.400 942.120 195.600 942.160 ;
        RECT 0.525 940.760 195.600 942.120 ;
        RECT 0.525 939.440 196.000 940.760 ;
        RECT 4.400 938.040 195.600 939.440 ;
        RECT 0.525 936.720 196.000 938.040 ;
        RECT 0.525 935.360 195.600 936.720 ;
        RECT 4.400 935.320 195.600 935.360 ;
        RECT 4.400 934.000 196.000 935.320 ;
        RECT 4.400 933.960 195.600 934.000 ;
        RECT 0.525 932.600 195.600 933.960 ;
        RECT 0.525 931.280 196.000 932.600 ;
        RECT 4.400 929.880 195.600 931.280 ;
        RECT 0.525 928.560 196.000 929.880 ;
        RECT 0.525 927.200 195.600 928.560 ;
        RECT 4.400 927.160 195.600 927.200 ;
        RECT 4.400 925.840 196.000 927.160 ;
        RECT 4.400 925.800 195.600 925.840 ;
        RECT 0.525 924.440 195.600 925.800 ;
        RECT 0.525 923.120 196.000 924.440 ;
        RECT 4.400 921.720 195.600 923.120 ;
        RECT 0.525 920.400 196.000 921.720 ;
        RECT 0.525 919.040 195.600 920.400 ;
        RECT 4.400 919.000 195.600 919.040 ;
        RECT 4.400 917.680 196.000 919.000 ;
        RECT 4.400 917.640 195.600 917.680 ;
        RECT 0.525 916.280 195.600 917.640 ;
        RECT 0.525 914.960 196.000 916.280 ;
        RECT 4.400 913.560 195.600 914.960 ;
        RECT 0.525 912.240 196.000 913.560 ;
        RECT 0.525 910.880 195.600 912.240 ;
        RECT 4.400 910.840 195.600 910.880 ;
        RECT 4.400 909.520 196.000 910.840 ;
        RECT 4.400 909.480 195.600 909.520 ;
        RECT 0.525 908.120 195.600 909.480 ;
        RECT 0.525 906.800 196.000 908.120 ;
        RECT 4.400 905.400 195.600 906.800 ;
        RECT 0.525 904.080 196.000 905.400 ;
        RECT 0.525 902.720 195.600 904.080 ;
        RECT 4.400 902.680 195.600 902.720 ;
        RECT 4.400 901.360 196.000 902.680 ;
        RECT 4.400 901.320 195.600 901.360 ;
        RECT 0.525 899.960 195.600 901.320 ;
        RECT 0.525 898.640 196.000 899.960 ;
        RECT 4.400 897.240 195.600 898.640 ;
        RECT 0.525 895.920 196.000 897.240 ;
        RECT 0.525 894.560 195.600 895.920 ;
        RECT 4.400 894.520 195.600 894.560 ;
        RECT 4.400 893.200 196.000 894.520 ;
        RECT 4.400 893.160 195.600 893.200 ;
        RECT 0.525 891.800 195.600 893.160 ;
        RECT 0.525 890.480 196.000 891.800 ;
        RECT 4.400 889.080 195.600 890.480 ;
        RECT 0.525 887.760 196.000 889.080 ;
        RECT 0.525 886.400 195.600 887.760 ;
        RECT 4.400 886.360 195.600 886.400 ;
        RECT 4.400 885.040 196.000 886.360 ;
        RECT 4.400 885.000 195.600 885.040 ;
        RECT 0.525 883.640 195.600 885.000 ;
        RECT 0.525 882.320 196.000 883.640 ;
        RECT 4.400 880.920 195.600 882.320 ;
        RECT 0.525 879.600 196.000 880.920 ;
        RECT 0.525 878.240 195.600 879.600 ;
        RECT 4.400 878.200 195.600 878.240 ;
        RECT 4.400 876.880 196.000 878.200 ;
        RECT 4.400 876.840 195.600 876.880 ;
        RECT 0.525 875.480 195.600 876.840 ;
        RECT 0.525 874.160 196.000 875.480 ;
        RECT 4.400 872.760 195.600 874.160 ;
        RECT 0.525 871.440 196.000 872.760 ;
        RECT 0.525 870.080 195.600 871.440 ;
        RECT 4.400 870.040 195.600 870.080 ;
        RECT 4.400 868.720 196.000 870.040 ;
        RECT 4.400 868.680 195.600 868.720 ;
        RECT 0.525 867.320 195.600 868.680 ;
        RECT 0.525 866.000 196.000 867.320 ;
        RECT 4.400 864.600 195.600 866.000 ;
        RECT 0.525 863.280 196.000 864.600 ;
        RECT 0.525 861.920 195.600 863.280 ;
        RECT 4.400 861.880 195.600 861.920 ;
        RECT 4.400 860.560 196.000 861.880 ;
        RECT 4.400 860.520 195.600 860.560 ;
        RECT 0.525 859.160 195.600 860.520 ;
        RECT 0.525 857.840 196.000 859.160 ;
        RECT 4.400 856.440 195.600 857.840 ;
        RECT 0.525 855.120 196.000 856.440 ;
        RECT 0.525 853.760 195.600 855.120 ;
        RECT 4.400 853.720 195.600 853.760 ;
        RECT 4.400 852.400 196.000 853.720 ;
        RECT 4.400 852.360 195.600 852.400 ;
        RECT 0.525 851.000 195.600 852.360 ;
        RECT 0.525 849.680 196.000 851.000 ;
        RECT 4.400 848.280 195.600 849.680 ;
        RECT 0.525 846.960 196.000 848.280 ;
        RECT 0.525 845.600 195.600 846.960 ;
        RECT 4.400 845.560 195.600 845.600 ;
        RECT 4.400 844.240 196.000 845.560 ;
        RECT 4.400 844.200 195.600 844.240 ;
        RECT 0.525 842.840 195.600 844.200 ;
        RECT 0.525 841.520 196.000 842.840 ;
        RECT 4.400 840.120 195.600 841.520 ;
        RECT 0.525 838.800 196.000 840.120 ;
        RECT 0.525 837.440 195.600 838.800 ;
        RECT 4.400 837.400 195.600 837.440 ;
        RECT 4.400 836.080 196.000 837.400 ;
        RECT 4.400 836.040 195.600 836.080 ;
        RECT 0.525 834.680 195.600 836.040 ;
        RECT 0.525 833.360 196.000 834.680 ;
        RECT 4.400 831.960 195.600 833.360 ;
        RECT 0.525 830.640 196.000 831.960 ;
        RECT 0.525 829.280 195.600 830.640 ;
        RECT 4.400 829.240 195.600 829.280 ;
        RECT 4.400 827.920 196.000 829.240 ;
        RECT 4.400 827.880 195.600 827.920 ;
        RECT 0.525 826.520 195.600 827.880 ;
        RECT 0.525 825.200 196.000 826.520 ;
        RECT 4.400 823.800 195.600 825.200 ;
        RECT 0.525 822.480 196.000 823.800 ;
        RECT 0.525 821.120 195.600 822.480 ;
        RECT 4.400 821.080 195.600 821.120 ;
        RECT 4.400 819.760 196.000 821.080 ;
        RECT 4.400 819.720 195.600 819.760 ;
        RECT 0.525 818.360 195.600 819.720 ;
        RECT 0.525 817.040 196.000 818.360 ;
        RECT 4.400 815.640 195.600 817.040 ;
        RECT 0.525 814.320 196.000 815.640 ;
        RECT 0.525 812.960 195.600 814.320 ;
        RECT 4.400 812.920 195.600 812.960 ;
        RECT 4.400 811.600 196.000 812.920 ;
        RECT 4.400 811.560 195.600 811.600 ;
        RECT 0.525 810.200 195.600 811.560 ;
        RECT 0.525 808.880 196.000 810.200 ;
        RECT 4.400 807.480 195.600 808.880 ;
        RECT 0.525 806.160 196.000 807.480 ;
        RECT 0.525 804.800 195.600 806.160 ;
        RECT 4.400 804.760 195.600 804.800 ;
        RECT 4.400 803.440 196.000 804.760 ;
        RECT 4.400 803.400 195.600 803.440 ;
        RECT 0.525 802.040 195.600 803.400 ;
        RECT 0.525 800.720 196.000 802.040 ;
        RECT 4.400 799.320 195.600 800.720 ;
        RECT 0.525 798.000 196.000 799.320 ;
        RECT 0.525 796.640 195.600 798.000 ;
        RECT 4.400 796.600 195.600 796.640 ;
        RECT 4.400 795.280 196.000 796.600 ;
        RECT 4.400 795.240 195.600 795.280 ;
        RECT 0.525 793.880 195.600 795.240 ;
        RECT 0.525 792.560 196.000 793.880 ;
        RECT 4.400 791.160 195.600 792.560 ;
        RECT 0.525 789.840 196.000 791.160 ;
        RECT 0.525 788.480 195.600 789.840 ;
        RECT 4.400 788.440 195.600 788.480 ;
        RECT 4.400 787.120 196.000 788.440 ;
        RECT 4.400 787.080 195.600 787.120 ;
        RECT 0.525 785.720 195.600 787.080 ;
        RECT 0.525 784.400 196.000 785.720 ;
        RECT 4.400 783.000 195.600 784.400 ;
        RECT 0.525 781.680 196.000 783.000 ;
        RECT 0.525 780.320 195.600 781.680 ;
        RECT 4.400 780.280 195.600 780.320 ;
        RECT 4.400 778.960 196.000 780.280 ;
        RECT 4.400 778.920 195.600 778.960 ;
        RECT 0.525 777.560 195.600 778.920 ;
        RECT 0.525 776.240 196.000 777.560 ;
        RECT 4.400 774.840 195.600 776.240 ;
        RECT 0.525 773.520 196.000 774.840 ;
        RECT 0.525 772.160 195.600 773.520 ;
        RECT 4.400 772.120 195.600 772.160 ;
        RECT 4.400 770.800 196.000 772.120 ;
        RECT 4.400 770.760 195.600 770.800 ;
        RECT 0.525 769.400 195.600 770.760 ;
        RECT 0.525 768.080 196.000 769.400 ;
        RECT 4.400 766.680 195.600 768.080 ;
        RECT 0.525 765.360 196.000 766.680 ;
        RECT 0.525 764.000 195.600 765.360 ;
        RECT 4.400 763.960 195.600 764.000 ;
        RECT 4.400 762.640 196.000 763.960 ;
        RECT 4.400 762.600 195.600 762.640 ;
        RECT 0.525 761.240 195.600 762.600 ;
        RECT 0.525 759.920 196.000 761.240 ;
        RECT 4.400 758.520 195.600 759.920 ;
        RECT 0.525 757.200 196.000 758.520 ;
        RECT 0.525 755.840 195.600 757.200 ;
        RECT 4.400 755.800 195.600 755.840 ;
        RECT 4.400 754.480 196.000 755.800 ;
        RECT 4.400 754.440 195.600 754.480 ;
        RECT 0.525 753.080 195.600 754.440 ;
        RECT 0.525 751.760 196.000 753.080 ;
        RECT 4.400 750.360 195.600 751.760 ;
        RECT 0.525 749.040 196.000 750.360 ;
        RECT 0.525 747.680 195.600 749.040 ;
        RECT 4.400 747.640 195.600 747.680 ;
        RECT 4.400 746.320 196.000 747.640 ;
        RECT 4.400 746.280 195.600 746.320 ;
        RECT 0.525 744.920 195.600 746.280 ;
        RECT 0.525 743.600 196.000 744.920 ;
        RECT 4.400 742.200 195.600 743.600 ;
        RECT 0.525 740.880 196.000 742.200 ;
        RECT 0.525 739.520 195.600 740.880 ;
        RECT 4.400 739.480 195.600 739.520 ;
        RECT 4.400 738.160 196.000 739.480 ;
        RECT 4.400 738.120 195.600 738.160 ;
        RECT 0.525 736.760 195.600 738.120 ;
        RECT 0.525 735.440 196.000 736.760 ;
        RECT 4.400 734.040 195.600 735.440 ;
        RECT 0.525 732.720 196.000 734.040 ;
        RECT 0.525 731.360 195.600 732.720 ;
        RECT 4.400 731.320 195.600 731.360 ;
        RECT 4.400 730.000 196.000 731.320 ;
        RECT 4.400 729.960 195.600 730.000 ;
        RECT 0.525 728.600 195.600 729.960 ;
        RECT 0.525 727.280 196.000 728.600 ;
        RECT 4.400 725.880 195.600 727.280 ;
        RECT 0.525 724.560 196.000 725.880 ;
        RECT 0.525 723.200 195.600 724.560 ;
        RECT 4.400 723.160 195.600 723.200 ;
        RECT 4.400 721.840 196.000 723.160 ;
        RECT 4.400 721.800 195.600 721.840 ;
        RECT 0.525 720.440 195.600 721.800 ;
        RECT 0.525 719.120 196.000 720.440 ;
        RECT 4.400 717.720 195.600 719.120 ;
        RECT 0.525 716.400 196.000 717.720 ;
        RECT 0.525 715.040 195.600 716.400 ;
        RECT 4.400 715.000 195.600 715.040 ;
        RECT 4.400 713.680 196.000 715.000 ;
        RECT 4.400 713.640 195.600 713.680 ;
        RECT 0.525 712.280 195.600 713.640 ;
        RECT 0.525 710.960 196.000 712.280 ;
        RECT 4.400 709.560 195.600 710.960 ;
        RECT 0.525 708.240 196.000 709.560 ;
        RECT 0.525 706.880 195.600 708.240 ;
        RECT 4.400 706.840 195.600 706.880 ;
        RECT 4.400 705.520 196.000 706.840 ;
        RECT 4.400 705.480 195.600 705.520 ;
        RECT 0.525 704.120 195.600 705.480 ;
        RECT 0.525 702.800 196.000 704.120 ;
        RECT 4.400 701.400 195.600 702.800 ;
        RECT 0.525 700.080 196.000 701.400 ;
        RECT 0.525 698.720 195.600 700.080 ;
        RECT 4.400 698.680 195.600 698.720 ;
        RECT 4.400 697.360 196.000 698.680 ;
        RECT 4.400 697.320 195.600 697.360 ;
        RECT 0.525 695.960 195.600 697.320 ;
        RECT 0.525 694.640 196.000 695.960 ;
        RECT 4.400 693.240 195.600 694.640 ;
        RECT 0.525 691.920 196.000 693.240 ;
        RECT 0.525 690.560 195.600 691.920 ;
        RECT 4.400 690.520 195.600 690.560 ;
        RECT 4.400 689.200 196.000 690.520 ;
        RECT 4.400 689.160 195.600 689.200 ;
        RECT 0.525 687.800 195.600 689.160 ;
        RECT 0.525 686.480 196.000 687.800 ;
        RECT 4.400 685.080 195.600 686.480 ;
        RECT 0.525 683.760 196.000 685.080 ;
        RECT 0.525 682.400 195.600 683.760 ;
        RECT 4.400 682.360 195.600 682.400 ;
        RECT 4.400 681.040 196.000 682.360 ;
        RECT 4.400 681.000 195.600 681.040 ;
        RECT 0.525 679.640 195.600 681.000 ;
        RECT 0.525 678.320 196.000 679.640 ;
        RECT 4.400 676.920 195.600 678.320 ;
        RECT 0.525 675.600 196.000 676.920 ;
        RECT 0.525 674.240 195.600 675.600 ;
        RECT 4.400 674.200 195.600 674.240 ;
        RECT 4.400 672.880 196.000 674.200 ;
        RECT 4.400 672.840 195.600 672.880 ;
        RECT 0.525 671.480 195.600 672.840 ;
        RECT 0.525 670.160 196.000 671.480 ;
        RECT 4.400 668.760 195.600 670.160 ;
        RECT 0.525 667.440 196.000 668.760 ;
        RECT 0.525 666.080 195.600 667.440 ;
        RECT 4.400 666.040 195.600 666.080 ;
        RECT 4.400 664.720 196.000 666.040 ;
        RECT 4.400 664.680 195.600 664.720 ;
        RECT 0.525 663.320 195.600 664.680 ;
        RECT 0.525 662.000 196.000 663.320 ;
        RECT 4.400 660.600 195.600 662.000 ;
        RECT 0.525 659.280 196.000 660.600 ;
        RECT 0.525 657.920 195.600 659.280 ;
        RECT 4.400 657.880 195.600 657.920 ;
        RECT 4.400 656.560 196.000 657.880 ;
        RECT 4.400 656.520 195.600 656.560 ;
        RECT 0.525 655.160 195.600 656.520 ;
        RECT 0.525 653.840 196.000 655.160 ;
        RECT 4.400 652.440 195.600 653.840 ;
        RECT 0.525 651.120 196.000 652.440 ;
        RECT 0.525 649.760 195.600 651.120 ;
        RECT 4.400 649.720 195.600 649.760 ;
        RECT 4.400 648.400 196.000 649.720 ;
        RECT 4.400 648.360 195.600 648.400 ;
        RECT 0.525 647.000 195.600 648.360 ;
        RECT 0.525 645.680 196.000 647.000 ;
        RECT 4.400 644.280 195.600 645.680 ;
        RECT 0.525 642.960 196.000 644.280 ;
        RECT 0.525 641.600 195.600 642.960 ;
        RECT 4.400 641.560 195.600 641.600 ;
        RECT 4.400 640.240 196.000 641.560 ;
        RECT 4.400 640.200 195.600 640.240 ;
        RECT 0.525 638.840 195.600 640.200 ;
        RECT 0.525 637.520 196.000 638.840 ;
        RECT 4.400 636.120 195.600 637.520 ;
        RECT 0.525 634.800 196.000 636.120 ;
        RECT 0.525 633.440 195.600 634.800 ;
        RECT 4.400 633.400 195.600 633.440 ;
        RECT 4.400 632.080 196.000 633.400 ;
        RECT 4.400 632.040 195.600 632.080 ;
        RECT 0.525 630.680 195.600 632.040 ;
        RECT 0.525 629.360 196.000 630.680 ;
        RECT 4.400 627.960 195.600 629.360 ;
        RECT 0.525 626.640 196.000 627.960 ;
        RECT 0.525 625.280 195.600 626.640 ;
        RECT 4.400 625.240 195.600 625.280 ;
        RECT 4.400 623.920 196.000 625.240 ;
        RECT 4.400 623.880 195.600 623.920 ;
        RECT 0.525 622.520 195.600 623.880 ;
        RECT 0.525 621.200 196.000 622.520 ;
        RECT 4.400 619.800 195.600 621.200 ;
        RECT 0.525 618.480 196.000 619.800 ;
        RECT 0.525 617.120 195.600 618.480 ;
        RECT 4.400 617.080 195.600 617.120 ;
        RECT 4.400 615.760 196.000 617.080 ;
        RECT 4.400 615.720 195.600 615.760 ;
        RECT 0.525 614.360 195.600 615.720 ;
        RECT 0.525 613.040 196.000 614.360 ;
        RECT 4.400 611.640 195.600 613.040 ;
        RECT 0.525 610.320 196.000 611.640 ;
        RECT 0.525 608.960 195.600 610.320 ;
        RECT 4.400 608.920 195.600 608.960 ;
        RECT 4.400 607.600 196.000 608.920 ;
        RECT 4.400 607.560 195.600 607.600 ;
        RECT 0.525 606.200 195.600 607.560 ;
        RECT 0.525 604.880 196.000 606.200 ;
        RECT 4.400 603.480 195.600 604.880 ;
        RECT 0.525 602.160 196.000 603.480 ;
        RECT 0.525 600.800 195.600 602.160 ;
        RECT 4.400 600.760 195.600 600.800 ;
        RECT 4.400 599.440 196.000 600.760 ;
        RECT 4.400 599.400 195.600 599.440 ;
        RECT 0.525 598.040 195.600 599.400 ;
        RECT 0.525 596.720 196.000 598.040 ;
        RECT 4.400 595.320 195.600 596.720 ;
        RECT 0.525 594.000 196.000 595.320 ;
        RECT 0.525 592.640 195.600 594.000 ;
        RECT 4.400 592.600 195.600 592.640 ;
        RECT 4.400 591.280 196.000 592.600 ;
        RECT 4.400 591.240 195.600 591.280 ;
        RECT 0.525 589.880 195.600 591.240 ;
        RECT 0.525 588.560 196.000 589.880 ;
        RECT 4.400 587.160 195.600 588.560 ;
        RECT 0.525 585.840 196.000 587.160 ;
        RECT 0.525 584.480 195.600 585.840 ;
        RECT 4.400 584.440 195.600 584.480 ;
        RECT 4.400 583.120 196.000 584.440 ;
        RECT 4.400 583.080 195.600 583.120 ;
        RECT 0.525 581.720 195.600 583.080 ;
        RECT 0.525 580.400 196.000 581.720 ;
        RECT 4.400 579.000 195.600 580.400 ;
        RECT 0.525 577.680 196.000 579.000 ;
        RECT 0.525 576.320 195.600 577.680 ;
        RECT 4.400 576.280 195.600 576.320 ;
        RECT 4.400 574.960 196.000 576.280 ;
        RECT 4.400 574.920 195.600 574.960 ;
        RECT 0.525 573.560 195.600 574.920 ;
        RECT 0.525 572.240 196.000 573.560 ;
        RECT 4.400 570.840 195.600 572.240 ;
        RECT 0.525 569.520 196.000 570.840 ;
        RECT 0.525 568.160 195.600 569.520 ;
        RECT 4.400 568.120 195.600 568.160 ;
        RECT 4.400 566.800 196.000 568.120 ;
        RECT 4.400 566.760 195.600 566.800 ;
        RECT 0.525 565.400 195.600 566.760 ;
        RECT 0.525 564.080 196.000 565.400 ;
        RECT 4.400 562.680 195.600 564.080 ;
        RECT 0.525 561.360 196.000 562.680 ;
        RECT 0.525 560.000 195.600 561.360 ;
        RECT 4.400 559.960 195.600 560.000 ;
        RECT 4.400 558.640 196.000 559.960 ;
        RECT 4.400 558.600 195.600 558.640 ;
        RECT 0.525 557.240 195.600 558.600 ;
        RECT 0.525 555.920 196.000 557.240 ;
        RECT 4.400 554.520 195.600 555.920 ;
        RECT 0.525 553.200 196.000 554.520 ;
        RECT 0.525 551.840 195.600 553.200 ;
        RECT 4.400 551.800 195.600 551.840 ;
        RECT 4.400 550.480 196.000 551.800 ;
        RECT 4.400 550.440 195.600 550.480 ;
        RECT 0.525 549.080 195.600 550.440 ;
        RECT 0.525 547.760 196.000 549.080 ;
        RECT 4.400 546.360 195.600 547.760 ;
        RECT 0.525 545.040 196.000 546.360 ;
        RECT 0.525 543.680 195.600 545.040 ;
        RECT 4.400 543.640 195.600 543.680 ;
        RECT 4.400 542.320 196.000 543.640 ;
        RECT 4.400 542.280 195.600 542.320 ;
        RECT 0.525 540.920 195.600 542.280 ;
        RECT 0.525 539.600 196.000 540.920 ;
        RECT 4.400 538.200 195.600 539.600 ;
        RECT 0.525 536.880 196.000 538.200 ;
        RECT 0.525 535.520 195.600 536.880 ;
        RECT 4.400 535.480 195.600 535.520 ;
        RECT 4.400 534.160 196.000 535.480 ;
        RECT 4.400 534.120 195.600 534.160 ;
        RECT 0.525 532.760 195.600 534.120 ;
        RECT 0.525 531.440 196.000 532.760 ;
        RECT 4.400 530.040 195.600 531.440 ;
        RECT 0.525 528.720 196.000 530.040 ;
        RECT 0.525 527.360 195.600 528.720 ;
        RECT 4.400 527.320 195.600 527.360 ;
        RECT 4.400 526.000 196.000 527.320 ;
        RECT 4.400 525.960 195.600 526.000 ;
        RECT 0.525 524.600 195.600 525.960 ;
        RECT 0.525 523.280 196.000 524.600 ;
        RECT 4.400 521.880 195.600 523.280 ;
        RECT 0.525 520.560 196.000 521.880 ;
        RECT 0.525 519.200 195.600 520.560 ;
        RECT 4.400 519.160 195.600 519.200 ;
        RECT 4.400 517.840 196.000 519.160 ;
        RECT 4.400 517.800 195.600 517.840 ;
        RECT 0.525 516.440 195.600 517.800 ;
        RECT 0.525 515.120 196.000 516.440 ;
        RECT 4.400 513.720 195.600 515.120 ;
        RECT 0.525 512.400 196.000 513.720 ;
        RECT 0.525 511.040 195.600 512.400 ;
        RECT 4.400 511.000 195.600 511.040 ;
        RECT 4.400 509.680 196.000 511.000 ;
        RECT 4.400 509.640 195.600 509.680 ;
        RECT 0.525 508.280 195.600 509.640 ;
        RECT 0.525 506.960 196.000 508.280 ;
        RECT 4.400 505.560 195.600 506.960 ;
        RECT 0.525 504.240 196.000 505.560 ;
        RECT 0.525 502.880 195.600 504.240 ;
        RECT 4.400 502.840 195.600 502.880 ;
        RECT 4.400 501.520 196.000 502.840 ;
        RECT 4.400 501.480 195.600 501.520 ;
        RECT 0.525 500.120 195.600 501.480 ;
        RECT 0.525 498.800 196.000 500.120 ;
        RECT 4.400 497.400 195.600 498.800 ;
        RECT 0.525 496.080 196.000 497.400 ;
        RECT 0.525 494.720 195.600 496.080 ;
        RECT 4.400 494.680 195.600 494.720 ;
        RECT 4.400 493.360 196.000 494.680 ;
        RECT 4.400 493.320 195.600 493.360 ;
        RECT 0.525 491.960 195.600 493.320 ;
        RECT 0.525 490.640 196.000 491.960 ;
        RECT 4.400 489.240 195.600 490.640 ;
        RECT 0.525 487.920 196.000 489.240 ;
        RECT 0.525 486.560 195.600 487.920 ;
        RECT 4.400 486.520 195.600 486.560 ;
        RECT 4.400 485.200 196.000 486.520 ;
        RECT 4.400 485.160 195.600 485.200 ;
        RECT 0.525 483.800 195.600 485.160 ;
        RECT 0.525 482.480 196.000 483.800 ;
        RECT 4.400 481.080 195.600 482.480 ;
        RECT 0.525 479.760 196.000 481.080 ;
        RECT 0.525 478.400 195.600 479.760 ;
        RECT 4.400 478.360 195.600 478.400 ;
        RECT 4.400 477.040 196.000 478.360 ;
        RECT 4.400 477.000 195.600 477.040 ;
        RECT 0.525 475.640 195.600 477.000 ;
        RECT 0.525 474.320 196.000 475.640 ;
        RECT 4.400 472.920 195.600 474.320 ;
        RECT 0.525 471.600 196.000 472.920 ;
        RECT 0.525 470.240 195.600 471.600 ;
        RECT 4.400 470.200 195.600 470.240 ;
        RECT 4.400 468.880 196.000 470.200 ;
        RECT 4.400 468.840 195.600 468.880 ;
        RECT 0.525 467.480 195.600 468.840 ;
        RECT 0.525 466.160 196.000 467.480 ;
        RECT 4.400 464.760 195.600 466.160 ;
        RECT 0.525 463.440 196.000 464.760 ;
        RECT 0.525 462.080 195.600 463.440 ;
        RECT 4.400 462.040 195.600 462.080 ;
        RECT 4.400 460.720 196.000 462.040 ;
        RECT 4.400 460.680 195.600 460.720 ;
        RECT 0.525 459.320 195.600 460.680 ;
        RECT 0.525 458.000 196.000 459.320 ;
        RECT 4.400 456.600 195.600 458.000 ;
        RECT 0.525 455.280 196.000 456.600 ;
        RECT 0.525 453.920 195.600 455.280 ;
        RECT 4.400 453.880 195.600 453.920 ;
        RECT 4.400 452.560 196.000 453.880 ;
        RECT 4.400 452.520 195.600 452.560 ;
        RECT 0.525 451.160 195.600 452.520 ;
        RECT 0.525 449.840 196.000 451.160 ;
        RECT 4.400 448.440 195.600 449.840 ;
        RECT 0.525 447.120 196.000 448.440 ;
        RECT 0.525 445.760 195.600 447.120 ;
        RECT 4.400 445.720 195.600 445.760 ;
        RECT 4.400 444.400 196.000 445.720 ;
        RECT 4.400 444.360 195.600 444.400 ;
        RECT 0.525 443.000 195.600 444.360 ;
        RECT 0.525 441.680 196.000 443.000 ;
        RECT 4.400 440.280 195.600 441.680 ;
        RECT 0.525 438.960 196.000 440.280 ;
        RECT 0.525 437.600 195.600 438.960 ;
        RECT 4.400 437.560 195.600 437.600 ;
        RECT 4.400 436.240 196.000 437.560 ;
        RECT 4.400 436.200 195.600 436.240 ;
        RECT 0.525 434.840 195.600 436.200 ;
        RECT 0.525 433.520 196.000 434.840 ;
        RECT 4.400 432.120 195.600 433.520 ;
        RECT 0.525 430.800 196.000 432.120 ;
        RECT 0.525 429.440 195.600 430.800 ;
        RECT 4.400 429.400 195.600 429.440 ;
        RECT 4.400 428.080 196.000 429.400 ;
        RECT 4.400 428.040 195.600 428.080 ;
        RECT 0.525 426.680 195.600 428.040 ;
        RECT 0.525 425.360 196.000 426.680 ;
        RECT 4.400 423.960 195.600 425.360 ;
        RECT 0.525 422.640 196.000 423.960 ;
        RECT 0.525 421.280 195.600 422.640 ;
        RECT 4.400 421.240 195.600 421.280 ;
        RECT 4.400 419.920 196.000 421.240 ;
        RECT 4.400 419.880 195.600 419.920 ;
        RECT 0.525 418.520 195.600 419.880 ;
        RECT 0.525 417.200 196.000 418.520 ;
        RECT 4.400 415.800 195.600 417.200 ;
        RECT 0.525 414.480 196.000 415.800 ;
        RECT 0.525 413.120 195.600 414.480 ;
        RECT 4.400 413.080 195.600 413.120 ;
        RECT 4.400 411.760 196.000 413.080 ;
        RECT 4.400 411.720 195.600 411.760 ;
        RECT 0.525 410.360 195.600 411.720 ;
        RECT 0.525 409.040 196.000 410.360 ;
        RECT 4.400 407.640 195.600 409.040 ;
        RECT 0.525 406.320 196.000 407.640 ;
        RECT 0.525 404.960 195.600 406.320 ;
        RECT 4.400 404.920 195.600 404.960 ;
        RECT 4.400 403.600 196.000 404.920 ;
        RECT 4.400 403.560 195.600 403.600 ;
        RECT 0.525 402.200 195.600 403.560 ;
        RECT 0.525 400.880 196.000 402.200 ;
        RECT 4.400 399.480 195.600 400.880 ;
        RECT 0.525 398.160 196.000 399.480 ;
        RECT 0.525 396.800 195.600 398.160 ;
        RECT 4.400 396.760 195.600 396.800 ;
        RECT 4.400 395.440 196.000 396.760 ;
        RECT 4.400 395.400 195.600 395.440 ;
        RECT 0.525 394.040 195.600 395.400 ;
        RECT 0.525 392.720 196.000 394.040 ;
        RECT 4.400 391.320 195.600 392.720 ;
        RECT 0.525 390.000 196.000 391.320 ;
        RECT 0.525 388.640 195.600 390.000 ;
        RECT 4.400 388.600 195.600 388.640 ;
        RECT 4.400 387.280 196.000 388.600 ;
        RECT 4.400 387.240 195.600 387.280 ;
        RECT 0.525 385.880 195.600 387.240 ;
        RECT 0.525 384.560 196.000 385.880 ;
        RECT 4.400 383.160 195.600 384.560 ;
        RECT 0.525 381.840 196.000 383.160 ;
        RECT 0.525 380.480 195.600 381.840 ;
        RECT 4.400 380.440 195.600 380.480 ;
        RECT 4.400 379.120 196.000 380.440 ;
        RECT 4.400 379.080 195.600 379.120 ;
        RECT 0.525 377.720 195.600 379.080 ;
        RECT 0.525 376.400 196.000 377.720 ;
        RECT 4.400 375.000 195.600 376.400 ;
        RECT 0.525 373.680 196.000 375.000 ;
        RECT 0.525 372.320 195.600 373.680 ;
        RECT 4.400 372.280 195.600 372.320 ;
        RECT 4.400 370.960 196.000 372.280 ;
        RECT 4.400 370.920 195.600 370.960 ;
        RECT 0.525 369.560 195.600 370.920 ;
        RECT 0.525 368.240 196.000 369.560 ;
        RECT 4.400 366.840 195.600 368.240 ;
        RECT 0.525 365.520 196.000 366.840 ;
        RECT 0.525 364.160 195.600 365.520 ;
        RECT 4.400 364.120 195.600 364.160 ;
        RECT 4.400 362.800 196.000 364.120 ;
        RECT 4.400 362.760 195.600 362.800 ;
        RECT 0.525 361.400 195.600 362.760 ;
        RECT 0.525 360.080 196.000 361.400 ;
        RECT 4.400 358.680 195.600 360.080 ;
        RECT 0.525 357.360 196.000 358.680 ;
        RECT 0.525 356.000 195.600 357.360 ;
        RECT 4.400 355.960 195.600 356.000 ;
        RECT 4.400 354.640 196.000 355.960 ;
        RECT 4.400 354.600 195.600 354.640 ;
        RECT 0.525 353.240 195.600 354.600 ;
        RECT 0.525 351.920 196.000 353.240 ;
        RECT 4.400 350.520 195.600 351.920 ;
        RECT 0.525 349.200 196.000 350.520 ;
        RECT 0.525 347.840 195.600 349.200 ;
        RECT 4.400 347.800 195.600 347.840 ;
        RECT 4.400 346.480 196.000 347.800 ;
        RECT 4.400 346.440 195.600 346.480 ;
        RECT 0.525 345.080 195.600 346.440 ;
        RECT 0.525 343.760 196.000 345.080 ;
        RECT 4.400 342.360 195.600 343.760 ;
        RECT 0.525 341.040 196.000 342.360 ;
        RECT 0.525 339.680 195.600 341.040 ;
        RECT 4.400 339.640 195.600 339.680 ;
        RECT 4.400 338.320 196.000 339.640 ;
        RECT 4.400 338.280 195.600 338.320 ;
        RECT 0.525 336.920 195.600 338.280 ;
        RECT 0.525 335.600 196.000 336.920 ;
        RECT 4.400 334.200 195.600 335.600 ;
        RECT 0.525 332.880 196.000 334.200 ;
        RECT 0.525 331.520 195.600 332.880 ;
        RECT 4.400 331.480 195.600 331.520 ;
        RECT 4.400 330.160 196.000 331.480 ;
        RECT 4.400 330.120 195.600 330.160 ;
        RECT 0.525 328.760 195.600 330.120 ;
        RECT 0.525 327.440 196.000 328.760 ;
        RECT 4.400 326.040 195.600 327.440 ;
        RECT 0.525 324.720 196.000 326.040 ;
        RECT 0.525 323.360 195.600 324.720 ;
        RECT 4.400 323.320 195.600 323.360 ;
        RECT 4.400 322.000 196.000 323.320 ;
        RECT 4.400 321.960 195.600 322.000 ;
        RECT 0.525 320.600 195.600 321.960 ;
        RECT 0.525 319.280 196.000 320.600 ;
        RECT 4.400 317.880 195.600 319.280 ;
        RECT 0.525 316.560 196.000 317.880 ;
        RECT 0.525 315.200 195.600 316.560 ;
        RECT 4.400 315.160 195.600 315.200 ;
        RECT 4.400 313.840 196.000 315.160 ;
        RECT 4.400 313.800 195.600 313.840 ;
        RECT 0.525 312.440 195.600 313.800 ;
        RECT 0.525 311.120 196.000 312.440 ;
        RECT 4.400 309.720 195.600 311.120 ;
        RECT 0.525 308.400 196.000 309.720 ;
        RECT 0.525 307.040 195.600 308.400 ;
        RECT 4.400 307.000 195.600 307.040 ;
        RECT 4.400 305.680 196.000 307.000 ;
        RECT 4.400 305.640 195.600 305.680 ;
        RECT 0.525 304.280 195.600 305.640 ;
        RECT 0.525 302.960 196.000 304.280 ;
        RECT 4.400 301.560 195.600 302.960 ;
        RECT 0.525 300.240 196.000 301.560 ;
        RECT 0.525 298.880 195.600 300.240 ;
        RECT 4.400 298.840 195.600 298.880 ;
        RECT 4.400 297.520 196.000 298.840 ;
        RECT 4.400 297.480 195.600 297.520 ;
        RECT 0.525 296.120 195.600 297.480 ;
        RECT 0.525 294.800 196.000 296.120 ;
        RECT 4.400 293.400 195.600 294.800 ;
        RECT 0.525 292.080 196.000 293.400 ;
        RECT 0.525 290.720 195.600 292.080 ;
        RECT 4.400 290.680 195.600 290.720 ;
        RECT 4.400 289.360 196.000 290.680 ;
        RECT 4.400 289.320 195.600 289.360 ;
        RECT 0.525 287.960 195.600 289.320 ;
        RECT 0.525 286.640 196.000 287.960 ;
        RECT 4.400 285.240 195.600 286.640 ;
        RECT 0.525 283.920 196.000 285.240 ;
        RECT 0.525 282.560 195.600 283.920 ;
        RECT 4.400 282.520 195.600 282.560 ;
        RECT 4.400 281.200 196.000 282.520 ;
        RECT 4.400 281.160 195.600 281.200 ;
        RECT 0.525 279.800 195.600 281.160 ;
        RECT 0.525 278.480 196.000 279.800 ;
        RECT 4.400 277.080 195.600 278.480 ;
        RECT 0.525 275.760 196.000 277.080 ;
        RECT 0.525 274.400 195.600 275.760 ;
        RECT 4.400 274.360 195.600 274.400 ;
        RECT 4.400 273.040 196.000 274.360 ;
        RECT 4.400 273.000 195.600 273.040 ;
        RECT 0.525 271.640 195.600 273.000 ;
        RECT 0.525 270.320 196.000 271.640 ;
        RECT 4.400 268.920 195.600 270.320 ;
        RECT 0.525 267.600 196.000 268.920 ;
        RECT 0.525 266.240 195.600 267.600 ;
        RECT 4.400 266.200 195.600 266.240 ;
        RECT 4.400 264.880 196.000 266.200 ;
        RECT 4.400 264.840 195.600 264.880 ;
        RECT 0.525 263.480 195.600 264.840 ;
        RECT 0.525 262.160 196.000 263.480 ;
        RECT 4.400 260.760 195.600 262.160 ;
        RECT 0.525 259.440 196.000 260.760 ;
        RECT 0.525 258.080 195.600 259.440 ;
        RECT 4.400 258.040 195.600 258.080 ;
        RECT 4.400 256.720 196.000 258.040 ;
        RECT 4.400 256.680 195.600 256.720 ;
        RECT 0.525 255.320 195.600 256.680 ;
        RECT 0.525 254.000 196.000 255.320 ;
        RECT 4.400 252.600 195.600 254.000 ;
        RECT 0.525 251.280 196.000 252.600 ;
        RECT 0.525 249.920 195.600 251.280 ;
        RECT 4.400 249.880 195.600 249.920 ;
        RECT 4.400 248.560 196.000 249.880 ;
        RECT 4.400 248.520 195.600 248.560 ;
        RECT 0.525 247.160 195.600 248.520 ;
        RECT 0.525 245.840 196.000 247.160 ;
        RECT 4.400 244.440 195.600 245.840 ;
        RECT 0.525 243.120 196.000 244.440 ;
        RECT 0.525 241.760 195.600 243.120 ;
        RECT 4.400 241.720 195.600 241.760 ;
        RECT 4.400 240.400 196.000 241.720 ;
        RECT 4.400 240.360 195.600 240.400 ;
        RECT 0.525 239.000 195.600 240.360 ;
        RECT 0.525 237.680 196.000 239.000 ;
        RECT 4.400 236.280 195.600 237.680 ;
        RECT 0.525 234.960 196.000 236.280 ;
        RECT 0.525 233.600 195.600 234.960 ;
        RECT 4.400 233.560 195.600 233.600 ;
        RECT 4.400 232.240 196.000 233.560 ;
        RECT 4.400 232.200 195.600 232.240 ;
        RECT 0.525 230.840 195.600 232.200 ;
        RECT 0.525 229.520 196.000 230.840 ;
        RECT 4.400 228.120 195.600 229.520 ;
        RECT 0.525 226.800 196.000 228.120 ;
        RECT 0.525 225.440 195.600 226.800 ;
        RECT 4.400 225.400 195.600 225.440 ;
        RECT 4.400 224.080 196.000 225.400 ;
        RECT 4.400 224.040 195.600 224.080 ;
        RECT 0.525 222.680 195.600 224.040 ;
        RECT 0.525 221.360 196.000 222.680 ;
        RECT 4.400 219.960 195.600 221.360 ;
        RECT 0.525 218.640 196.000 219.960 ;
        RECT 0.525 217.280 195.600 218.640 ;
        RECT 4.400 217.240 195.600 217.280 ;
        RECT 4.400 215.920 196.000 217.240 ;
        RECT 4.400 215.880 195.600 215.920 ;
        RECT 0.525 214.520 195.600 215.880 ;
        RECT 0.525 213.200 196.000 214.520 ;
        RECT 4.400 211.800 195.600 213.200 ;
        RECT 0.525 210.480 196.000 211.800 ;
        RECT 0.525 209.120 195.600 210.480 ;
        RECT 4.400 209.080 195.600 209.120 ;
        RECT 4.400 207.760 196.000 209.080 ;
        RECT 4.400 207.720 195.600 207.760 ;
        RECT 0.525 206.360 195.600 207.720 ;
        RECT 0.525 205.040 196.000 206.360 ;
        RECT 4.400 203.640 195.600 205.040 ;
        RECT 0.525 202.320 196.000 203.640 ;
        RECT 0.525 200.960 195.600 202.320 ;
        RECT 4.400 200.920 195.600 200.960 ;
        RECT 4.400 199.600 196.000 200.920 ;
        RECT 4.400 199.560 195.600 199.600 ;
        RECT 0.525 198.200 195.600 199.560 ;
        RECT 0.525 196.880 196.000 198.200 ;
        RECT 4.400 195.480 195.600 196.880 ;
        RECT 0.525 194.160 196.000 195.480 ;
        RECT 0.525 192.800 195.600 194.160 ;
        RECT 4.400 192.760 195.600 192.800 ;
        RECT 4.400 191.440 196.000 192.760 ;
        RECT 4.400 191.400 195.600 191.440 ;
        RECT 0.525 190.040 195.600 191.400 ;
        RECT 0.525 188.720 196.000 190.040 ;
        RECT 4.400 187.320 195.600 188.720 ;
        RECT 0.525 186.000 196.000 187.320 ;
        RECT 0.525 184.640 195.600 186.000 ;
        RECT 4.400 184.600 195.600 184.640 ;
        RECT 4.400 183.280 196.000 184.600 ;
        RECT 4.400 183.240 195.600 183.280 ;
        RECT 0.525 181.880 195.600 183.240 ;
        RECT 0.525 180.560 196.000 181.880 ;
        RECT 4.400 179.160 195.600 180.560 ;
        RECT 0.525 177.840 196.000 179.160 ;
        RECT 0.525 176.480 195.600 177.840 ;
        RECT 4.400 176.440 195.600 176.480 ;
        RECT 4.400 175.120 196.000 176.440 ;
        RECT 4.400 175.080 195.600 175.120 ;
        RECT 0.525 173.720 195.600 175.080 ;
        RECT 0.525 172.400 196.000 173.720 ;
        RECT 4.400 171.000 195.600 172.400 ;
        RECT 0.525 169.680 196.000 171.000 ;
        RECT 0.525 168.320 195.600 169.680 ;
        RECT 4.400 168.280 195.600 168.320 ;
        RECT 4.400 166.960 196.000 168.280 ;
        RECT 4.400 166.920 195.600 166.960 ;
        RECT 0.525 165.560 195.600 166.920 ;
        RECT 0.525 164.240 196.000 165.560 ;
        RECT 4.400 162.840 195.600 164.240 ;
        RECT 0.525 161.520 196.000 162.840 ;
        RECT 0.525 160.160 195.600 161.520 ;
        RECT 4.400 160.120 195.600 160.160 ;
        RECT 4.400 158.800 196.000 160.120 ;
        RECT 4.400 158.760 195.600 158.800 ;
        RECT 0.525 157.400 195.600 158.760 ;
        RECT 0.525 156.080 196.000 157.400 ;
        RECT 4.400 154.680 195.600 156.080 ;
        RECT 0.525 153.360 196.000 154.680 ;
        RECT 0.525 152.000 195.600 153.360 ;
        RECT 4.400 151.960 195.600 152.000 ;
        RECT 4.400 150.600 196.000 151.960 ;
        RECT 0.525 147.920 196.000 150.600 ;
        RECT 4.400 146.520 196.000 147.920 ;
        RECT 0.525 143.840 196.000 146.520 ;
        RECT 4.400 142.440 196.000 143.840 ;
        RECT 0.525 139.760 196.000 142.440 ;
        RECT 4.400 138.360 196.000 139.760 ;
        RECT 0.525 135.680 196.000 138.360 ;
        RECT 4.400 134.280 196.000 135.680 ;
        RECT 0.525 131.600 196.000 134.280 ;
        RECT 4.400 130.200 196.000 131.600 ;
        RECT 0.525 127.520 196.000 130.200 ;
        RECT 4.400 126.120 196.000 127.520 ;
        RECT 0.525 123.440 196.000 126.120 ;
        RECT 4.400 122.040 196.000 123.440 ;
        RECT 0.525 119.360 196.000 122.040 ;
        RECT 4.400 117.960 196.000 119.360 ;
        RECT 0.525 115.280 196.000 117.960 ;
        RECT 4.400 113.880 196.000 115.280 ;
        RECT 0.525 111.200 196.000 113.880 ;
        RECT 4.400 109.800 196.000 111.200 ;
        RECT 0.525 107.120 196.000 109.800 ;
        RECT 4.400 105.720 196.000 107.120 ;
        RECT 0.525 103.040 196.000 105.720 ;
        RECT 4.400 101.640 196.000 103.040 ;
        RECT 0.525 98.960 196.000 101.640 ;
        RECT 4.400 97.560 196.000 98.960 ;
        RECT 0.525 10.715 196.000 97.560 ;
      LAYER met4 ;
        RECT 3.055 13.775 20.640 1080.345 ;
        RECT 23.040 13.775 97.440 1080.345 ;
        RECT 99.840 13.775 174.240 1080.345 ;
        RECT 176.640 13.775 191.065 1080.345 ;
  END
END multiplexer
END LIBRARY

