* NGSPICE file created from multiplexer.ext - technology: sky130B

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt multiplexer cap_addr[0] cap_addr[1] cap_addr[2] cap_addr[3] cap_addr[4] cap_addr[5]
+ cap_addr[6] cap_addr[7] cap_addr[8] cap_io_in[0] cap_io_in[1] cap_io_in[2] cap_io_in[3]
+ cap_io_in[4] cap_io_in[5] cap_io_in[6] cap_io_in[7] cap_io_in[8] custom_settings[0]
+ custom_settings[10] custom_settings[11] custom_settings[12] custom_settings[13]
+ custom_settings[14] custom_settings[15] custom_settings[16] custom_settings[17]
+ custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20] custom_settings[21]
+ custom_settings[22] custom_settings[23] custom_settings[24] custom_settings[25]
+ custom_settings[26] custom_settings[27] custom_settings[28] custom_settings[29]
+ custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3] custom_settings[4]
+ custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8] custom_settings[9]
+ io_in_0 io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2]
+ io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_oeb_6502
+ io_oeb_8x305[0] io_oeb_8x305[1] io_oeb_8x305[2] io_oeb_8x305[3] io_oeb_8x305[4]
+ io_oeb_as1802 io_oeb_scrapcpu[0] io_oeb_scrapcpu[10] io_oeb_scrapcpu[11] io_oeb_scrapcpu[12]
+ io_oeb_scrapcpu[13] io_oeb_scrapcpu[14] io_oeb_scrapcpu[15] io_oeb_scrapcpu[16]
+ io_oeb_scrapcpu[17] io_oeb_scrapcpu[18] io_oeb_scrapcpu[19] io_oeb_scrapcpu[1] io_oeb_scrapcpu[20]
+ io_oeb_scrapcpu[21] io_oeb_scrapcpu[22] io_oeb_scrapcpu[23] io_oeb_scrapcpu[24]
+ io_oeb_scrapcpu[25] io_oeb_scrapcpu[26] io_oeb_scrapcpu[27] io_oeb_scrapcpu[28]
+ io_oeb_scrapcpu[29] io_oeb_scrapcpu[2] io_oeb_scrapcpu[30] io_oeb_scrapcpu[31] io_oeb_scrapcpu[32]
+ io_oeb_scrapcpu[33] io_oeb_scrapcpu[34] io_oeb_scrapcpu[35] io_oeb_scrapcpu[3] io_oeb_scrapcpu[4]
+ io_oeb_scrapcpu[5] io_oeb_scrapcpu[6] io_oeb_scrapcpu[7] io_oeb_scrapcpu[8] io_oeb_scrapcpu[9]
+ io_oeb_vliw[0] io_oeb_vliw[10] io_oeb_vliw[11] io_oeb_vliw[12] io_oeb_vliw[13] io_oeb_vliw[14]
+ io_oeb_vliw[15] io_oeb_vliw[16] io_oeb_vliw[17] io_oeb_vliw[18] io_oeb_vliw[19]
+ io_oeb_vliw[1] io_oeb_vliw[20] io_oeb_vliw[21] io_oeb_vliw[22] io_oeb_vliw[23] io_oeb_vliw[24]
+ io_oeb_vliw[25] io_oeb_vliw[26] io_oeb_vliw[27] io_oeb_vliw[28] io_oeb_vliw[29]
+ io_oeb_vliw[2] io_oeb_vliw[30] io_oeb_vliw[31] io_oeb_vliw[32] io_oeb_vliw[33] io_oeb_vliw[34]
+ io_oeb_vliw[35] io_oeb_vliw[3] io_oeb_vliw[4] io_oeb_vliw[5] io_oeb_vliw[6] io_oeb_vliw[7]
+ io_oeb_vliw[8] io_oeb_vliw[9] io_oeb_z80[0] io_oeb_z80[10] io_oeb_z80[11] io_oeb_z80[12]
+ io_oeb_z80[13] io_oeb_z80[14] io_oeb_z80[15] io_oeb_z80[16] io_oeb_z80[17] io_oeb_z80[18]
+ io_oeb_z80[19] io_oeb_z80[1] io_oeb_z80[20] io_oeb_z80[21] io_oeb_z80[22] io_oeb_z80[23]
+ io_oeb_z80[24] io_oeb_z80[25] io_oeb_z80[26] io_oeb_z80[27] io_oeb_z80[28] io_oeb_z80[29]
+ io_oeb_z80[2] io_oeb_z80[30] io_oeb_z80[31] io_oeb_z80[32] io_oeb_z80[33] io_oeb_z80[34]
+ io_oeb_z80[35] io_oeb_z80[3] io_oeb_z80[4] io_oeb_z80[5] io_oeb_z80[6] io_oeb_z80[7]
+ io_oeb_z80[8] io_oeb_z80[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ io_out[9] io_out_6502[0] io_out_6502[10] io_out_6502[11] io_out_6502[12] io_out_6502[13]
+ io_out_6502[14] io_out_6502[15] io_out_6502[16] io_out_6502[17] io_out_6502[18]
+ io_out_6502[19] io_out_6502[1] io_out_6502[20] io_out_6502[21] io_out_6502[22] io_out_6502[23]
+ io_out_6502[24] io_out_6502[25] io_out_6502[26] io_out_6502[27] io_out_6502[28]
+ io_out_6502[29] io_out_6502[2] io_out_6502[30] io_out_6502[31] io_out_6502[32] io_out_6502[33]
+ io_out_6502[34] io_out_6502[35] io_out_6502[3] io_out_6502[4] io_out_6502[5] io_out_6502[6]
+ io_out_6502[7] io_out_6502[8] io_out_6502[9] io_out_8x305[0] io_out_8x305[10] io_out_8x305[11]
+ io_out_8x305[12] io_out_8x305[13] io_out_8x305[14] io_out_8x305[15] io_out_8x305[16]
+ io_out_8x305[17] io_out_8x305[18] io_out_8x305[19] io_out_8x305[1] io_out_8x305[20]
+ io_out_8x305[21] io_out_8x305[22] io_out_8x305[23] io_out_8x305[24] io_out_8x305[25]
+ io_out_8x305[26] io_out_8x305[27] io_out_8x305[28] io_out_8x305[29] io_out_8x305[2]
+ io_out_8x305[30] io_out_8x305[31] io_out_8x305[32] io_out_8x305[33] io_out_8x305[34]
+ io_out_8x305[35] io_out_8x305[3] io_out_8x305[4] io_out_8x305[5] io_out_8x305[6]
+ io_out_8x305[7] io_out_8x305[8] io_out_8x305[9] io_out_as1802[0] io_out_as1802[10]
+ io_out_as1802[11] io_out_as1802[12] io_out_as1802[13] io_out_as1802[14] io_out_as1802[15]
+ io_out_as1802[16] io_out_as1802[17] io_out_as1802[18] io_out_as1802[19] io_out_as1802[1]
+ io_out_as1802[20] io_out_as1802[21] io_out_as1802[22] io_out_as1802[23] io_out_as1802[24]
+ io_out_as1802[25] io_out_as1802[26] io_out_as1802[27] io_out_as1802[28] io_out_as1802[29]
+ io_out_as1802[2] io_out_as1802[30] io_out_as1802[31] io_out_as1802[32] io_out_as1802[33]
+ io_out_as1802[34] io_out_as1802[35] io_out_as1802[3] io_out_as1802[4] io_out_as1802[5]
+ io_out_as1802[6] io_out_as1802[7] io_out_as1802[8] io_out_as1802[9] io_out_scrapcpu[0]
+ io_out_scrapcpu[10] io_out_scrapcpu[11] io_out_scrapcpu[12] io_out_scrapcpu[13]
+ io_out_scrapcpu[14] io_out_scrapcpu[15] io_out_scrapcpu[16] io_out_scrapcpu[17]
+ io_out_scrapcpu[18] io_out_scrapcpu[19] io_out_scrapcpu[1] io_out_scrapcpu[20] io_out_scrapcpu[21]
+ io_out_scrapcpu[22] io_out_scrapcpu[23] io_out_scrapcpu[24] io_out_scrapcpu[25]
+ io_out_scrapcpu[26] io_out_scrapcpu[27] io_out_scrapcpu[28] io_out_scrapcpu[29]
+ io_out_scrapcpu[2] io_out_scrapcpu[30] io_out_scrapcpu[31] io_out_scrapcpu[32] io_out_scrapcpu[33]
+ io_out_scrapcpu[34] io_out_scrapcpu[35] io_out_scrapcpu[3] io_out_scrapcpu[4] io_out_scrapcpu[5]
+ io_out_scrapcpu[6] io_out_scrapcpu[7] io_out_scrapcpu[8] io_out_scrapcpu[9] io_out_vliw[0]
+ io_out_vliw[10] io_out_vliw[11] io_out_vliw[12] io_out_vliw[13] io_out_vliw[14]
+ io_out_vliw[15] io_out_vliw[16] io_out_vliw[17] io_out_vliw[18] io_out_vliw[19]
+ io_out_vliw[1] io_out_vliw[20] io_out_vliw[21] io_out_vliw[22] io_out_vliw[23] io_out_vliw[24]
+ io_out_vliw[25] io_out_vliw[26] io_out_vliw[27] io_out_vliw[28] io_out_vliw[29]
+ io_out_vliw[2] io_out_vliw[30] io_out_vliw[31] io_out_vliw[32] io_out_vliw[33] io_out_vliw[34]
+ io_out_vliw[35] io_out_vliw[3] io_out_vliw[4] io_out_vliw[5] io_out_vliw[6] io_out_vliw[7]
+ io_out_vliw[8] io_out_vliw[9] io_out_z80[0] io_out_z80[10] io_out_z80[11] io_out_z80[12]
+ io_out_z80[13] io_out_z80[14] io_out_z80[15] io_out_z80[16] io_out_z80[17] io_out_z80[18]
+ io_out_z80[19] io_out_z80[1] io_out_z80[20] io_out_z80[21] io_out_z80[22] io_out_z80[23]
+ io_out_z80[24] io_out_z80[25] io_out_z80[26] io_out_z80[27] io_out_z80[28] io_out_z80[29]
+ io_out_z80[2] io_out_z80[30] io_out_z80[31] io_out_z80[32] io_out_z80[33] io_out_z80[34]
+ io_out_z80[35] io_out_z80[3] io_out_z80[4] io_out_z80[5] io_out_z80[6] io_out_z80[7]
+ io_out_z80[8] io_out_z80[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] rst_6502 rst_8x305 rst_as1802 rst_scrapcpu
+ rst_vliw rst_z80 vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i
XFILLER_0_280_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_300_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_300_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 hold675/X vssd1 vssd1 vccd1 vccd1 _1090_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 hold691/X vssd1 vssd1 vccd1 vccd1 _0983_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold351 _1224_/Q vssd1 vssd1 vccd1 vccd1 _0851_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold384 hold789/X vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 hold785/X vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 hold744/X vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_244_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_244_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_341_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output513_A _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0892__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0985_ hold562/X _0987_/B _0996_/A vssd1 vssd1 vccd1 vccd1 _0985_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_313_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput401 _1106_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[19] sky130_fd_sc_hd__buf_12
XFILLER_0_285_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput412 _1116_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[29] sky130_fd_sc_hd__buf_12
Xoutput423 _1239_/A vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput434 _1249_/A vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput456 _1236_/A vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__buf_12
Xoutput467 _0673_/X vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
Xoutput445 hold78/A vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__buf_12
Xoutput478 _0713_/X vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_12
XFILLER_0_226_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput489 _1181_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_226_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1073__B _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0883__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold170 hold528/X vssd1 vssd1 vccd1 vccd1 _1112_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1264__A _1264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 _0936_/Y vssd1 vssd1 vccd1 vccd1 _1148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _0905_/Y vssd1 vssd1 vccd1 vccd1 _0906_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_386_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0770_ _0851_/A _0841_/B _0851_/B vssd1 vssd1 vccd1 vccd1 _0770_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA_output463_A _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_310_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1253_ _1253_/A vssd1 vssd1 vccd1 vccd1 _1253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1184_ _1184_/CLK _1184_/D vssd1 vssd1 vccd1 vccd1 _1184_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0518__A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_377_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_345_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0968_ _0967_/A _1157_/Q _0967_/C hold600/A vssd1 vssd1 vccd1 vccd1 _0968_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0899_ hold240/X _0880_/A _0898_/X vssd1 vssd1 vccd1 vccd1 _0899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_258_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_357_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_258_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_373_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_387_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_306_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_322_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0623__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_311_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_359_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_374_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0822_ hold235/X _0775_/Y _0821_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0822_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_126_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0753_ _0767_/A _0767_/B _0753_/C vssd1 vssd1 vccd1 vccd1 _0753_/X sky130_fd_sc_hd__and3_4
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0684_ _0684_/A1 _0732_/A2 _0696_/B1 _0684_/B2 vssd1 vssd1 vccd1 vccd1 _0685_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_381_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_263_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0550__A1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1236_ _1236_/A vssd1 vssd1 vccd1 vccd1 _1236_/X sky130_fd_sc_hd__buf_1
XFILLER_0_223_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1167_ _1167_/CLK _1167_/D vssd1 vssd1 vccd1 vccd1 _1167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1098_ _1224_/CLK _1098_/D vssd1 vssd1 vccd1 vccd1 _1098_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0541__A1 _0541_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_292_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output426_A _1242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1021_ _1021_/A _1021_/B vssd1 vssd1 vccd1 vccd1 _1021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0599__A1 _0599_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold703 _1215_/Q vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
X_0805_ _0805_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0805_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0736_ _0736_/A1 _0508_/B _0748_/B1 _0736_/B2 vssd1 vssd1 vccd1 vccd1 _0737_/C sky130_fd_sc_hd__a22o_1
Xhold725 _1181_/Q vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _0818_/X vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 _1129_/Q vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold769 _1183_/Q vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _1170_/Q vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold747 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_295_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0667_ _0667_/A1 _0514_/B _0683_/B1 _0667_/B2 vssd1 vssd1 vccd1 vccd1 _0669_/B sky130_fd_sc_hd__a22o_1
X_0598_ input43/X _0598_/A2 _0598_/B1 input79/X vssd1 vssd1 vccd1 vccd1 _0598_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_354_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1219_ _1221_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 _1219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0826__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_380_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_274_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0762__A1 _1093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput301 io_out_vliw[5] vssd1 vssd1 vccd1 vccd1 _0628_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_274_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput312 io_out_z80[15] vssd1 vssd1 vccd1 vccd1 _0666_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_264_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput334 io_out_z80[35] vssd1 vssd1 vccd1 vccd1 _0746_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_227_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput323 io_out_z80[25] vssd1 vssd1 vccd1 vccd1 _0706_/A1 sky130_fd_sc_hd__buf_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput345 hold414/X vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__clkbuf_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput367 hold519/X vssd1 vssd1 vccd1 vccd1 hold520/A sky130_fd_sc_hd__clkbuf_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput378 hold465/X vssd1 vssd1 vccd1 vccd1 hold466/A sky130_fd_sc_hd__clkbuf_1
Xinput356 hold468/X vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_388_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__buf_1
XFILLER_0_199_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_388_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_280_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_356_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_312_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0521_ hold93/X hold87/X _0767_/B hold77/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_277_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output543_A hold303/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_280_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0808__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1004_ _1004_/A _1008_/C vssd1 vssd1 vccd1 vccd1 _1007_/B sky130_fd_sc_hd__and2_1
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0526__A _0526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_362_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_343_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold511 hold511/A vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1076__B _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 _0832_/X vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _1062_/Y vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _1023_/Y vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0744__B2 _0744_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0719_ _0719_/A1 _0593_/A _0516_/B _0719_/B2 vssd1 vssd1 vccd1 vccd1 _0721_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_256_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold555 _1069_/Y vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _1031_/X vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 _1009_/Y vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold566 hold738/X vssd1 vssd1 vccd1 vccd1 _0851_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold599 _1159_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_271_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout574_A _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1267__A _1267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0735__B2 _0735_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0735__A1 _0735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput120 io_oeb_z80[4] vssd1 vssd1 vccd1 vccd1 _0533_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_275_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput153 io_out_6502[34] vssd1 vssd1 vccd1 vccd1 _0743_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput142 io_out_6502[24] vssd1 vssd1 vccd1 vccd1 _0703_/A1 sky130_fd_sc_hd__buf_2
Xinput131 io_out_6502[14] vssd1 vssd1 vccd1 vccd1 _0663_/A1 sky130_fd_sc_hd__buf_2
Xinput186 io_out_8x305[31] vssd1 vssd1 vccd1 vccd1 _0730_/B2 sky130_fd_sc_hd__buf_2
Xinput175 io_out_8x305[21] vssd1 vssd1 vccd1 vccd1 _0690_/B2 sky130_fd_sc_hd__buf_2
Xinput164 io_out_8x305[11] vssd1 vssd1 vccd1 vccd1 _0650_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_215_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput197 io_out_8x305[9] vssd1 vssd1 vccd1 vccd1 _0642_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_270_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0671__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output493_A _0629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_344_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_325_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0726__B2 _0726_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0504_ hold76/X hold92/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__or2_1
XFILLER_0_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_280_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_288_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold341 _1122_/Q vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 hold673/X vssd1 vssd1 vccd1 vccd1 _1102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _0882_/C vssd1 vssd1 vccd1 vccd1 _1082_/C sky130_fd_sc_hd__buf_2
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold385 hold783/X vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 hold734/X vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _0779_/A vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _0974_/Y vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_256_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_244_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_392_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_261_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_381_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0708__B2 _0708_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0507__C _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_360_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0984_ _1017_/A _1017_/B vssd1 vssd1 vccd1 vccd1 _0987_/B sky130_fd_sc_hd__and2_1
XFILLER_0_320_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0947__A1 hold217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput402 _1088_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[1] sky130_fd_sc_hd__buf_12
Xoutput413 _1089_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[2] sky130_fd_sc_hd__buf_12
Xoutput424 _1240_/A vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput435 _1250_/A vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__buf_12
Xoutput457 _1237_/A vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput468 _0677_/X vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
Xoutput446 _0592_/X vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__buf_12
XFILLER_0_285_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput479 _0717_/X vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_346_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_355_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0635__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0938__A1 hold185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold160 _1121_/Q vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold775/X vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold182 hold383/X vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__clkbuf_2
Xhold193 _0906_/Y vssd1 vssd1 vccd1 vccd1 _1138_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_244_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0929__A1 hold173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1051__B1 _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output456_A _1236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1252_ _1252_/A vssd1 vssd1 vccd1 vccd1 _1252_/X sky130_fd_sc_hd__buf_1
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1175_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1183_ _1184_/CLK _1183_/D vssd1 vssd1 vccd1 vccd1 _1183_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0518__B _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_392_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0967_ _0967_/A _0967_/B _0967_/C _0967_/D vssd1 vssd1 vccd1 vccd1 _1017_/A sky130_fd_sc_hd__and4_2
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0898_ hold260/X _0776_/A hold605/A _1016_/B _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0898_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_357_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_306_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_395_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0792__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_283_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_374_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0821_ _0821_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0821_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0752_ input2/X _1088_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0753_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0683_ _0683_/A1 _0747_/A2 _0683_/B1 _0683_/B2 vssd1 vssd1 vccd1 vccd1 _0685_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_177_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0801__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1235_ _1235_/A vssd1 vssd1 vccd1 vccd1 _1235_/X sky130_fd_sc_hd__buf_1
XFILLER_0_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1166_ _1224_/CLK _1166_/D vssd1 vssd1 vccd1 vccd1 _1166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_384_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1097_ _1204_/CLK _1097_/D vssd1 vssd1 vccd1 vccd1 _1097_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_392_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_286_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold447_A hold19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_371_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0780__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_292_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output419_A _1093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1020_ _1024_/A _1037_/B vssd1 vssd1 vccd1 vccd1 _1020_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_374_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0804_ hold260/X _0810_/A2 _0803_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0804_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_330_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_287_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0735_ _0735_/A1 _0747_/A2 _0516_/B _0735_/B2 vssd1 vssd1 vccd1 vccd1 _0737_/B sky130_fd_sc_hd__a22o_1
Xhold704 _1059_/X vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 _1124_/Q vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 _1209_/Q vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 _1225_/Q vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_330_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0666_ _0666_/A1 _0674_/A2 _0674_/B1 _0666_/B2 vssd1 vssd1 vccd1 vccd1 _0669_/A sky130_fd_sc_hd__a22o_1
Xhold759 _1167_/Q vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold748 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_295_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0597_ _0597_/A1 _0605_/A2 hold95/X _0596_/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__a211o_4
XANTENNA__0523__A2 hold82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1218_ _1221_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _1218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1149_ _1154_/CLK _1149_/D vssd1 vssd1 vccd1 vccd1 _1149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout617_A _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_380_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_306_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput302 io_out_vliw[6] vssd1 vssd1 vccd1 vccd1 _0632_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_328_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput324 io_out_z80[26] vssd1 vssd1 vccd1 vccd1 _0710_/A1 sky130_fd_sc_hd__buf_1
Xinput313 io_out_z80[16] vssd1 vssd1 vccd1 vccd1 _0670_/A1 sky130_fd_sc_hd__buf_1
Xinput335 io_out_z80[3] vssd1 vssd1 vccd1 vccd1 _0618_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput368 hold513/X vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__buf_1
Xinput357 hold471/X vssd1 vssd1 vccd1 vccd1 hold472/A sky130_fd_sc_hd__clkbuf_1
Xinput346 hold417/X vssd1 vssd1 vccd1 vccd1 hold418/A sky130_fd_sc_hd__clkbuf_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput379 hold453/X vssd1 vssd1 vccd1 vccd1 hold454/A sky130_fd_sc_hd__clkbuf_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_388_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_12
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__buf_2
XFILLER_0_388_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_371_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_289_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0520_ hold99/A hold86/X vssd1 vssd1 vccd1 vccd1 _0767_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output536_A _0516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0910__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1003_ _1004_/A _1008_/C vssd1 vssd1 vccd1 vccd1 _1003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_362_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold501 hold59/X vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_0718_ _0718_/A1 _0505_/Y _0518_/B _0718_/B2 vssd1 vssd1 vccd1 vccd1 _0721_/A sky130_fd_sc_hd__a22o_1
Xhold523 _1116_/Q vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _1063_/X vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _1026_/Y vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold556 _1070_/X vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _1179_/Q vssd1 vssd1 vccd1 vccd1 _1050_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold567 _0770_/Y vssd1 vssd1 vccd1 vccd1 _0775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_365_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0649_ _0649_/A _0649_/B _0649_/C vssd1 vssd1 vccd1 vccd1 _0649_/X sky130_fd_sc_hd__or3_4
Xhold589 _1010_/X vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0901__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0680__B2 _0680_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_353_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput110 io_oeb_z80[28] vssd1 vssd1 vccd1 vccd1 _0588_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_247_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput121 io_oeb_z80[5] vssd1 vssd1 vccd1 vccd1 _0535_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput154 io_out_6502[35] vssd1 vssd1 vccd1 vccd1 _0747_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput143 io_out_6502[25] vssd1 vssd1 vccd1 vccd1 _0707_/A1 sky130_fd_sc_hd__buf_2
Xinput132 io_out_6502[15] vssd1 vssd1 vccd1 vccd1 _0667_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_355_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput187 io_out_8x305[32] vssd1 vssd1 vccd1 vccd1 _0734_/B2 sky130_fd_sc_hd__buf_2
Xinput176 io_out_8x305[22] vssd1 vssd1 vccd1 vccd1 _0694_/B2 sky130_fd_sc_hd__buf_2
Xinput165 io_out_8x305[12] vssd1 vssd1 vccd1 vccd1 _0654_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput198 io_out_as1802[0] vssd1 vssd1 vccd1 vccd1 _0607_/B2 sky130_fd_sc_hd__buf_1
XFILLER_0_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0671__A1 _0671_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_317_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0671__B2 _0671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output486_A _0741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_344_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0503_ hold76/X hold92/X vssd1 vssd1 vccd1 vccd1 _0767_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_238_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_280_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold19_A hold19/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_367_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0662__B2 _0662_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold320 _1106_/Q vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 hold342/A vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _0845_/X vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _1093_/Q vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold386 hold792/X vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _1084_/X vssd1 vssd1 vccd1 vccd1 _1085_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _0976_/Y vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 hold793/X vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_314_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0613__C _0613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0644__B2 _0644_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_372_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ _0983_/A _0983_/B _0983_/C _0983_/D vssd1 vssd1 vccd1 vccd1 _1017_/B sky130_fd_sc_hd__and4_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput414 _1117_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[30] sky130_fd_sc_hd__buf_12
Xoutput403 _1107_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[20] sky130_fd_sc_hd__buf_12
Xoutput425 _1241_/A vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput458 _1238_/A vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput469 _0609_/X vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
Xoutput436 _1251_/A vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__buf_12
Xoutput447 _1261_/A vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__buf_12
XFILLER_0_238_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0635__B2 _0635_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0635__A1 _0635_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_363_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_308_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_323_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold150 hold685/X vssd1 vssd1 vccd1 vccd1 _0789_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold194 hold696/X vssd1 vssd1 vccd1 vccd1 _1065_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _0932_/Y vssd1 vssd1 vccd1 vccd1 _0933_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold682/X vssd1 vssd1 vccd1 vccd1 _1098_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_244_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0626__B2 _0626_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_354_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output449_A hold89/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1251_ _1251_/A vssd1 vssd1 vccd1 vccd1 _1251_/X sky130_fd_sc_hd__buf_1
XFILLER_0_246_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1182_ _1184_/CLK _1182_/D vssd1 vssd1 vccd1 vccd1 _1182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_389_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_392_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_360_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0966_ _0956_/Y hold378/X _0965_/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0966_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_360_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0897_ _1085_/A _0897_/B vssd1 vssd1 vccd1 vccd1 _0897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_373_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_395_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_368_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0608__B2 _0608_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_336_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_386_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0820_ hold276/X _0840_/A2 _0819_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0820_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0751_ _0767_/A _0767_/B _0751_/C vssd1 vssd1 vccd1 vccd1 _0751_/X sky130_fd_sc_hd__and3_4
XFILLER_0_141_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output566_A hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0682_ _0682_/A1 _0746_/A2 _0746_/B1 _0682_/B2 vssd1 vssd1 vccd1 vccd1 _0685_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_367_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1234_ _1234_/A vssd1 vssd1 vccd1 vccd1 _1234_/X sky130_fd_sc_hd__buf_1
XFILLER_0_223_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1165_ _1224_/CLK _1165_/D vssd1 vssd1 vccd1 vccd1 _1165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_273_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1096_ _1224_/CLK _1096_/D vssd1 vssd1 vccd1 vccd1 _1096_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_392_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_365_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0949_ hold529/X _0952_/A2 _0952_/B1 _1078_/C _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0949_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout597_A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_324_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0621__C _0621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_292_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_292_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_374_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0803_ _0803_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0803_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0734_ _0734_/A1 _0746_/A2 _0518_/B _0734_/B2 vssd1 vssd1 vccd1 vccd1 _0737_/A sky130_fd_sc_hd__a22o_1
XANTENNA__0756__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 _0816_/X vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold705 _1208_/Q vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 _0882_/A vssd1 vssd1 vccd1 vccd1 _0772_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_295_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0665_ _0665_/A _0665_/B _0665_/C vssd1 vssd1 vccd1 vccd1 _0665_/X sky130_fd_sc_hd__or3_4
Xhold749 _1185_/Q vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 _1222_/Q vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0596_ input42/X _0598_/A2 _0598_/B1 input78/X vssd1 vssd1 vccd1 vccd1 _0596_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_283_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1217_ _1221_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _1217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1148_ _1154_/CLK _1148_/D vssd1 vssd1 vccd1 vccd1 _1148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_338_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1079_ _1078_/C _1078_/B hold322/X vssd1 vssd1 vccd1 vccd1 _1079_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0747__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_395_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_274_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput303 io_out_vliw[7] vssd1 vssd1 vccd1 vccd1 _0636_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_395_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_274_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput325 io_out_z80[27] vssd1 vssd1 vccd1 vccd1 _0714_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_227_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput314 io_out_z80[17] vssd1 vssd1 vccd1 vccd1 _0674_/A1 sky130_fd_sc_hd__buf_1
Xinput336 io_out_z80[4] vssd1 vssd1 vccd1 vccd1 _0622_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput347 hold694/X vssd1 vssd1 vccd1 vccd1 _0768_/B sky130_fd_sc_hd__clkbuf_1
Xinput369 hold510/X vssd1 vssd1 vccd1 vccd1 hold511/A sky130_fd_sc_hd__clkbuf_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput358 hold474/X vssd1 vssd1 vccd1 vccd1 hold475/A sky130_fd_sc_hd__clkbuf_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__buf_2
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_356_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output431_A _1247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1002_ _0799_/A _0996_/A hold549/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_254_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0807__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_335_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold502 hold502/A vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_303_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0717_ _0717_/A _0717_/B _0717_/C vssd1 vssd1 vccd1 vccd1 _0717_/X sky130_fd_sc_hd__or3_4
Xhold524 _0836_/X vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 hold599/X vssd1 vssd1 vccd1 vccd1 hold600/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 hold65/X vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_256_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold579 _1049_/Y vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _1027_/X vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _0879_/X vssd1 vssd1 vccd1 vccd1 _0880_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _1162_/Q vssd1 vssd1 vccd1 vccd1 _0983_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0648_ _0648_/A1 _0660_/A2 _0696_/B1 _0648_/B2 vssd1 vssd1 vccd1 vccd1 _0649_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_256_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0579_ _0579_/A1 _0590_/A2 _0604_/A2 input34/X vssd1 vssd1 vccd1 vccd1 _0579_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_256_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput111 io_oeb_z80[29] vssd1 vssd1 vccd1 vccd1 _0590_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput100 io_oeb_z80[19] vssd1 vssd1 vccd1 vccd1 _0568_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_274_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput122 io_oeb_z80[6] vssd1 vssd1 vccd1 vccd1 _0537_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput144 io_out_6502[26] vssd1 vssd1 vccd1 vccd1 _0711_/A1 sky130_fd_sc_hd__buf_2
Xinput133 io_out_6502[16] vssd1 vssd1 vccd1 vccd1 _0671_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput177 io_out_8x305[23] vssd1 vssd1 vccd1 vccd1 _0698_/B2 sky130_fd_sc_hd__buf_2
Xinput166 io_out_8x305[13] vssd1 vssd1 vccd1 vccd1 _0658_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput155 io_out_6502[3] vssd1 vssd1 vccd1 vccd1 _0619_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_355_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput188 io_out_8x305[33] vssd1 vssd1 vccd1 vccd1 _0738_/B2 sky130_fd_sc_hd__buf_2
Xinput199 io_out_as1802[10] vssd1 vssd1 vccd1 vccd1 _0647_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_291_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0671__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_325_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output479_A _0717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_340_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0502_ hold99/X _0517_/B vssd1 vssd1 vccd1 vccd1 _0505_/A sky130_fd_sc_hd__or2_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_265_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0895__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold310 hold398/X vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_376_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold343 hold76/X vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold716/X vssd1 vssd1 vccd1 vccd1 _1106_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold686/X vssd1 vssd1 vccd1 vccd1 _1093_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold387 hold782/X vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _1085_/X vssd1 vssd1 vccd1 vccd1 _1189_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _0846_/X vssd1 vssd1 vccd1 vccd1 _1120_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 hold754/X vssd1 vssd1 vccd1 vccd1 _1161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold398 hold736/X vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_271_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0886__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_279_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0810__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_322_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0982_ _0983_/C _0979_/B _0983_/D vssd1 vssd1 vccd1 vccd1 _0982_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput415 _1118_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[31] sky130_fd_sc_hd__buf_12
Xoutput404 _1108_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[21] sky130_fd_sc_hd__buf_12
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput426 _1242_/A vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__buf_12
XFILLER_0_285_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput459 _0641_/X vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
Xoutput437 _1252_/A vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__buf_12
Xoutput448 hold96/A vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__buf_12
XFILLER_0_238_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0635__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_311_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_304_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold162 hold92/X vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold151 hold560/X vssd1 vssd1 vccd1 vccd1 _1162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 hold550/X vssd1 vssd1 vccd1 vccd1 _1167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _0831_/X vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _0933_/Y vssd1 vssd1 vccd1 vccd1 _1147_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold385/X vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0571__A1 _0571_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout620 input342/X vssd1 vssd1 vccd1 vccd1 _1085_/A sky130_fd_sc_hd__buf_4
XFILLER_0_232_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0859__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1250_ _1250_/A vssd1 vssd1 vccd1 vccd1 _1250_/X sky130_fd_sc_hd__buf_1
XFILLER_0_235_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output511_A _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1181_ _1187_/CLK _1181_/D vssd1 vssd1 vccd1 vccd1 _1181_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_393_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0815__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0965_ _0965_/A _1021_/A vssd1 vssd1 vccd1 vccd1 _0965_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_360_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0896_ hold254/X _0880_/A _0895_/X vssd1 vssd1 vccd1 vccd1 _0896_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0709__C _0709_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_368_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_322_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0750_ input1/X _1087_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0751_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_141_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output461_A _0649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0681_ _0681_/A _0681_/B _0681_/C vssd1 vssd1 vccd1 vccd1 _0681_/X sky130_fd_sc_hd__or3_4
XANTENNA_output559_A hold185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0535__A1 _0535_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1233_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1233_/X sky130_fd_sc_hd__buf_1
XFILLER_0_223_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0838__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1164_ _1225_/CLK _1164_/D vssd1 vssd1 vccd1 vccd1 _1164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_273_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1095_ _1225_/CLK _1095_/D vssd1 vssd1 vccd1 vccd1 _1095_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_392_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_373_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0948_ _1036_/A _0948_/B vssd1 vssd1 vccd1 vccd1 _0948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_368_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0879_ hold212/X _0776_/A hold605/A _0983_/D vssd1 vssd1 vccd1 vccd1 _0879_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0802_ hold227/X _0810_/A2 _0801_/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0802_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0733_ _0733_/A _0733_/B _0733_/C vssd1 vssd1 vccd1 vccd1 _0733_/X sky130_fd_sc_hd__or3_4
Xhold717 _1110_/Q vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 _0814_/X vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold728 _0772_/X vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0664_ _0664_/A1 _0732_/A2 _0696_/B1 _0664_/B2 vssd1 vssd1 vccd1 vccd1 _0665_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_268_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold739 _1084_/S vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_283_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0595_ _0595_/A1 _0605_/A2 _0593_/X _0594_/X vssd1 vssd1 vccd1 vccd1 _1261_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_236_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1216_ _1221_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 _1216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1147_ _1154_/CLK _1147_/D vssd1 vssd1 vccd1 vccd1 _1147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1078_ hold322/X _1078_/B _1078_/C vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0747__A1 _0747_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0747__B2 _0747_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput304 io_out_vliw[8] vssd1 vssd1 vccd1 vccd1 _0640_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_328_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput326 io_out_z80[28] vssd1 vssd1 vccd1 vccd1 _0718_/A1 sky130_fd_sc_hd__buf_1
Xinput315 io_out_z80[18] vssd1 vssd1 vccd1 vccd1 _0678_/A1 sky130_fd_sc_hd__buf_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput337 io_out_z80[5] vssd1 vssd1 vccd1 vccd1 _0626_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput359 hold429/X vssd1 vssd1 vccd1 vccd1 hold430/A sky130_fd_sc_hd__clkbuf_1
Xinput348 hold435/X vssd1 vssd1 vccd1 vccd1 hold436/A sky130_fd_sc_hd__clkbuf_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold88 hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__buf_4
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__buf_2
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0683__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_371_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0738__A1 _0738_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0738__B2 _0738_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_292_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_292_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output424_A _1240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_379_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1001_ hold548/X _1008_/C _0996_/A vssd1 vssd1 vccd1 vccd1 _1001_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_347_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_390_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_350_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0823__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0716_ _0716_/A1 _0508_/B _0748_/B1 _0716_/B2 vssd1 vssd1 vccd1 vccd1 _0717_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_279_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold525 _1118_/Q vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _0968_/Y vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _0880_/X vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _0978_/Y vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 hold759/X vssd1 vssd1 vccd1 vccd1 _0999_/D sky130_fd_sc_hd__buf_1
XFILLER_0_268_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0647_ _0647_/A1 _0514_/B _0695_/B1 _0647_/B2 vssd1 vssd1 vccd1 vccd1 _0649_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0578_ input69/X _0586_/B1 _0574_/X _0577_/X vssd1 vssd1 vccd1 vccd1 _1254_/A sky130_fd_sc_hd__a211o_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_381_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_314_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0717__C _0717_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_353_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_274_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput101 io_oeb_z80[1] vssd1 vssd1 vccd1 vccd1 _0525_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput123 io_oeb_z80[7] vssd1 vssd1 vccd1 vccd1 _0539_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput112 io_oeb_z80[2] vssd1 vssd1 vccd1 vccd1 _0528_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput145 io_out_6502[27] vssd1 vssd1 vccd1 vccd1 _0715_/A1 sky130_fd_sc_hd__buf_2
Xinput134 io_out_6502[17] vssd1 vssd1 vccd1 vccd1 _0675_/A1 sky130_fd_sc_hd__buf_2
Xinput178 io_out_8x305[24] vssd1 vssd1 vccd1 vccd1 _0702_/B2 sky130_fd_sc_hd__buf_2
Xinput167 io_out_8x305[14] vssd1 vssd1 vccd1 vccd1 _0662_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput156 io_out_6502[4] vssd1 vssd1 vccd1 vccd1 _0623_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput189 io_out_8x305[34] vssd1 vssd1 vccd1 vccd1 _0742_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_291_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_371_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0501_ _1267_/A hold647/X _0852_/A vssd1 vssd1 vccd1 vccd1 _0518_/A sky130_fd_sc_hd__mux2_8
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1180_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA_output541_A hold252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_253_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0512__C_N _0868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_367_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0647__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_382_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold300 hold712/X vssd1 vssd1 vccd1 vccd1 _1104_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _0878_/X vssd1 vssd1 vccd1 vccd1 _1129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold322 _1187_/Q vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 hold650/X vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold344 hold743/X vssd1 vssd1 vccd1 vccd1 _0845_/A sky130_fd_sc_hd__buf_1
XFILLER_0_376_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0583__C1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold377 hold689/X vssd1 vssd1 vccd1 vccd1 _0967_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold355 hold724/X vssd1 vssd1 vccd1 vccd1 _0849_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold366 hold726/X vssd1 vssd1 vccd1 vccd1 _0882_/A sky130_fd_sc_hd__buf_1
XFILLER_0_256_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold388 hold786/X vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 hold794/X vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_271_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_325_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_314_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_364_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0981_ _0789_/A _1021_/A hold559/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0981_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output491_A _0621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput405 _1109_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[22] sky130_fd_sc_hd__buf_12
Xoutput416 _1090_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[3] sky130_fd_sc_hd__buf_12
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput427 _1243_/A vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput438 _1253_/A vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__buf_12
Xoutput449 hold89/A vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__buf_12
XFILLER_0_281_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_293_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold141 hold713/X vssd1 vssd1 vccd1 vccd1 _0817_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 hold711/X vssd1 vssd1 vccd1 vccd1 _0811_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold589/X vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold163 hold699/X vssd1 vssd1 vccd1 vccd1 _1076_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold386/X vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__clkbuf_2
Xhold174 _0929_/Y vssd1 vssd1 vccd1 vccd1 _0930_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0571__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 hold522/X vssd1 vssd1 vccd1 vccd1 _1114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 hold604/X vssd1 vssd1 vccd1 vccd1 hold605/A sky130_fd_sc_hd__buf_4
XFILLER_0_217_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1180_ _1180_/CLK _1180_/D vssd1 vssd1 vccd1 vccd1 _1180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_389_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_246_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0964_ _0967_/C _0964_/B vssd1 vssd1 vccd1 vccd1 _0964_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0831__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0786__C1 _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0895_ hold227/X _0776_/A hold605/A _1004_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0895_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_383_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_322_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0792__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_299_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_302_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0680_ _0680_/A1 _0732_/A2 _0696_/B1 _0680_/B2 vssd1 vssd1 vccd1 vccd1 _0681_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_153_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output454_A _1234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0535__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1232_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1232_/X sky130_fd_sc_hd__buf_1
XANTENNA__0940__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1163_ _1225_/CLK _1163_/D vssd1 vssd1 vccd1 vccd1 _1163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_255_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1094_ _1225_/CLK _1094_/D vssd1 vssd1 vccd1 vccd1 _1094_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_365_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_380_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0947_ hold217/X _0953_/A2 _0946_/X vssd1 vssd1 vccd1 vccd1 _0947_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_286_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0878_ hold310/X hold729/A hold607/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0878_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1184_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_294_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_347_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_362_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output571_A hold280/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0801_ _0801_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0801_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0732_ _0732_/A1 _0732_/A2 _0748_/B1 _0732_/B2 vssd1 vssd1 vccd1 vccd1 _0733_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_268_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold718 _0824_/X vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold707 _1211_/Q vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0663_ _0663_/A1 _0514_/B _0683_/B1 _0663_/B2 vssd1 vssd1 vccd1 vccd1 _0665_/B sky130_fd_sc_hd__a22o_1
Xhold729 hold729/A vssd1 vssd1 vccd1 vccd1 _0774_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0594_ input41/X _0604_/A2 _0510_/B input77/X vssd1 vssd1 vccd1 vccd1 _0594_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_372_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1215_ _1215_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 _1215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1146_ _1154_/CLK _1146_/D vssd1 vssd1 vccd1 vccd1 _1146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_370_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0692__B2 _0692_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1077_ _0956_/Y hold284/X _1076_/X _0500_/Y vssd1 vssd1 vccd1 vccd1 _1077_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_365_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_361_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput305 io_out_vliw[9] vssd1 vssd1 vccd1 vccd1 _0644_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_328_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput327 io_out_z80[29] vssd1 vssd1 vccd1 vccd1 _0722_/A1 sky130_fd_sc_hd__buf_1
Xinput316 io_out_z80[19] vssd1 vssd1 vccd1 vccd1 _0682_/A1 sky130_fd_sc_hd__buf_1
XANTENNA__0904__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_328_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput338 io_out_z80[6] vssd1 vssd1 vccd1 vccd1 _0630_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput349 hold444/X vssd1 vssd1 vccd1 vccd1 hold445/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_242_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__buf_1
XFILLER_0_199_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_344_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0683__A1 _0683_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0683__B2 _0683_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_344_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0986__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_9 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_369_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1000_ _1017_/A _1017_/B _1017_/C vssd1 vssd1 vccd1 vccd1 _1008_/C sky130_fd_sc_hd__and3_1
XFILLER_0_344_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_387_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0674__B2 _0674_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0977__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0715_ _0715_/A1 _0593_/A _0516_/B _0715_/B2 vssd1 vssd1 vccd1 vccd1 _0717_/B sky130_fd_sc_hd__a22o_1
Xhold526 _0840_/X vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 hold61/X vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold537 _0969_/Y vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold559 _0980_/X vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _0998_/Y vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0646_ _0646_/A1 _0506_/B _0526_/A _0646_/B2 vssd1 vssd1 vccd1 vccd1 _0649_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0577_ _0577_/A1 _0590_/A2 _0604_/A2 input33/X vssd1 vssd1 vccd1 vccd1 _0577_/X sky130_fd_sc_hd__a22o_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_295_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1129_ _1157_/CLK _1129_/D vssd1 vssd1 vccd1 vccd1 _1129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_326_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_353_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout615_A _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_275_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput102 io_oeb_z80[20] vssd1 vssd1 vccd1 vccd1 _0571_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_274_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput113 io_oeb_z80[30] vssd1 vssd1 vccd1 vccd1 _0595_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput124 io_oeb_z80[8] vssd1 vssd1 vccd1 vccd1 _0541_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput135 io_out_6502[18] vssd1 vssd1 vccd1 vccd1 _0679_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput168 io_out_8x305[15] vssd1 vssd1 vccd1 vccd1 _0666_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput146 io_out_6502[28] vssd1 vssd1 vccd1 vccd1 _0719_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput157 io_out_6502[5] vssd1 vssd1 vccd1 vccd1 _0627_/A1 sky130_fd_sc_hd__buf_2
Xinput179 io_out_8x305[25] vssd1 vssd1 vccd1 vccd1 _0706_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_291_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0656__B2 _0656_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0959__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_325_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1081__A1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0500_ _1085_/A vssd1 vssd1 vccd1 vccd1 _0500_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_265_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output534_A _0514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0647__B2 _0647_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0647__A1 _0647_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_390_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_390_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold301 hold409/X vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold323 _1079_/Y vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 hold719/X vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _0786_/X vssd1 vssd1 vccd1 vccd1 _1091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _0849_/X vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 hold728/X vssd1 vssd1 vccd1 vccd1 hold729/A sky130_fd_sc_hd__buf_2
Xhold345 hold538/X vssd1 vssd1 vccd1 vccd1 _1159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _0964_/Y vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0629_ _0629_/A _0629_/B _0629_/C vssd1 vssd1 vccd1 vccd1 _0629_/X sky130_fd_sc_hd__or3_4
Xhold389 hold784/X vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_271_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_325_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0638__B2 _0638_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_366_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_366_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_251_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0980_ hold558/X _0979_/X _0956_/Y vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_372_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output484_A _0733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput406 _1110_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[23] sky130_fd_sc_hd__buf_12
Xoutput417 _1091_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[4] sky130_fd_sc_hd__buf_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput428 _1244_/A vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput439 _1254_/A vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_0_238_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0829__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_348_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_304_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold131 hold700/X vssd1 vssd1 vccd1 vccd1 _0833_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold542/X vssd1 vssd1 vccd1 vccd1 _1176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold546/X vssd1 vssd1 vccd1 vccd1 _1173_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold120 hold564/X vssd1 vssd1 vccd1 vccd1 hold565/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _0837_/X vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _0938_/Y vssd1 vssd1 vccd1 vccd1 _0939_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _0930_/Y vssd1 vssd1 vccd1 vccd1 _1146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 hold82/X vssd1 vssd1 vccd1 vccd1 _0598_/B1 sky130_fd_sc_hd__buf_2
XFILLER_0_217_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout611 _0851_/X vssd1 vssd1 vccd1 vccd1 _0952_/B1 sky130_fd_sc_hd__buf_4
Xhold197 hold405/X vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_336_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0859__A1 hold220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold260_A _1100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0755__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_386_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_322_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_282_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_377_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_377_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0963_ _0779_/A _1021_/A hold635/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0894_ _1085_/A _0894_/B vssd1 vssd1 vccd1 vccd1 _0894_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0710__B1 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_395_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_395_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_383_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_336_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_304_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_386_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_359_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output447_A _1261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1231_ hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__buf_1
X_1162_ _1167_/CLK _1162_/D vssd1 vssd1 vccd1 vccd1 _1162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1093_ _1167_/CLK _1093_/D vssd1 vssd1 vccd1 vccd1 _1093_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_365_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0842__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0946_ hold523/X _0952_/A2 _0952_/B1 _1072_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0946_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_333_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0877_ _0880_/A _0877_/B vssd1 vssd1 vccd1 vccd1 _0877_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_289_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_347_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0989__B1 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output397_A _1102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0800_ hold171/X _0810_/A2 _0799_/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0800_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_370_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0731_ _0731_/A1 _0747_/A2 _0516_/B _0731_/B2 vssd1 vssd1 vccd1 vccd1 _0733_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_268_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output564_A hold229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold708 _0820_/X vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 _1092_/Q vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_268_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0662_ _0662_/A1 _0674_/A2 _0674_/B1 _0662_/B2 vssd1 vssd1 vccd1 vccd1 _0665_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0593_ _0593_/A hold95/A vssd1 vssd1 vccd1 vccd1 _0593_/X sky130_fd_sc_hd__or2_2
XFILLER_0_228_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0837__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1214_ _1214_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 _1214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ _1154_/CLK _1145_/D vssd1 vssd1 vccd1 vccd1 _1145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1076_ _1076_/A _1076_/B vssd1 vssd1 vccd1 vccd1 _1076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0929_ hold173/X _0953_/A2 _0928_/X vssd1 vssd1 vccd1 vccd1 _0929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_395_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_286_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout595_A _0515_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput317 io_out_z80[1] vssd1 vssd1 vccd1 vccd1 _0610_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput306 io_out_z80[0] vssd1 vssd1 vccd1 vccd1 _0606_/A1 sky130_fd_sc_hd__clkbuf_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput339 io_out_z80[7] vssd1 vssd1 vccd1 vccd1 _0634_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput328 io_out_z80[2] vssd1 vssd1 vccd1 vccd1 _0614_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_344_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0763__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_371_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_265_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_280_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_343_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_303_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0714_ _0714_/A1 _0505_/Y _0746_/B1 _0714_/B2 vssd1 vssd1 vccd1 vccd1 _0717_/A sky130_fd_sc_hd__a22o_1
Xhold527 _1112_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 hold69/X vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_268_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0645_ _0645_/A _0645_/B _0645_/C vssd1 vssd1 vccd1 vccd1 _0645_/X sky130_fd_sc_hd__or3_4
Xhold538 _0970_/X vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 _1001_/Y vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0576_ input68/X _0586_/B1 _0574_/X _0575_/X vssd1 vssd1 vccd1 vccd1 _1253_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_110_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_295_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0898__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1128_ _1175_/CLK _1128_/D vssd1 vssd1 vccd1 vccd1 _1128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1059_ _0956_/Y hold327/X _1058_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _1059_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_334_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_247_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput114 io_oeb_z80[31] vssd1 vssd1 vccd1 vccd1 _0597_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput103 io_oeb_z80[21] vssd1 vssd1 vccd1 vccd1 _0573_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_255_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput125 io_oeb_z80[9] vssd1 vssd1 vccd1 vccd1 _0543_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__0889__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput136 io_out_6502[19] vssd1 vssd1 vccd1 vccd1 _0683_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput169 io_out_8x305[16] vssd1 vssd1 vccd1 vccd1 _0670_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput147 io_out_6502[29] vssd1 vssd1 vccd1 vccd1 _0723_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput158 io_out_6502[6] vssd1 vssd1 vccd1 vccd1 _0631_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_371_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_369_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_261_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0647__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_390_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_390_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0804__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold302 hold730/X vssd1 vssd1 vccd1 vccd1 _1127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold324 hold656/X vssd1 vssd1 vccd1 vccd1 _1187_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 hold720/X vssd1 vssd1 vccd1 vccd1 _1092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold676/X vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0583__A1 _0583_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold357 _0850_/X vssd1 vssd1 vccd1 vccd1 _1122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 hold742/X vssd1 vssd1 vccd1 vccd1 _1082_/B sky130_fd_sc_hd__buf_2
Xhold346 hold626/X vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0628_ _0628_/A1 _0660_/A2 _0628_/B1 _0628_/B2 vssd1 vssd1 vccd1 vccd1 _0629_/C sky130_fd_sc_hd__a22o_2
Xhold379 _0966_/X vssd1 vssd1 vccd1 vccd1 _1158_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0559_ _0565_/A _0559_/B _0559_/C vssd1 vssd1 vccd1 vccd1 _1247_/A sky130_fd_sc_hd__or3_4
XFILLER_0_244_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_271_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1063__A2 _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0810__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0574__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_243_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_317_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_372_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_372_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output477_A _0709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput407 _1111_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[24] sky130_fd_sc_hd__buf_12
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput418 _1092_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[5] sky130_fd_sc_hd__buf_12
Xoutput429 _1245_/A vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__buf_12
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_292_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_304_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold110 hold112/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0556__A1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 hold556/X vssd1 vssd1 vccd1 vccd1 _1184_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold715/X vssd1 vssd1 vccd1 vccd1 _0815_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold662/X vssd1 vssd1 vccd1 vccd1 _0797_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold530/X vssd1 vssd1 vccd1 vccd1 _1117_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold380/X vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__clkbuf_2
Xhold154 hold657/X vssd1 vssd1 vccd1 vccd1 _0825_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout601 _0628_/B1 vssd1 vssd1 vccd1 vccd1 _0696_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_229_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold187 _0939_/Y vssd1 vssd1 vccd1 vccd1 _1149_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _0908_/Y vssd1 vssd1 vccd1 vccd1 _0909_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _0775_/A vssd1 vssd1 vccd1 vccd1 _0776_/A sky130_fd_sc_hd__buf_4
XFILLER_0_336_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0755__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_354_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0649__C _0649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0962_ hold634/X _0961_/X _0956_/Y vssd1 vssd1 vccd1 vccd1 _0962_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0893_ hold303/X _0880_/A hold760/X vssd1 vssd1 vccd1 vccd1 _0893_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_266_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0710__B2 _0710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_383_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_336_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0529__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_272_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1161_ _1167_/CLK _1161_/D vssd1 vssd1 vccd1 vccd1 _1161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_377_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1092_ _1175_/CLK _1092_/D vssd1 vssd1 vccd1 vccd1 _1092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_380_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0945_ _1036_/A _0945_/B vssd1 vssd1 vccd1 vccd1 _0945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0876_ hold331/X _0776_/A hold605/A _0983_/C vssd1 vssd1 vccd1 vccd1 _0876_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_254_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_368_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0695__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_362_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ _0730_/A1 _0746_/A2 _0746_/B1 _0730_/B2 vssd1 vssd1 vccd1 vccd1 _0733_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold709 _1216_/Q vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_268_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0661_ _0661_/A _0661_/B _0661_/C vssd1 vssd1 vccd1 vccd1 _0661_/X sky130_fd_sc_hd__or3_4
XANTENNA_output557_A hold182/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_283_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0592_ _0592_/A _0592_/B _0515_/B vssd1 vssd1 vccd1 vccd1 _0592_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_283_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1213_ _1215_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 _1213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1144_ _1154_/CLK _1144_/D vssd1 vssd1 vccd1 vccd1 _1144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1075_ _1078_/C _1078_/B vssd1 vssd1 vccd1 vccd1 _1075_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0601__B1 hold95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0928_ hold248/X _0952_/A2 _0952_/B1 _1050_/C _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0928_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0859_ hold220/X hold729/A hold645/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0859_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_286_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput318 io_out_z80[20] vssd1 vssd1 vccd1 vccd1 _0686_/A1 sky130_fd_sc_hd__buf_1
Xinput307 io_out_z80[10] vssd1 vssd1 vccd1 vccd1 _0646_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_328_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput329 io_out_z80[30] vssd1 vssd1 vccd1 vccd1 _0726_/A1 sky130_fd_sc_hd__buf_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_384_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_344_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0763__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_360_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_360_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_265_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_273_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0657__C _0657_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0659__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_394_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0954__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_362_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0713_ _0713_/A _0713_/B _0713_/C vssd1 vssd1 vccd1 vccd1 _0713_/X sky130_fd_sc_hd__or3_4
Xhold517 hold517/A vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0644_ _0644_/A1 _0660_/A2 _0696_/B1 _0644_/B2 vssd1 vssd1 vccd1 vccd1 _0645_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_268_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold528 _0828_/X vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 hold755/X vssd1 vssd1 vccd1 vccd1 _1038_/A sky130_fd_sc_hd__buf_1
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_283_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0575_ _0575_/A1 _0590_/A2 _0604_/A2 input32/X vssd1 vssd1 vccd1 vccd1 _0575_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1127_ _1189_/CLK _1127_/D vssd1 vssd1 vccd1 vccd1 _1127_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0864__A hold99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1058_ _1058_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_247_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput115 io_oeb_z80[32] vssd1 vssd1 vccd1 vccd1 _0599_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput104 io_oeb_z80[22] vssd1 vssd1 vccd1 vccd1 _0575_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput126 io_out_6502[0] vssd1 vssd1 vccd1 vccd1 _0607_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_355_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput137 io_out_6502[1] vssd1 vssd1 vccd1 vccd1 _0611_/A1 sky130_fd_sc_hd__buf_2
Xinput148 io_out_6502[2] vssd1 vssd1 vccd1 vccd1 _0615_/A1 sky130_fd_sc_hd__buf_2
Xinput159 io_out_6502[7] vssd1 vssd1 vccd1 vccd1 _0635_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_270_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_344_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output422_A _1096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_300_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold314 hold702/X vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 hold765/X vssd1 vssd1 vccd1 vccd1 _1060_/A sky130_fd_sc_hd__buf_1
XFILLER_0_142_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold303 hold401/X vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold369 _0847_/X vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _0780_/X vssd1 vssd1 vccd1 vccd1 _1088_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 hold627/X vssd1 vssd1 vccd1 vccd1 _1087_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold358 hold722/X vssd1 vssd1 vccd1 vccd1 _0847_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_229_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0627_ _0627_/A1 _0514_/B _0695_/B1 _0627_/B2 vssd1 vssd1 vccd1 vccd1 _0629_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0558_ input97/X _0590_/A2 _0510_/B input61/X vssd1 vssd1 vccd1 vccd1 _0559_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_252_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_366_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout620_A input342/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0574__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_251_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput408 _1112_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[25] sky130_fd_sc_hd__buf_12
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput419 _1093_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[6] sky130_fd_sc_hd__buf_12
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0970__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0845__C _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_363_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 _0507_/X vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__buf_2
XFILLER_0_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold144 _1035_/Y vssd1 vssd1 vccd1 vccd1 _1036_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _0769_/X vssd1 vssd1 vccd1 vccd1 _1086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 hold625/X vssd1 vssd1 vccd1 vccd1 _1166_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold666/X vssd1 vssd1 vccd1 vccd1 _0805_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold155 hold658/X vssd1 vssd1 vccd1 vccd1 _1180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _0923_/Y vssd1 vssd1 vccd1 vccd1 _0924_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold771/X vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__buf_1
Xfanout602 _0628_/B1 vssd1 vssd1 vccd1 vccd1 _0748_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold188 hold387/X vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__clkbuf_2
Xfanout613 _0775_/A vssd1 vssd1 vccd1 vccd1 _0952_/A2 sky130_fd_sc_hd__buf_4
Xhold199 _0909_/Y vssd1 vssd1 vccd1 vccd1 _1139_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1214_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_394_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_314_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_322_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0499__A _0860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0952__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_243_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0665__C _0665_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_392_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ _0967_/A _0961_/B vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_298_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0786__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0892_ hold171/X _0776_/A hold605/A _0999_/D _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0892_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_301_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_298_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0943__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0856__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0710__A2 _0505_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_383_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0872__A hold76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0529__A2 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_272_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_327_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1160_ _1225_/CLK _1160_/D vssd1 vssd1 vccd1 vccd1 _1160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1091_ _1175_/CLK _1091_/D vssd1 vssd1 vccd1 vccd1 _1091_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_377_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_365_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0944_ hold188/X _0953_/A2 _0943_/X vssd1 vssd1 vccd1 vccd1 _0944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0875_ hold272/X hold729/A hold693/X _0500_/Y vssd1 vssd1 vccd1 vccd1 _0875_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_125_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0695__A1 _0695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0695__B2 _0695_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_383_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_358_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0907__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_374_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0686__B2 _0686_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_347_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0610__B2 _0610_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0660_ _0660_/A1 _0660_/A2 _0696_/B1 _0660_/B2 vssd1 vssd1 vccd1 vccd1 _0661_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0591_ input75/X hold82/X hold95/X vssd1 vssd1 vccd1 vccd1 _0592_/B sky130_fd_sc_hd__a21o_1
XANTENNA_output452_A _1266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1212_ _1215_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 _1212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_284_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1143_ _1189_/CLK _1143_/D vssd1 vssd1 vccd1 vccd1 _1143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_338_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1074_ _0956_/Y hold287/X _1073_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1074_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_365_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ _1036_/A _0927_/B vssd1 vssd1 vccd1 vccd1 _0927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0601__A1 _0601_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0858_ _0880_/A _0858_/B vssd1 vssd1 vccd1 vccd1 _0858_/X sky130_fd_sc_hd__or2_1
XFILLER_0_395_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0789_ _0789_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0789_/X sky130_fd_sc_hd__or2_1
XFILLER_0_286_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput308 io_out_z80[11] vssd1 vssd1 vccd1 vccd1 _0650_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput319 io_out_z80[21] vssd1 vssd1 vccd1 vccd1 _0690_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0668__B2 _0668_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_360_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_385_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0659__A1 _0659_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0659__B2 _0659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_387_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0673__C _0673_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_270_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0712_ _0712_/A1 _0508_/B _0748_/B1 _0712_/B2 vssd1 vssd1 vccd1 vccd1 _0713_/C sky130_fd_sc_hd__a22o_1
Xhold518 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 hold63/X vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_268_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0643_ _0643_/A1 _0514_/B _0695_/B1 _0643_/B2 vssd1 vssd1 vccd1 vccd1 _0645_/B sky130_fd_sc_hd__a22o_1
Xhold529 _1117_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_283_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0574_ input11/X _0593_/A _0526_/X vssd1 vssd1 vccd1 vccd1 _0574_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_148_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1221_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_378_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1126_ _1157_/CLK _1126_/D vssd1 vssd1 vccd1 vccd1 _1126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0864__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1057_ _1181_/Q _1057_/B vssd1 vssd1 vccd1 vccd1 _1057_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_381_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_319_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_334_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput116 io_oeb_z80[33] vssd1 vssd1 vccd1 vccd1 _0601_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput105 io_oeb_z80[23] vssd1 vssd1 vccd1 vccd1 _0577_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_255_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput127 io_out_6502[10] vssd1 vssd1 vccd1 vccd1 _0647_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_355_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput149 io_out_6502[30] vssd1 vssd1 vccd1 vccd1 _0727_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput138 io_out_6502[20] vssd1 vssd1 vccd1 vccd1 _0687_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_270_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_369_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_384_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1066__A1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_337_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_297_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0501__A0 _1267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_363_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold315 _0826_/X vssd1 vssd1 vccd1 vccd1 _1111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _1054_/Y vssd1 vssd1 vccd1 vccd1 _1057_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _0893_/Y vssd1 vssd1 vccd1 vccd1 _0894_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold337 hold664/X vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 hold723/X vssd1 vssd1 vccd1 vccd1 _0965_/A sky130_fd_sc_hd__buf_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold359 hold641/X vssd1 vssd1 vccd1 vccd1 _1160_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0626_ _0626_/A1 _0674_/A2 _0674_/B1 _0626_/B2 vssd1 vssd1 vccd1 vccd1 _0629_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_159_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0557_ input25/X hold100/X _0518_/B input13/X vssd1 vssd1 vccd1 vccd1 _0559_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_244_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1109_ _1221_/CLK _1109_/D vssd1 vssd1 vccd1 vccd1 _1109_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_366_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout613_A _0775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_334_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_366_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0731__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_382_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_382_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput409 _1113_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[26] sky130_fd_sc_hd__buf_12
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_276_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_348_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_348_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold101 _0600_/X vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold112 _1086_/Q vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold585/X vssd1 vssd1 vccd1 vccd1 _1170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold670/X vssd1 vssd1 vccd1 vccd1 _0801_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold145 _1036_/Y vssd1 vssd1 vccd1 vccd1 _1175_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold705/X vssd1 vssd1 vccd1 vccd1 _0813_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold684/X vssd1 vssd1 vccd1 vccd1 _1096_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_284_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout603 _0510_/B vssd1 vssd1 vccd1 vccd1 _0628_/B1 sky130_fd_sc_hd__buf_2
X_0609_ _0609_/A _0609_/B _0609_/C vssd1 vssd1 vccd1 vccd1 _0609_/X sky130_fd_sc_hd__or3_4
XFILLER_0_229_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold189 _0944_/Y vssd1 vssd1 vccd1 vccd1 _0945_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _0924_/Y vssd1 vssd1 vccd1 vccd1 _1144_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _0966_/C1 vssd1 vssd1 vccd1 vccd1 _1006_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_244_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold775_A _1098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold690 _0862_/X vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_290_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_290_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0681__C _0681_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0960_ _0967_/A _0961_/B vssd1 vssd1 vccd1 vccd1 _0964_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_345_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output482_A _0725_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0891_ _1085_/A _0891_/B vssd1 vssd1 vccd1 vccd1 _0891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_395_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0872__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0934__B1 _0851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_272_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_359_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_263_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_377_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ _1188_/CLK _1090_/D vssd1 vssd1 vccd1 vccd1 _1090_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_333_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0943_ hold278/X _0952_/A2 _0952_/B1 _1071_/B _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0943_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0874_ _0880_/A _0874_/B vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__or2_1
XFILLER_0_301_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_333_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_364_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput570 hold316/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_245_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0777__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_374_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_390_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0590_ _0590_/A1 _0590_/A2 _0604_/A2 input39/X vssd1 vssd1 vccd1 vccd1 _0592_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output445_A hold78/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_291_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1211_ _1215_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 _1211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_251_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1142_ _1189_/CLK _1142_/D vssd1 vssd1 vccd1 vccd1 _1142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1073_ _1073_/A _1076_/B vssd1 vssd1 vccd1 vccd1 _1073_/X sky130_fd_sc_hd__or2_1
XFILLER_0_365_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_346_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0926_ hold269/X _0953_/A2 _0925_/X vssd1 vssd1 vccd1 vccd1 _0926_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0857_ hold335/X _0776_/A hold605/A _0961_/B _0856_/X vssd1 vssd1 vccd1 vccd1 _0857_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0788_ hold312/X _0840_/A2 _0787_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput309 io_out_z80[12] vssd1 vssd1 vccd1 vccd1 _0654_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_360_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0840__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_273_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0659__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output395_A _1100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0711_ _0711_/A1 _0593_/A _0516_/B _0711_/B2 vssd1 vssd1 vccd1 vccd1 _0713_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_154_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0595__A1 _0595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output562_A hold217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 hold508/A vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0642_ _0642_/A1 _0674_/A2 _0674_/B1 _0642_/B2 vssd1 vssd1 vccd1 vccd1 _0645_/A sky130_fd_sc_hd__a22o_1
Xhold519 hold71/X vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_256_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0573_ _0573_/A1 _0506_/B _0569_/A _0572_/X vssd1 vssd1 vccd1 vccd1 _1252_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_283_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_363_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1125_ _1189_/CLK _1125_/D vssd1 vssd1 vccd1 vccd1 _1125_/Q sky130_fd_sc_hd__dfxtp_1
X_1056_ _0825_/A _1080_/B _1055_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _1056_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_334_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0586__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0909_ _1036_/A _0909_/B vssd1 vssd1 vccd1 vccd1 _0909_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout593_A _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput117 io_oeb_z80[34] vssd1 vssd1 vccd1 vccd1 _0603_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput106 io_oeb_z80[24] vssd1 vssd1 vccd1 vccd1 _0579_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_355_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_255_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput139 io_out_6502[21] vssd1 vssd1 vccd1 vccd1 _0691_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput128 io_out_6502[11] vssd1 vssd1 vccd1 vccd1 _0651_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_215_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1232__A _1232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_384_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0577__A1 _0577_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_90 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0804__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_316_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0568__A1 _0568_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 _0894_/Y vssd1 vssd1 vccd1 vccd1 _1134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 hold402/X vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0625_ _0625_/A _0625_/B _0625_/C vssd1 vssd1 vccd1 vccd1 _0625_/X sky130_fd_sc_hd__or3_4
Xhold327 _1057_/Y vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _0843_/X vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold665/X vssd1 vssd1 vccd1 vccd1 _1089_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0556_ input96/X _0590_/A2 _0565_/A _0555_/X vssd1 vssd1 vccd1 vccd1 _1246_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_252_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0740__B2 _0740_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1108_ _1214_/CLK _1108_/D vssd1 vssd1 vccd1 vccd1 _1108_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_366_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1039_ _1080_/B _1039_/B vssd1 vssd1 vccd1 vccd1 _1039_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__0891__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_A hold100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_247_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0731__B2 _0731_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0731__A1 _0731_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0785__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_382_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_382_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0722__B2 _0722_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_292_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 _0601_/X vssd1 vssd1 vccd1 vccd1 _1264_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold135 hold709/X vssd1 vssd1 vccd1 vccd1 _0829_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 _0955_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold620/X vssd1 vssd1 vccd1 vccd1 hold621/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold157 hold577/X vssd1 vssd1 vccd1 vccd1 _1174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold703/X vssd1 vssd1 vccd1 vccd1 _1058_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hold672/X vssd1 vssd1 vccd1 vccd1 _0807_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0608_ _0608_/A1 _0660_/A2 _0628_/B1 _0608_/B2 vssd1 vssd1 vccd1 vccd1 _0609_/C sky130_fd_sc_hd__a22o_1
Xfanout604 hold82/X vssd1 vssd1 vccd1 vccd1 _0510_/B sky130_fd_sc_hd__buf_4
Xhold179 hold381/X vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__clkbuf_2
Xfanout615 _0966_/C1 vssd1 vssd1 vccd1 vccd1 _1083_/C1 sky130_fd_sc_hd__buf_4
X_0539_ _0539_/A1 _0605_/A2 _0529_/X _0538_/X vssd1 vssd1 vccd1 vccd1 _1238_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_379_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold680 _0792_/X vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _1161_/Q vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0704__B2 _0704_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0890_ hold291/X _0880_/A _0889_/X vssd1 vssd1 vccd1 vccd1 _0890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output475_A _0701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_395_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0631__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_304_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1240__A _1240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_388_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0942_ _1036_/A _0942_/B vssd1 vssd1 vccd1 vccd1 _0942_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_144_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0873_ hold312/X _0952_/A2 _0952_/B1 _0983_/B _0872_/X vssd1 vssd1 vccd1 vccd1 _0873_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_301_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_391_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0604__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_277_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput560 hold203/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput571 hold280/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_12
XANTENNA__1235__A _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_374_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_359_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0793__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_390_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output438_A _1253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1210_ _1215_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 _1210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_291_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_284_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1141_ _1189_/CLK _1141_/D vssd1 vssd1 vccd1 vccd1 _1141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_260_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1072_ _1072_/A _1072_/B vssd1 vssd1 vccd1 vccd1 _1072_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_180 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_380_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0925_ hold235/X _0952_/A2 _0952_/B1 _1050_/B _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0925_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0856_ hold73/X _1082_/C vssd1 vssd1 vccd1 vccd1 _0856_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0787_ _0849_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0787_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_267_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_388_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0894__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput390 _0767_/X vssd1 vssd1 vccd1 vccd1 cap_addr[8] sky130_fd_sc_hd__buf_12
XFILLER_0_233_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_362_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_370_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0710_ _0710_/A1 _0505_/Y _0518_/B _0710_/B2 vssd1 vssd1 vccd1 vccd1 _0713_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_154_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output388_A _0763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold509 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0641_ _0641_/A _0641_/B _0641_/C vssd1 vssd1 vccd1 vccd1 _0641_/X sky130_fd_sc_hd__or3_4
XANTENNA_output555_A hold269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0572_ input31/X _0598_/A2 _0586_/B1 input67/X vssd1 vssd1 vccd1 vccd1 _0572_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_291_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1124_ _1188_/CLK _1124_/D vssd1 vssd1 vccd1 vccd1 _1124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1055_ _1053_/X _1057_/B _0956_/Y vssd1 vssd1 vccd1 vccd1 _1055_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_393_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0908_ hold197/X _0953_/A2 _0907_/X vssd1 vssd1 vccd1 vccd1 _0908_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_302_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0839_ _1080_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0839_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput118 io_oeb_z80[35] vssd1 vssd1 vccd1 vccd1 _0605_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput107 io_oeb_z80[25] vssd1 vssd1 vccd1 vccd1 _0581_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_215_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput129 io_out_6502[12] vssd1 vssd1 vccd1 vccd1 _0655_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_270_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold331_A _1093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_80 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_91 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_375_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_316_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_316_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold306 _1101_/Q vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _0881_/X vssd1 vssd1 vccd1 vccd1 _1130_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0624_ _0624_/A1 _0660_/A2 _0628_/B1 _0624_/B2 vssd1 vssd1 vccd1 vccd1 _0625_/C sky130_fd_sc_hd__a22o_2
XANTENNA__0502__A hold99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold328 hold704/X vssd1 vssd1 vccd1 vccd1 _1181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 hold674/X vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0555_ input24/X _0604_/A2 _0586_/B1 input60/X vssd1 vssd1 vccd1 vccd1 _0555_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_252_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1107_ _1214_/CLK _1107_/D vssd1 vssd1 vccd1 vccd1 _1107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_366_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1038_ _1038_/A _1038_/B vssd1 vssd1 vccd1 vccd1 _1038_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_366_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_381_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_366_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1243__A _1243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_382_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0798__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_313_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_276_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output420_A _1094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0946__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold653/X vssd1 vssd1 vccd1 vccd1 _0821_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _0955_/X vssd1 vssd1 vccd1 vccd1 _1155_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold136 hold534/X vssd1 vssd1 vccd1 vccd1 _1182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _1213_/Q vssd1 vssd1 vccd1 vccd1 _0823_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold598/X vssd1 vssd1 vccd1 vccd1 _1171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0607_ _0607_/A1 _0747_/A2 _0516_/B _0607_/B2 vssd1 vssd1 vccd1 vccd1 _0609_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_229_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout605 hold100/X vssd1 vssd1 vccd1 vccd1 _0598_/A2 sky130_fd_sc_hd__buf_4
Xhold169 _0827_/X vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0538_ input51/X _0598_/A2 _0598_/B1 input87/X vssd1 vssd1 vccd1 vccd1 _0538_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout616 _0500_/Y vssd1 vssd1 vccd1 vccd1 _0966_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1238__A _1238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0937__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold681 _1201_/Q vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold670 _1202_/Q vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _0873_/X vssd1 vssd1 vccd1 vccd1 _0874_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_246_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_389_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0640__B2 _0640_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output468_A _0677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput290 io_out_vliw[28] vssd1 vssd1 vccd1 vccd1 _0720_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_368_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0631__B2 _0631_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0631__A1 _0631_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_304_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0934__A2 _0775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0897__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0698__B2 _0698_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_359_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0622__B2 _0622_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_388_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ hold203/X _0953_/A2 _0940_/X vssd1 vssd1 vccd1 vccd1 _0941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0872_ hold76/X _1082_/C vssd1 vssd1 vccd1 vccd1 _0872_/X sky130_fd_sc_hd__or2_1
XFILLER_0_341_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_301_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1157_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_386_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0510__A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_333_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1060__B _1181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_364_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0604__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput561 hold188/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput550 hold222/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_12
Xoutput572 hold262/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_245_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_359_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1251__A _1251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_390_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_382_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_251_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1140_ _1175_/CLK _1140_/D vssd1 vssd1 vccd1 vccd1 _1140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_358_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1071_ _1071_/A _1071_/B _1072_/A _1071_/D vssd1 vssd1 vccd1 vccd1 _1078_/B sky130_fd_sc_hd__and4_1
XFILLER_0_393_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_181 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0924_ _1036_/A _0924_/B vssd1 vssd1 vccd1 vccd1 _0924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0855_ hold252/X hold729/A hold661/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0855_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0786_ hold333/X _0840_/A2 _0785_/X _0500_/Y vssd1 vssd1 vccd1 vccd1 _0786_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1246__A _1246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput391 _1087_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[0] sky130_fd_sc_hd__buf_12
XFILLER_0_233_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_254_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0640_ _0640_/A1 _0660_/A2 _0696_/B1 _0640_/B2 vssd1 vssd1 vccd1 vccd1 _0641_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_256_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0571_ _0571_/A1 _0506_/B _0569_/A _0570_/X vssd1 vssd1 vccd1 vccd1 _1251_/A sky130_fd_sc_hd__a211o_4
XANTENNA_output548_A hold197/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output450_A _0601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0752__A0 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_378_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1123_ _1157_/CLK _1123_/D vssd1 vssd1 vccd1 vccd1 _1123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1054_ _1060_/A _1060_/D vssd1 vssd1 vccd1 vccd1 _1054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0907_ hold308/X _0952_/A2 _0952_/B1 _1024_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0907_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0838_ hold529/X _0840_/A2 hold164/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0838_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_101_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0769_ _0955_/A hold695/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_339_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0743__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput108 io_oeb_z80[26] vssd1 vssd1 vccd1 vccd1 _0583_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_270_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput119 io_oeb_z80[3] vssd1 vssd1 vccd1 vccd1 _0531_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout579_A _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_304_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_81 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_92 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_70 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0799__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0734__B1 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_375_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_331_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold307 hold667/X vssd1 vssd1 vccd1 vccd1 _1101_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0623_ _0623_/A1 _0514_/B _0695_/B1 _0623_/B2 vssd1 vssd1 vccd1 vccd1 _0625_/B sky130_fd_sc_hd__a22o_1
Xhold318 _1113_/Q vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _1102_/Q vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_256_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0554_ input95/X _0590_/A2 _0565_/A _0553_/X vssd1 vssd1 vccd1 vccd1 _1245_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_110_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_252_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_252_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1106_ _1214_/CLK _1106_/D vssd1 vssd1 vccd1 vccd1 _1106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1037_ _1038_/A _1037_/B _1037_/C _1037_/D vssd1 vssd1 vccd1 vccd1 _1050_/D sky130_fd_sc_hd__and4_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput90 io_oeb_z80[0] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_293_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0707__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0513__A _0860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold104 hold86/X vssd1 vssd1 vccd1 vccd1 _0860_/A sky130_fd_sc_hd__buf_2
Xhold115 hold341/X vssd1 vssd1 vccd1 vccd1 hold342/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold594/X vssd1 vssd1 vccd1 vccd1 _1178_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 hold581/X vssd1 vssd1 vccd1 vccd1 _1179_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold707/X vssd1 vssd1 vccd1 vccd1 _0819_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 hold677/X vssd1 vssd1 vccd1 vccd1 _0809_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0606_ _0606_/A1 _0746_/A2 _0746_/B1 _0606_/B2 vssd1 vssd1 vccd1 vccd1 _0609_/A sky130_fd_sc_hd__a22o_1
Xfanout606 hold100/X vssd1 vssd1 vccd1 vccd1 _0604_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0537_ _0537_/A1 _0506_/B _0529_/X _0536_/X vssd1 vssd1 vccd1 vccd1 _1237_/A sky130_fd_sc_hd__a211o_4
Xfanout617 _0500_/Y vssd1 vssd1 vccd1 vccd1 _0955_/B sky130_fd_sc_hd__buf_4
XFILLER_0_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout611_A _0851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold660 _0853_/X vssd1 vssd1 vccd1 vccd1 _0854_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _0802_/X vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold693 _0874_/X vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _0800_/X vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1254__A _1254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_389_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_266_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput280 io_out_vliw[19] vssd1 vssd1 vccd1 vccd1 _0684_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_306_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput291 io_out_vliw[29] vssd1 vssd1 vccd1 vccd1 _0724_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_236_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0508__A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0631__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1224__D hold4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_363_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0855__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_327_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1249__A _1249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_295_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold490 hold490/A vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_263_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_271_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0587__C_N hold99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_377_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0846__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_385_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ hold521/X _0952_/A2 _0952_/B1 _1071_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0940_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0871_ hold301/X hold729/A hold652/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0871_/X sky130_fd_sc_hd__o211a_1
XANTENNA_output480_A _0613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0510__B _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_379_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_364_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1014__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput562 hold217/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_12
Xoutput551 hold209/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_12
Xoutput540 hold412/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_12
XFILLER_0_285_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_295_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0531__A1 _0531_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1070_ _0833_/A _1076_/B hold555/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1070_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0834__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_160 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_182 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0598__A1 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0923_ hold176/X _0953_/A2 _0922_/X vssd1 vssd1 vccd1 vccd1 _0923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_302_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0854_ _0880_/A _0854_/B vssd1 vssd1 vccd1 vccd1 _0854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_259_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0785_ _0847_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0785_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_328_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_282_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0522__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1199_ _1204_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 _1199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold102_A _0601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1002__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput392 _1097_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[10] sky130_fd_sc_hd__buf_12
XFILLER_0_254_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1262__A hold96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0816__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_370_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0570_ input30/X _0598_/A2 _0586_/B1 input66/X vssd1 vssd1 vccd1 vccd1 _0570_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_122_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output443_A _1258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1122_ _1175_/CLK _1122_/D vssd1 vssd1 vccd1 vccd1 _1122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1053_ _1060_/A _1060_/D vssd1 vssd1 vccd1 vccd1 _1053_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_346_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0516__A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0906_ _1085_/A _0906_/B vssd1 vssd1 vccd1 vccd1 _0906_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0837_ _1076_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__or2_1
XFILLER_0_302_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0768_ _0768_/A _0768_/B vssd1 vssd1 vccd1 vccd1 _0771_/B sky130_fd_sc_hd__and2_1
XANTENNA__0743__A1 _0743_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0743__B2 _0743_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput109 io_oeb_z80[27] vssd1 vssd1 vccd1 vccd1 _0585_/A1 sky130_fd_sc_hd__clkbuf_2
X_0699_ _0699_/A1 _0747_/A2 _0515_/Y _0699_/B2 vssd1 vssd1 vccd1 vccd1 _0701_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_371_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_60 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_93 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_71 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1257__A _1257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_249_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0734__B2 _0734_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output393_A _1098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output560_A hold203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold308 _1103_/Q vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_296_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0622_ _0622_/A1 _0674_/A2 _0674_/B1 _0622_/B2 vssd1 vssd1 vccd1 vccd1 _0625_/A sky130_fd_sc_hd__a22o_1
Xhold319 hold710/X vssd1 vssd1 vccd1 vccd1 _1113_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0553_ input23/X _0604_/A2 _0586_/B1 input59/X vssd1 vssd1 vccd1 vccd1 _0553_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_249_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_264_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1105_ _1214_/CLK _1105_/D vssd1 vssd1 vccd1 vccd1 _1105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1036_ _1036_/A _1036_/B vssd1 vssd1 vccd1 vccd1 _1036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_381_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_334_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput91 io_oeb_z80[10] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_2
Xinput80 io_oeb_vliw[33] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0716__B2 _0716_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_A _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_306_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0707__A1 _0707_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0707__B2 _0707_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0643__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_371_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold105 _0505_/Y vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__buf_1
Xhold116 hold343/X vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__buf_1
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold149 hold611/X vssd1 vssd1 vccd1 vccd1 _1177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold573/X vssd1 vssd1 vccd1 vccd1 _1172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold687/X vssd1 vssd1 vccd1 vccd1 _0793_/A sky130_fd_sc_hd__dlygate4sd3_1
X_0605_ _0605_/A1 _0605_/A2 _0593_/X _0604_/X vssd1 vssd1 vccd1 vccd1 _1266_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout607 _0508_/B vssd1 vssd1 vccd1 vccd1 _0732_/A2 sky130_fd_sc_hd__buf_4
X_0536_ input50/X _0598_/A2 _0598_/B1 input86/X vssd1 vssd1 vccd1 vccd1 _0536_/X sky130_fd_sc_hd__a22o_1
Xfanout618 _0500_/Y vssd1 vssd1 vccd1 vccd1 _1081_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_336_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1019_ _0807_/A _1021_/A hold597/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _1019_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_394_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_307_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout604_A hold82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 _1091_/Q vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _0854_/X vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _1205_/Q vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_275_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _1199_/Q vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_353_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput281 io_out_vliw[1] vssd1 vssd1 vccd1 vccd1 _0612_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput270 io_out_vliw[0] vssd1 vssd1 vccd1 vccd1 _0608_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_368_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput292 io_out_vliw[2] vssd1 vssd1 vccd1 vccd1 _0616_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_395_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_289_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0519_ hold99/A hold86/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__nand2_1
XFILLER_0_213_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_382_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0607__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_382_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1265__A _1265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 hold35/X vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_263_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_263_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_310_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0870_ _0880_/A _0870_/B vssd1 vssd1 vccd1 vccd1 _0870_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output473_A _0693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0782__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0519__A hold99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_368_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_364_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_364_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0999_ _0999_/A _1165_/Q _1166_/Q _0999_/D vssd1 vssd1 vccd1 vccd1 _1017_/C sky130_fd_sc_hd__and4_1
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput530 _1235_/X vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__1085__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput552 hold220/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput563 hold297/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_12
Xoutput541 hold252/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_0_285_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_245_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmultiplexer_621 vssd1 vssd1 vccd1 vccd1 multiplexer_621/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_0_374_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_295_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0531__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_161 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_150 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_172 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 hold37/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0922_ hold276/X _0952_/A2 _0952_/B1 _1050_/A _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0922_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_314_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0853_ hold346/X _0776_/A hold604/X _0967_/A _0852_/X vssd1 vssd1 vccd1 vccd1 _0853_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_140_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0784_ hold339/X _0810_/A2 _0783_/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0784_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_87_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_391_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput1 cap_io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_0_344_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0522__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1267_ _1267_/A vssd1 vssd1 vccd1 vccd1 _1267_/X sky130_fd_sc_hd__buf_1
XFILLER_0_356_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1198_ _1224_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 _1198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_349_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_364_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_258_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput393 _1098_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[11] sky130_fd_sc_hd__buf_12
Xoutput382 _0751_/X vssd1 vssd1 vccd1 vccd1 cap_addr[0] sky130_fd_sc_hd__buf_12
XFILLER_0_273_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_318_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_343_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_370_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output436_A _1251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1121_ _1175_/CLK _1121_/D vssd1 vssd1 vccd1 vccd1 _1121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1052_ _0823_/A _1080_/B hold580/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1052_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0516__B _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0905_ hold191/X _0880_/A _0904_/X vssd1 vssd1 vccd1 vccd1 _0905_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_259_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0836_ hold523/X _0840_/A2 hold246/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0836_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0767_ _0767_/A _0767_/B _0767_/C vssd1 vssd1 vccd1 vccd1 _0767_/X sky130_fd_sc_hd__and3_4
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_302_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0698_ _0698_/A1 _0746_/A2 _0746_/B1 _0698_/B2 vssd1 vssd1 vccd1 vccd1 _0701_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_282_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_325_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_50 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold212_A _1094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_72 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_94 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_246_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0670__B2 _0670_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_343_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output386_A _0759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0621_ _0621_/A _0621_/B _0621_/C vssd1 vssd1 vccd1 vccd1 _0621_/X sky130_fd_sc_hd__or3_4
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output553_A hold232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 hold678/X vssd1 vssd1 vccd1 vccd1 _1103_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0973__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0552_ input94/X _0605_/A2 _0565_/A _0551_/X vssd1 vssd1 vccd1 vccd1 _1244_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_249_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_264_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1104_ _1180_/CLK _1104_/D vssd1 vssd1 vccd1 vccd1 _1104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1035_ _0815_/A _0956_/Y _1034_/X vssd1 vssd1 vccd1 vccd1 _1035_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_322_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0949__C1 _0952_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput81 io_oeb_vliw[34] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_1
Xinput70 io_oeb_vliw[24] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
X_0819_ _0819_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0819_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput92 io_oeb_z80[11] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_228_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_270_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_270_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_315_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_357_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0652__B2 _0652_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0900__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0643__A1 _0643_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0643__B2 _0643_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_371_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_304_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold106 hold160/X vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold117 hold683/X vssd1 vssd1 vccd1 vccd1 _0795_/A sky130_fd_sc_hd__dlygate4sd3_1
X_0604_ input46/X _0604_/A2 _0510_/B input82/X vssd1 vssd1 vccd1 vccd1 _0604_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold128 hold615/X vssd1 vssd1 vccd1 vccd1 hold616/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold681/X vssd1 vssd1 vccd1 vccd1 _0799_/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout608 _0660_/A2 vssd1 vssd1 vccd1 vccd1 _0508_/B sky130_fd_sc_hd__buf_2
X_0535_ _0535_/A1 _0506_/B _0529_/X _0534_/X vssd1 vssd1 vccd1 vccd1 _1236_/A sky130_fd_sc_hd__a211o_4
Xfanout619 _1085_/A vssd1 vssd1 vccd1 vccd1 _1036_/A sky130_fd_sc_hd__buf_4
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_252_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1018_ hold596/X _1037_/B _1021_/A vssd1 vssd1 vccd1 vccd1 _1018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_347_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0634__B2 _0634_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_362_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold651 _0869_/X vssd1 vssd1 vccd1 vccd1 _0870_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _1200_/Q vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 _0971_/Y vssd1 vssd1 vccd1 vccd1 _0972_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold673 _0808_/X vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _0771_/B vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _0796_/X vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_353_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0561__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput271 io_out_vliw[10] vssd1 vssd1 vccd1 vccd1 _0648_/B2 sky130_fd_sc_hd__buf_2
Xinput260 io_out_scrapcpu[33] vssd1 vssd1 vccd1 vccd1 _0740_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_269_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output516_A _1258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput293 io_out_vliw[30] vssd1 vssd1 vccd1 vccd1 _0728_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput282 io_out_vliw[20] vssd1 vssd1 vccd1 vccd1 _0688_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_376_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0616__B2 _0616_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0518_ _0518_/A _0518_/B vssd1 vssd1 vccd1 vccd1 _0518_/X sky130_fd_sc_hd__and2_2
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_379_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0855__A1 hold252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_394_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_382_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0607__A1 _0607_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_312_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_312_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_350_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold470 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold481 hold481/A vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_263_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold492 hold51/X vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0846__A1 hold99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output466_A _0669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_364_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_289_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0998_ _1166_/Q _0995_/B _0999_/D vssd1 vssd1 vccd1 vccd1 _0998_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_332_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput520 _1261_/X vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_12
XFILLER_0_131_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0701__C _0701_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput531 _1236_/X vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_12
Xoutput553 hold232/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput542 hold291/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_12
XFILLER_0_300_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput564 hold229/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0525__B1 hold95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmultiplexer_622 vssd1 vssd1 vccd1 vccd1 multiplexer_622/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_0_213_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0764__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_151 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_140 hold477/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_173 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_162 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 hold63/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_361_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0921_ _1036_/A _0921_/B vssd1 vssd1 vccd1 vccd1 _0921_/Y sky130_fd_sc_hd__nor2_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0852_ _0852_/A _1082_/C vssd1 vssd1 vccd1 vccd1 _0852_/X sky130_fd_sc_hd__or2_1
XFILLER_0_314_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0783_ _0845_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0783_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_384_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 cap_io_in[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
XFILLER_0_369_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1266_ _1266_/A vssd1 vssd1 vccd1 vccd1 _1266_/X sky130_fd_sc_hd__buf_1
XFILLER_0_250_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1197_ _1224_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 _1197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_364_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput394 _1099_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[12] sky130_fd_sc_hd__buf_12
Xoutput383 _0753_/X vssd1 vssd1 vccd1 vccd1 cap_addr[1] sky130_fd_sc_hd__buf_12
XFILLER_0_387_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1188_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_395_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_270_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0903__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0985__B1 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_295_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1120_ _1188_/CLK _1120_/D vssd1 vssd1 vccd1 vccd1 _1120_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output429_A _1245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1051_ hold579/X _1060_/D _1076_/B vssd1 vssd1 vccd1 vccd1 _1051_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0904_ hold329/X _0776_/A hold605/A _1016_/D _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0904_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0835_ _1073_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0835_/X sky130_fd_sc_hd__or2_1
XANTENNA__0976__B1 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_339_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0766_ input9/X _1095_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0767_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0697_ _0697_/A _0697_/B _0697_/C vssd1 vssd1 vccd1 vccd1 _0697_/X sky130_fd_sc_hd__or3_4
XFILLER_0_121_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_282_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1082__C _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1249_ _1249_/A vssd1 vssd1 vccd1 vccd1 _1249_/X sky130_fd_sc_hd__buf_1
XFILLER_0_369_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_40 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_84 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_95 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0719__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_265_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0620_ _0620_/A1 _0660_/A2 _0628_/B1 _0620_/B2 vssd1 vssd1 vccd1 vccd1 _0621_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_296_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0551_ input22/X _0604_/A2 _0598_/B1 input58/X vssd1 vssd1 vccd1 vccd1 _0551_/X sky130_fd_sc_hd__a22o_1
XANTENNA_output546_A hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_264_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1103_ _1180_/CLK _1103_/D vssd1 vssd1 vccd1 vccd1 _1103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1034_ _1032_/B _1028_/X _1038_/B _1080_/B vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_220_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput82 io_oeb_vliw[35] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
Xinput71 io_oeb_vliw[25] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput60 io_oeb_vliw[15] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_1
X_0818_ hold289/X _0840_/A2 _0817_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0818_/X sky130_fd_sc_hd__o211a_1
Xhold800 _1136_/Q vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput93 io_oeb_z80[12] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_366_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0749_ _0749_/A _0749_/B _0749_/C vssd1 vssd1 vccd1 vccd1 _0749_/X sky130_fd_sc_hd__or3_4
XFILLER_0_228_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout577_A _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_251_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_325_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_321_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_388_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0643__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 hold162/X vssd1 vssd1 vccd1 vccd1 _0868_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0603_ _0603_/A1 _0605_/A2 _0593_/X _0602_/X vssd1 vssd1 vccd1 vccd1 _1265_/A sky130_fd_sc_hd__a211o_4
Xhold118 hold631/X vssd1 vssd1 vccd1 vccd1 hold632/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold668/X vssd1 vssd1 vccd1 vccd1 _0803_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout609 _0507_/X vssd1 vssd1 vccd1 vccd1 _0660_/A2 sky130_fd_sc_hd__clkbuf_4
X_0534_ input49/X _0598_/A2 _0598_/B1 input85/X vssd1 vssd1 vccd1 vccd1 _0534_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0867__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_339_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1017_ _1017_/A _1017_/B _1017_/C _1017_/D vssd1 vssd1 vccd1 vccd1 _1037_/B sky130_fd_sc_hd__and4_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_303_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 _0993_/Y vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_377_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold652 _0870_/X vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _0798_/X vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _0973_/X vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 _1217_/Q vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _1090_/Q vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _1196_/Q vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_283_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0570__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_393_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0561__A1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput272 io_out_vliw[11] vssd1 vssd1 vccd1 vccd1 _0652_/B2 sky130_fd_sc_hd__buf_2
Xinput261 io_out_scrapcpu[34] vssd1 vssd1 vccd1 vccd1 _0744_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput250 io_out_scrapcpu[24] vssd1 vssd1 vccd1 vccd1 _0704_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput294 io_out_vliw[31] vssd1 vssd1 vccd1 vccd1 _0732_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput283 io_out_vliw[21] vssd1 vssd1 vccd1 vccd1 _0692_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_234_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_376_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0805__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0517_ hold99/X _0517_/B hold93/X vssd1 vssd1 vccd1 vccd1 _0526_/A sky130_fd_sc_hd__and3_4
XFILLER_0_265_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0552__A1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold471 hold41/X vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 hold460/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold482 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 hold493/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0543__A1 _0543_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0906__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_381_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output459_A _0641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_393_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_376_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_263_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold96_A hold96/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_332_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0997_ _0797_/A _0996_/A hold624/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0997_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_332_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput510 _1252_/X vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_12
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput521 hold97/X vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_12
Xoutput532 _1237_/X vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_12
Xoutput554 hold176/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput543 hold303/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput565 hold257/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_12
XFILLER_0_374_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0525__A1 _0525_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_307_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_253_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmultiplexer_623 vssd1 vssd1 vccd1 vccd1 multiplexer_623/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XFILLER_0_213_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0828__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0764__A1 _1094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold771_A _1096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_291_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold290 hold714/X vssd1 vssd1 vccd1 vccd1 _1107_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_244_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_130 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_152 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_141 hold498/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_174 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_373_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_163 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ hold232/X _0953_/A2 _0919_/X vssd1 vssd1 vccd1 vccd1 _0920_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0851_ _0851_/A _0851_/B _0841_/B vssd1 vssd1 vccd1 vccd1 _0851_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_314_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0782_ hold337/X _0810_/A2 _0781_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0782_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_377_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1265_ _1265_/A vssd1 vssd1 vccd1 vccd1 _1265_/X sky130_fd_sc_hd__buf_1
Xinput3 cap_io_in[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
XFILLER_0_344_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1196_ _1224_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 _1196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0691__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_364_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_369_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0746__A1 _0746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0746__B2 _0746_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput395 _1100_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[13] sky130_fd_sc_hd__buf_12
Xoutput384 _0755_/X vssd1 vssd1 vccd1 vccd1 cap_addr[2] sky130_fd_sc_hd__buf_12
XFILLER_0_318_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_343_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1050_ _1050_/A _1050_/B _1050_/C _1050_/D vssd1 vssd1 vccd1 vccd1 _1060_/D sky130_fd_sc_hd__and4_2
XFILLER_0_393_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0813__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0903_ _1085_/A _0903_/B vssd1 vssd1 vccd1 vccd1 _0903_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0834_ hold278/X _0840_/A2 _0833_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0834_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_153_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0728__B2 _0728_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0765_ _0767_/A _0767_/B _0765_/C vssd1 vssd1 vccd1 vccd1 _0765_/X sky130_fd_sc_hd__and3_4
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0696_ _0696_/A1 _0732_/A2 _0696_/B1 _0696_/B2 vssd1 vssd1 vccd1 vccd1 _0697_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_269_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_369_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1248_ _1248_/A vssd1 vssd1 vccd1 vccd1 _1248_/X sky130_fd_sc_hd__buf_1
XFILLER_0_371_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1179_ _1184_/CLK _1179_/D vssd1 vssd1 vccd1 vccd1 _1179_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_41 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_52 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold100_A _0507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_320_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0719__A1 _0719_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0719__B2 _0719_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_265_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0655__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0617__C _0617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0550_ input93/X _0605_/A2 _0565_/A _0549_/X vssd1 vssd1 vccd1 vccd1 _1243_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output441_A _1256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1102_ _1188_/CLK _1102_/D vssd1 vssd1 vccd1 vccd1 _1102_/Q sky130_fd_sc_hd__dfxtp_1
X_1033_ _1033_/A _1037_/D vssd1 vssd1 vccd1 vccd1 _1038_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_319_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0646__B1 _0526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_322_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 io_oeb_scrapcpu[6] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xinput72 io_oeb_vliw[26] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
Xinput61 io_oeb_vliw[16] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_1
X_0817_ _0817_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0817_/X sky130_fd_sc_hd__or2_1
Xhold801 _1135_/Q vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
X_0748_ _0748_/A1 _0508_/B _0748_/B1 _0748_/B2 vssd1 vssd1 vccd1 vccd1 _0749_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_287_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput94 io_oeb_z80[13] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_2
Xinput83 io_oeb_vliw[3] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_1
XFILLER_0_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0679_ _0679_/A1 _0747_/A2 _0683_/B1 _0679_/B2 vssd1 vssd1 vccd1 vccd1 _0681_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_228_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_304_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output489_A _1181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold108 _0512_/X vssd1 vssd1 vccd1 vccd1 _0515_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0602_ input45/X _0604_/A2 _0510_/B input81/X vssd1 vssd1 vccd1 vccd1 _0602_/X sky130_fd_sc_hd__a22o_1
Xhold119 hold679/X vssd1 vssd1 vccd1 vccd1 _0791_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0533_ _0533_/A1 _0506_/B _0529_/X _0532_/X vssd1 vssd1 vccd1 vccd1 _1235_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0619__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1016_ _1168_/Q _1016_/B _1016_/C _1016_/D vssd1 vssd1 vccd1 vccd1 _1017_/D sky130_fd_sc_hd__and4_1
XFILLER_0_354_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold620 _1006_/X vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_275_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold653 _1212_/Q vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 _1157_/Q vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold631 _0994_/X vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_275_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold697 _1066_/X vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _1089_/Q vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _0784_/X vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _0790_/X vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_283_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold265_A _1095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_326_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_367_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput262 io_out_scrapcpu[35] vssd1 vssd1 vccd1 vccd1 _0748_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput251 io_out_scrapcpu[25] vssd1 vssd1 vccd1 vccd1 _0708_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput240 io_out_scrapcpu[15] vssd1 vssd1 vccd1 vccd1 _0668_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput295 io_out_vliw[32] vssd1 vssd1 vccd1 vccd1 _0736_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput284 io_out_vliw[22] vssd1 vssd1 vccd1 vccd1 _0696_/B2 sky130_fd_sc_hd__buf_2
Xinput273 io_out_vliw[12] vssd1 vssd1 vccd1 vccd1 _0656_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_236_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_376_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_344_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0821__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_257_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_300_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0516_ _0518_/A _0516_/B vssd1 vssd1 vccd1 vccd1 _0516_/X sky130_fd_sc_hd__and2_2
XFILLER_0_277_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_379_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_394_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_257_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold450 hold25/X vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold483 hold47/X vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0625__C _0625_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_239_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0782__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_294_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold89_A hold89/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_332_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0996_ _0996_/A _0996_/B vssd1 vssd1 vccd1 vccd1 _0996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput511 _1253_/X vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_12
Xoutput500 _1243_/X vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_12
XFILLER_0_300_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput522 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__buf_6
Xoutput533 _1238_/X vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_12
Xoutput544 hold254/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput555 hold269/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput566 hold250/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_300_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0525__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_374_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmultiplexer_624 vssd1 vssd1 vccd1 vccd1 io_oeb[0] multiplexer_624/LO sky130_fd_sc_hd__conb_1
XFILLER_0_213_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_370_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold280 hold399/X vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_348_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold291 hold397/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_131 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_120 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_142 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_175 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_153 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_164 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_361_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_314_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0850_ hold116/X hold739/X hold356/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0850_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output569_A hold310/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0781_ _0965_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0781_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output471_A _0685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1264_ _1264_/A vssd1 vssd1 vccd1 vccd1 _1264_/X sky130_fd_sc_hd__buf_1
Xinput4 cap_io_in[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_0_344_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_250_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1195_ _1204_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _1195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_360_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0691__B2 _0691_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0691__A1 _0691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_364_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0994__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0979_ _0983_/C _0979_/B vssd1 vssd1 vccd1 vccd1 _0979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput396 _1101_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[14] sky130_fd_sc_hd__buf_12
Xoutput385 _0757_/X vssd1 vssd1 vccd1 vccd1 cap_addr[3] sky130_fd_sc_hd__buf_12
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_318_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_387_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0682__B2 _0682_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout590 _0526_/A vssd1 vssd1 vccd1 vccd1 _0674_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_164_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_334_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0902_ hold237/X _0880_/A _0901_/X vssd1 vssd1 vccd1 vccd1 _0902_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0833_ _0833_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0833_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0764_ input8/X _1094_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0765_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0695_ _0695_/A1 _0747_/A2 _0695_/B1 _0695_/B2 vssd1 vssd1 vccd1 vccd1 _0697_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_369_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1247_ _1247_/A vssd1 vssd1 vccd1 vccd1 _1247_/X sky130_fd_sc_hd__buf_1
XFILLER_0_2_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1178_ _1221_/CLK _1178_/D vssd1 vssd1 vccd1 vccd1 _1178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_377_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0664__B2 _0664_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_392_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_304_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_53 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_42 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_86 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0719__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0655__A1 _0655_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0655__B2 _0655_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_383_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_316_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0633__C _0633_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0591__B1 hold95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output434_A _1249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1101_ _1205_/CLK _1101_/D vssd1 vssd1 vccd1 vccd1 _1101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_260_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1032_ _1032_/A _1032_/B vssd1 vssd1 vccd1 vccd1 _1037_/D sky130_fd_sc_hd__and2_1
XFILLER_0_359_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0646__B2 _0646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_374_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput40 io_oeb_scrapcpu[2] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_330_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput51 io_oeb_scrapcpu[7] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput73 io_oeb_vliw[27] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
Xinput62 io_oeb_vliw[17] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_1
Xhold802 _1143_/Q vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
X_0816_ hold320/X _0840_/A2 _0815_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0816_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_330_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0747_ _0747_/A1 _0747_/A2 _0516_/B _0747_/B2 vssd1 vssd1 vccd1 vccd1 _0749_/B sky130_fd_sc_hd__a22o_1
Xinput95 io_oeb_z80[14] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_2
Xinput84 io_oeb_vliw[4] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0678_ _0678_/A1 _0746_/A2 _0746_/B1 _0678_/B2 vssd1 vssd1 vccd1 vccd1 _0681_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_380_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_380_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold308_A _1103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_333_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_246_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_246_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_388_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0628__B2 _0628_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output384_A _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0601_ _0601_/A1 _0605_/A2 hold95/X hold101/X vssd1 vssd1 vccd1 vccd1 _0601_/X sky130_fd_sc_hd__a211o_4
Xhold109 _0592_/X vssd1 vssd1 vccd1 vccd1 _1260_/A sky130_fd_sc_hd__buf_1
X_0532_ input48/X _0598_/A2 _0598_/B1 input84/X vssd1 vssd1 vccd1 vccd1 _0532_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0564__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0819__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0867__A1 hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0619__B2 _0619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0619__A1 _0619_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1015_ _1016_/D _1015_/B vssd1 vssd1 vccd1 vccd1 _1015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_362_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold610 _1043_/Y vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold621 hold621/A vssd1 vssd1 vccd1 vccd1 _1168_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_330_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold654 _0822_/X vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 _0961_/B vssd1 vssd1 vccd1 vccd1 _0967_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 hold632/A vssd1 vssd1 vccd1 vccd1 _1165_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold665 _0782_/X vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 _1088_/Q vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 _1198_/Q vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_290_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold698 _1219_/Q vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_243_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput230 io_out_as1802[6] vssd1 vssd1 vccd1 vccd1 _0631_/B2 sky130_fd_sc_hd__buf_2
Xinput252 io_out_scrapcpu[26] vssd1 vssd1 vccd1 vccd1 _0712_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput241 io_out_scrapcpu[16] vssd1 vssd1 vccd1 vccd1 _0672_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput263 io_out_scrapcpu[3] vssd1 vssd1 vccd1 vccd1 _0620_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput296 io_out_vliw[33] vssd1 vssd1 vccd1 vccd1 _0740_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput285 io_out_vliw[23] vssd1 vssd1 vccd1 vccd1 _0700_/B2 sky130_fd_sc_hd__buf_2
Xinput274 io_out_vliw[13] vssd1 vssd1 vccd1 vccd1 _0660_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_383_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_388_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_252_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_312_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0515_ _0517_/B _0515_/B vssd1 vssd1 vccd1 vccd1 _0515_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_265_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_367_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold462 hold33/X vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 hold451/A vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold484 hold484/A vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold55/X vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0641__C _0641_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_239_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_294_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output514_A _1256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_376_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0995_ _0995_/A _0995_/B vssd1 vssd1 vccd1 vccd1 _0995_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__0758__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput501 _1244_/X vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_12
XFILLER_0_300_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput523 _1264_/X vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_12
Xoutput512 _1254_/X vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_12
Xoutput545 hold240/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput534 _0514_/X vssd1 vssd1 vccd1 vccd1 rst_6502 sky130_fd_sc_hd__buf_12
XFILLER_0_300_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput556 hold173/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput567 hold301/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_285_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmultiplexer_625 vssd1 vssd1 vccd1 vccd1 la_data_out[0] multiplexer_625/LO sky130_fd_sc_hd__conb_1
XFILLER_0_390_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_308_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_276_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_268_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_276_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold270 _0926_/Y vssd1 vssd1 vccd1 vccd1 _0927_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold292 _0890_/Y vssd1 vssd1 vccd1 vccd1 _0891_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _0884_/Y vssd1 vssd1 vccd1 vccd1 _0885_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_132 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_110 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_121 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_143 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_176 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_373_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_165 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_154 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0780_ hold335/X _0810_/A2 _0779_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0780_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output464_A _0661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1263_ hold89/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__clkbuf_1
Xinput5 cap_io_in[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1194_ _1204_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 _1194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_337_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_369_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0978_ _0983_/C _0979_/B vssd1 vssd1 vccd1 vccd1 _0978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput386 _0759_/X vssd1 vssd1 vccd1 vccd1 cap_addr[4] sky130_fd_sc_hd__buf_12
XFILLER_0_273_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput397 _1102_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[15] sky130_fd_sc_hd__buf_12
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_387_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0753__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_311_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_276_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_272_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout591 _0518_/B vssd1 vssd1 vccd1 vccd1 _0746_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout580 _0775_/Y vssd1 vssd1 vccd1 vccd1 _0810_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_232_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_260_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0901_ hold306/X _0776_/A hold605/A _1016_/C _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0901_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1083__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0832_ hold521/X _0840_/A2 hold195/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0832_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0763_ _0767_/A _0767_/B _0763_/C vssd1 vssd1 vccd1 vccd1 _0763_/X sky130_fd_sc_hd__and3_4
XFILLER_0_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0694_ _0694_/A1 _0746_/A2 _0746_/B1 _0694_/B2 vssd1 vssd1 vccd1 vccd1 _0697_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1246_ _1246_/A vssd1 vssd1 vccd1 vccd1 _1246_/X sky130_fd_sc_hd__buf_1
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1177_ _1214_/CLK _1177_/D vssd1 vssd1 vccd1 vccd1 _1177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_10 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_87 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_98 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0655__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_324_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_245_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1100_ _1205_/CLK _1100_/D vssd1 vssd1 vccd1 vccd1 _1100_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_output427_A _1243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1031_ _0813_/A _1080_/B hold576/X _0955_/B vssd1 vssd1 vccd1 vccd1 _1031_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0646__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput30 io_oeb_scrapcpu[20] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput41 io_oeb_scrapcpu[30] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
XFILLER_0_287_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput52 io_oeb_scrapcpu[8] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput63 io_oeb_vliw[18] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_1
XFILLER_0_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0815_ _0815_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0815_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0746_ _0746_/A1 _0746_/A2 _0746_/B1 _0746_/B2 vssd1 vssd1 vccd1 vccd1 _0749_/A sky130_fd_sc_hd__a22o_1
Xinput96 io_oeb_z80[15] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
Xinput74 io_oeb_vliw[28] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_1
Xinput85 io_oeb_vliw[5] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1225_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_366_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0677_ _0677_/A _0677_/B _0677_/C vssd1 vssd1 vccd1 vccd1 _0677_/X sky130_fd_sc_hd__or3_4
XFILLER_0_149_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_255_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_380_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0573__A1 _0573_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_261_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_388_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_372_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0800__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0600_ input44/X _0604_/A2 _0510_/B input80/X vssd1 vssd1 vccd1 vccd1 _0600_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0531_ _0531_/A1 _0506_/B _0529_/X _0530_/X vssd1 vssd1 vccd1 vccd1 _1234_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0564__A1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output544_A hold254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0619__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0835__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1014_ _0805_/A _1021_/A hold584/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_362_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold611 _1044_/X vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold600 hold600/A vssd1 vssd1 vccd1 vccd1 _0967_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold644 _0857_/X vssd1 vssd1 vccd1 vccd1 _0858_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 hold642/X vssd1 vssd1 vccd1 vccd1 _0961_/B sky130_fd_sc_hd__buf_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold622 hold774/X vssd1 vssd1 vccd1 vccd1 _0995_/A sky130_fd_sc_hd__buf_1
X_0729_ _0729_/A _0729_/B _0729_/C vssd1 vssd1 vccd1 vccd1 _0729_/X sky130_fd_sc_hd__or3_4
Xhold655 _1221_/Q vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _1204_/Q vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _1206_/Q vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _0794_/X vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold699 _1220_/Q vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_283_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout575_A _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0729__C _0729_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_342_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0761__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1035__A2 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0546__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput220 io_out_as1802[2] vssd1 vssd1 vccd1 vccd1 _0615_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_219_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput231 io_out_as1802[7] vssd1 vssd1 vccd1 vccd1 _0635_/B2 sky130_fd_sc_hd__buf_2
Xinput253 io_out_scrapcpu[27] vssd1 vssd1 vccd1 vccd1 _0716_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput242 io_out_scrapcpu[17] vssd1 vssd1 vccd1 vccd1 _0676_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_236_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput297 io_out_vliw[34] vssd1 vssd1 vccd1 vccd1 _0744_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput286 io_out_vliw[24] vssd1 vssd1 vccd1 vccd1 _0704_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput275 io_out_vliw[14] vssd1 vssd1 vccd1 vccd1 _0664_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_388_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput264 io_out_scrapcpu[4] vssd1 vssd1 vccd1 vccd1 _0624_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_383_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output494_A _0633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0537__A1 _0537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0514_ _0518_/A _0514_/B vssd1 vssd1 vccd1 vccd1 _0514_/X sky130_fd_sc_hd__and2_4
XFILLER_0_265_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_375_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_388_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0528__A1 _0528_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 hold463/A vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 hold9/X vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 hold430/A vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold485 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold496/A vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 hold45/X vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_337_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0700__B2 _0700_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold702_A _1111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_381_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_262_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_357_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0994_ _0795_/A _0996_/A hold630/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0994_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput502 _1245_/X vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_12
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput535 _0518_/X vssd1 vssd1 vccd1 vccd1 rst_8x305 sky130_fd_sc_hd__buf_12
XFILLER_0_300_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput524 _1265_/X vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_12
Xoutput513 _1255_/X vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_12
XFILLER_0_300_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput557 hold182/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput546 hold237/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_12
Xoutput568 hold272/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_238_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_374_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_307_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_367_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_348_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold271 _0927_/Y vssd1 vssd1 vccd1 vccd1 _1145_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _1100_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_348_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold293 _0891_/Y vssd1 vssd1 vccd1 vccd1 _1133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _0885_/Y vssd1 vssd1 vccd1 vccd1 _1131_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_244_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_111 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_133 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_358_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_166 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_155 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_144 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_380_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output457_A _1237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1262_ hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__clkbuf_1
Xinput6 cap_io_in[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_0_349_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1193_ _1204_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _1193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_392_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_352_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0977_ _0849_/A _0996_/A hold364/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0977_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0600__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_258_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput387 _0761_/X vssd1 vssd1 vccd1 vccd1 cap_addr[5] sky130_fd_sc_hd__buf_12
XFILLER_0_273_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput398 _1103_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[16] sky130_fd_sc_hd__buf_12
XFILLER_0_318_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0667__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_395_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0753__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout592 _0526_/A vssd1 vssd1 vccd1 vccd1 _0518_/B sky130_fd_sc_hd__buf_4
Xfanout581 _0506_/B vssd1 vssd1 vccd1 vccd1 _0674_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_244_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_334_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0900_ _1085_/A _0900_/B vssd1 vssd1 vccd1 vccd1 _0900_/Y sky130_fd_sc_hd__nor2_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0831_ _1065_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0831_/X sky130_fd_sc_hd__or2_1
XFILLER_0_299_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0762_ input7/X _1093_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0763_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0693_ _0693_/A _0693_/B _0693_/C vssd1 vssd1 vccd1 vccd1 _0693_/X sky130_fd_sc_hd__or3_4
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1245_ _1245_/A vssd1 vssd1 vccd1 vccd1 _1245_/X sky130_fd_sc_hd__buf_1
XFILLER_0_223_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1176_ _1214_/CLK _1176_/D vssd1 vssd1 vccd1 vccd1 _1176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_22 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_55 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_88 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_356_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_316_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_351_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0591__A2 hold82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1030_ _1028_/X hold575/X _1080_/B vssd1 vssd1 vccd1 vccd1 _1030_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_366_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_334_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput31 io_oeb_scrapcpu[21] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 io_oeb_scrapcpu[11] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0814_ hold274/X _0840_/A2 _0813_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0814_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput42 io_oeb_scrapcpu[31] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_287_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput53 io_oeb_scrapcpu[9] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_1
Xinput64 io_oeb_vliw[19] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0745_ _0745_/A _0745_/B _0745_/C vssd1 vssd1 vccd1 vccd1 _0745_/X sky130_fd_sc_hd__or3_4
Xinput97 io_oeb_z80[16] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_2
Xinput75 io_oeb_vliw[29] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
Xinput86 io_oeb_vliw[6] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0676_ _0676_/A1 _0732_/A2 _0696_/B1 _0676_/B2 vssd1 vssd1 vccd1 vccd1 _0677_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_283_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_295_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1159_ _1188_/CLK _1159_/D vssd1 vssd1 vccd1 vccd1 _1159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout618_A _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1047__B1 _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0573__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0759__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_292_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_261_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_388_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_388_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_356_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0530_ input47/X _0598_/A2 _0598_/B1 input83/X vssd1 vssd1 vccd1 vccd1 _0530_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_277_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output537_A _0508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1013_ _1015_/B hold583/X _1021_/A vssd1 vssd1 vccd1 vccd1 _1013_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold601 _0865_/X vssd1 vssd1 vccd1 vccd1 _0866_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 hold767/X vssd1 vssd1 vccd1 vccd1 _0999_/A sky130_fd_sc_hd__buf_1
XFILLER_0_303_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0728_ _0728_/A1 _0732_/A2 _0748_/B1 _0728_/B2 vssd1 vssd1 vccd1 vccd1 _0729_/C sky130_fd_sc_hd__a22o_1
Xhold645 _0858_/X vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _0964_/B vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 _0995_/Y vssd1 vssd1 vccd1 vccd1 _0996_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_330_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold656 _1081_/X vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _0810_/X vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 _0806_/X vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0659_ _0659_/A1 _0593_/A _0695_/B1 _0659_/B2 vssd1 vssd1 vccd1 vccd1 _0661_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold689 _1158_/Q vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_393_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0511__A_N hold76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_342_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0761__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0794__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_367_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0546__A2 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput210 io_out_as1802[20] vssd1 vssd1 vccd1 vccd1 _0687_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput221 io_out_as1802[30] vssd1 vssd1 vccd1 vccd1 _0727_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput232 io_out_as1802[8] vssd1 vssd1 vccd1 vccd1 _0639_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput254 io_out_scrapcpu[28] vssd1 vssd1 vccd1 vccd1 _0720_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput243 io_out_scrapcpu[18] vssd1 vssd1 vccd1 vccd1 _0680_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_236_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput287 io_out_vliw[25] vssd1 vssd1 vccd1 vccd1 _0708_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput276 io_out_vliw[15] vssd1 vssd1 vccd1 vccd1 _0668_/B2 sky130_fd_sc_hd__buf_2
Xinput265 io_out_scrapcpu[5] vssd1 vssd1 vccd1 vccd1 _0628_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput298 io_out_vliw[35] vssd1 vssd1 vccd1 vccd1 _0748_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_388_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_391_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_344_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output487_A _0745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0537__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0513_ _0860_/A _0515_/B vssd1 vssd1 vccd1 vccd1 _0513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_288_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_382_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold420 hold5/X vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0528__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold431 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 hold27/X vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 hold442/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 hold53/X vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold475/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_337_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold497 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_262_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_376_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_364_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_391_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0993_ hold629/X _0995_/B _0996_/A vssd1 vssd1 vccd1 vccd1 _0993_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput536 _0516_/X vssd1 vssd1 vccd1 vccd1 rst_as1802 sky130_fd_sc_hd__buf_12
XFILLER_0_288_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput525 _1266_/X vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_12
Xoutput514 _1256_/X vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_12
Xoutput503 _1246_/X vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_12
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput558 hold179/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput547 hold191/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput569 hold310/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XFILLER_0_300_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0694__B2 _0694_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0592__A _0592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0997__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_363_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout600_A hold82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold109_A _0592_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold250 hold391/X vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__clkbuf_2
Xhold261 hold669/X vssd1 vssd1 vccd1 vccd1 _1100_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold283 hold751/X vssd1 vssd1 vccd1 vccd1 _1078_/C sky130_fd_sc_hd__buf_1
Xhold294 hold655/X vssd1 vssd1 vccd1 vccd1 _1080_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold396/X vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_348_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0767__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_364_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_112 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_123 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_134 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_101 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_167 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_156 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_145 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_178 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_373_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_258_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1261_ _1261_/A vssd1 vssd1 vccd1 vccd1 _1261_/X sky130_fd_sc_hd__buf_1
Xinput7 cap_io_in[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_0_274_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1192_ _1204_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _1192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_389_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0676__B2 _0676_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0843__C _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ hold363/X _0979_/B _0996_/A vssd1 vssd1 vccd1 vccd1 _0976_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_360_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0600__A1 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput399 _1104_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[17] sky130_fd_sc_hd__buf_12
Xoutput388 _0763_/X vssd1 vssd1 vccd1 vccd1 cap_addr[6] sky130_fd_sc_hd__buf_12
XFILLER_0_226_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0667__A1 _0667_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0667__B2 _0667_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_276_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_291_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout582 hold105/X vssd1 vssd1 vccd1 vccd1 _0506_/B sky130_fd_sc_hd__buf_6
Xfanout593 _0683_/B1 vssd1 vssd1 vccd1 vccd1 _0695_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__0658__B2 _0658_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_386_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0830_ hold318/X _0840_/A2 _0829_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0830_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_342_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0761_ _0767_/A _0767_/B _0761_/C vssd1 vssd1 vccd1 vccd1 _0761_/X sky130_fd_sc_hd__and3_4
XFILLER_0_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output567_A hold301/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0692_ _0692_/A1 _0732_/A2 _0748_/B1 _0692_/B2 vssd1 vssd1 vccd1 vccd1 _0693_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_267_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0594__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_270_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1244_ _1244_/A vssd1 vssd1 vccd1 vccd1 _1244_/X sky130_fd_sc_hd__buf_1
XFILLER_0_223_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1175_ _1175_/CLK _1175_/D vssd1 vssd1 vccd1 vccd1 _1175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_377_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1074__A1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_34 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_67 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0959_ _1082_/A _0996_/A hold201/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0959_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_258_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0585__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_258_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_273_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_254_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold343_A hold76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_386_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_374_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 io_in_0 vssd1 vssd1 vccd1 vccd1 _1267_/A sky130_fd_sc_hd__clkbuf_8
Xinput21 io_oeb_scrapcpu[12] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
X_0813_ _0813_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0813_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput43 io_oeb_scrapcpu[32] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_287_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput32 io_oeb_scrapcpu[22] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_1
Xinput54 io_oeb_vliw[0] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0744_ _0744_/A1 _0508_/B _0748_/B1 _0744_/B2 vssd1 vssd1 vccd1 vccd1 _0745_/C sky130_fd_sc_hd__a22o_1
Xinput98 io_oeb_z80[17] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0567__B1 _0526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput87 io_oeb_vliw[7] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_1
Xinput76 io_oeb_vliw[2] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_1
Xinput65 io_oeb_vliw[1] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0675_ _0675_/A1 _0514_/B _0683_/B1 _0675_/B2 vssd1 vssd1 vccd1 vccd1 _0677_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_296_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1158_ _1167_/CLK _1158_/D vssd1 vssd1 vccd1 vccd1 _1158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1089_ _1205_/CLK _1089_/D vssd1 vssd1 vccd1 vccd1 _1089_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_353_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_306_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0558__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0759__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0775__A _0775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_372_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold725_A _1181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_372_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output432_A _1248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_379_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1012_ _1016_/C _1012_/B vssd1 vssd1 vccd1 vccd1 _1012_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 _0866_/X vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_330_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0727_ _0727_/A1 _0747_/A2 _0516_/B _0727_/B2 vssd1 vssd1 vccd1 vccd1 _0729_/B sky130_fd_sc_hd__a22o_1
Xhold635 _0962_/X vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 _0996_/Y vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 _0987_/Y vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _1189_/Q vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _1214_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold679 _1197_/Q vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _1203_/Q vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
X_0658_ _0658_/A1 _0674_/A2 _0674_/B1 _0658_/B2 vssd1 vssd1 vccd1 vccd1 _0661_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_216_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0589_ hold77/X _0589_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__or2_4
XFILLER_0_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_338_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_342_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_338_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold306_A _1101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput211 io_out_as1802[21] vssd1 vssd1 vccd1 vccd1 _0691_/B2 sky130_fd_sc_hd__buf_2
Xinput200 io_out_as1802[11] vssd1 vssd1 vccd1 vccd1 _0651_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_274_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput222 io_out_as1802[31] vssd1 vssd1 vccd1 vccd1 _0731_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput233 io_out_as1802[9] vssd1 vssd1 vccd1 vccd1 _0643_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput244 io_out_scrapcpu[19] vssd1 vssd1 vccd1 vccd1 _0684_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_234_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput288 io_out_vliw[26] vssd1 vssd1 vccd1 vccd1 _0712_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput277 io_out_vliw[16] vssd1 vssd1 vccd1 vccd1 _0672_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_388_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput255 io_out_scrapcpu[29] vssd1 vssd1 vccd1 vccd1 _0724_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput266 io_out_scrapcpu[6] vssd1 vssd1 vccd1 vccd1 _0632_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0703__B1 _0515_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput299 io_out_vliw[3] vssd1 vssd1 vccd1 vccd1 _0620_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_388_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output382_A _0751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0512_ hold76/X hold99/X _0868_/A vssd1 vssd1 vccd1 vccd1 _0512_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_390_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_388_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 hold800/X vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold17/X vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 hold454/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 hold487/A vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 hold43/X vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold498 hold57/X vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_337_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_271_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_341_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_262_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_391_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_372_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ _0992_/A _0992_/B vssd1 vssd1 vccd1 vccd1 _0995_/B sky130_fd_sc_hd__and2_1
XFILLER_0_317_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput526 _1267_/X vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_12
Xoutput515 _1257_/X vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_12
Xoutput504 _1247_/X vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_12
XFILLER_0_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput537 _0508_/X vssd1 vssd1 vccd1 vccd1 rst_scrapcpu sky130_fd_sc_hd__buf_12
XFILLER_0_285_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput559 hold185/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput548 hold197/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_238_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold240 hold410/X vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__clkbuf_2
Xhold251 _0867_/X vssd1 vssd1 vccd1 vccd1 _1126_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold395/X vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_348_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold284 hold752/X vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _0839_/X vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _0875_/X vssd1 vssd1 vccd1 vccd1 _1128_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_244_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0767__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_364_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_102 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_124 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_113 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_380_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_157 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_146 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_135 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_380_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_168 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1260_ _1260_/A vssd1 vssd1 vccd1 vccd1 _1260_/X sky130_fd_sc_hd__buf_1
Xinput8 cap_io_in[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_0_274_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output512_A _1254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1191_ _1204_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _1191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_349_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0975_ _0983_/A _0983_/B _1017_/A vssd1 vssd1 vccd1 vccd1 _0979_/B sky130_fd_sc_hd__and3_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_360_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1010__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0868__A _0868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput389 _0765_/X vssd1 vssd1 vccd1 vccd1 cap_addr[7] sky130_fd_sc_hd__buf_12
XFILLER_0_226_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0587__B _0587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0667__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_355_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_395_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1077__C1 _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_355_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_363_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_291_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout583 _0590_/A2 vssd1 vssd1 vccd1 vccd1 _0605_/A2 sky130_fd_sc_hd__buf_6
Xfanout594 _0515_/Y vssd1 vssd1 vccd1 vccd1 _0683_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_391_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0830__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0760_ input6/X _1092_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0761_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output462_A _0653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0691_ _0691_/A1 _0747_/A2 _0695_/B1 _0691_/B2 vssd1 vssd1 vccd1 vccd1 _0693_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_267_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_263_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1243_ _1243_/A vssd1 vssd1 vccd1 vccd1 _1243_/X sky130_fd_sc_hd__buf_1
XFILLER_0_263_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1174_ _1180_/CLK _1174_/D vssd1 vssd1 vccd1 vccd1 _1174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_392_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0806__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_392_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_79 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0958_ _0967_/A _0996_/A vssd1 vssd1 vccd1 vccd1 _0958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_68 hold35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0585__A1 _0585_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0889_ hold267/X _0776_/A hold605/A _0995_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0889_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_273_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0812__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_249_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_255_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_374_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput22 io_oeb_scrapcpu[13] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
XFILLER_0_181_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0812_ hold299/X _0840_/A2 _0811_/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0812_/X sky130_fd_sc_hd__o211a_1
Xinput11 io_oeb_6502 vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 io_oeb_scrapcpu[33] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
Xinput33 io_oeb_scrapcpu[23] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
Xinput55 io_oeb_vliw[10] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0743_ _0743_/A1 _0747_/A2 _0516_/B _0743_/B2 vssd1 vssd1 vccd1 vccd1 _0745_/B sky130_fd_sc_hd__a22o_1
Xinput77 io_oeb_vliw[30] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
Xinput66 io_oeb_vliw[20] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0567__B2 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput88 io_oeb_vliw[8] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput99 io_oeb_z80[18] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_2
X_0674_ _0674_/A1 _0674_/A2 _0674_/B1 _0674_/B2 vssd1 vssd1 vccd1 vccd1 _0677_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_228_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0849__C _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1157_ _1157_/CLK _1157_/D vssd1 vssd1 vccd1 vccd1 _1157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1088_ _1188_/CLK _1088_/D vssd1 vssd1 vccd1 vccd1 _1088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0558__A1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0730__B2 _0730_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_292_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0669__C _0669_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output425_A _1241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1011_ _1016_/C _1012_/B vssd1 vssd1 vccd1 vccd1 _1015_/B sky130_fd_sc_hd__and2_1
XFILLER_0_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_260_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_387_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold603 _1223_/Q vssd1 vssd1 vccd1 vccd1 _0841_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_330_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0726_ _0726_/A1 _0746_/A2 _0746_/B1 _0726_/B2 vssd1 vssd1 vccd1 vccd1 _0729_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold636 _1190_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _0997_/X vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 _0989_/Y vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold647 hold73/X vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _1056_/X vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 _0804_/X vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
X_0657_ _0657_/A _0657_/B _0657_/C vssd1 vssd1 vccd1 vccd1 _0657_/X sky130_fd_sc_hd__or3_4
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0588_ _0588_/A1 _0505_/A hold87/A input74/X _0587_/X vssd1 vssd1 vccd1 vccd1 _0589_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0712__B2 _0712_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1209_ _1215_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 _1209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_259_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_274_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput201 io_out_as1802[12] vssd1 vssd1 vccd1 vccd1 _0655_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_274_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput223 io_out_as1802[32] vssd1 vssd1 vccd1 vccd1 _0735_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput212 io_out_as1802[22] vssd1 vssd1 vccd1 vccd1 _0695_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput245 io_out_scrapcpu[1] vssd1 vssd1 vccd1 vccd1 _0612_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput234 io_out_scrapcpu[0] vssd1 vssd1 vccd1 vccd1 _0608_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0703__A1 _0703_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput278 io_out_vliw[17] vssd1 vssd1 vccd1 vccd1 _0676_/B2 sky130_fd_sc_hd__buf_2
Xinput267 io_out_scrapcpu[7] vssd1 vssd1 vccd1 vccd1 _0636_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput256 io_out_scrapcpu[2] vssd1 vssd1 vccd1 vccd1 _0616_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0703__B2 _0703_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput289 io_out_vliw[27] vssd1 vssd1 vccd1 vccd1 _0716_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_388_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_388_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1167_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_369_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_312_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0511_ hold76/X hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__and2b_1
XANTENNA_output542_A hold291/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_382_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold400 hold798/X vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 hold733/X vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold433 hold433/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold762/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 hold21/X vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0709_ _0709_/A _0709_/B _0709_/C vssd1 vssd1 vccd1 vccd1 _0709_/X sky130_fd_sc_hd__or3_4
Xhold477 hold39/X vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/A vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_378_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output492_A _0625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0991_ _0992_/A _0992_/B vssd1 vssd1 vccd1 vccd1 _0991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput527 hold649/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__buf_6
Xoutput516 _1258_/X vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_12
Xoutput505 _1248_/X vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_12
Xoutput538 _0510_/X vssd1 vssd1 vccd1 vccd1 rst_vliw sky130_fd_sc_hd__buf_12
XFILLER_0_285_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput549 hold206/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_0_238_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0679__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold230 _0950_/Y vssd1 vssd1 vccd1 vccd1 _0951_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _0899_/Y vssd1 vssd1 vccd1 vccd1 _0900_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold252 hold392/X vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold285 _1077_/X vssd1 vssd1 vccd1 vccd1 _1186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold526/X vssd1 vssd1 vccd1 vccd1 _1118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _1105_/Q vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _0887_/Y vssd1 vssd1 vccd1 vccd1 _0888_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_364_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_103 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_114 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_158 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_147 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_136 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0783__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_380_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_169 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_380_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_381_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_267_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_267_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0958__B _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0677__C _0677_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1190_ _1204_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 _1190_/Q sky130_fd_sc_hd__dfxtp_1
Xinput9 cap_io_in[8] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_4
XFILLER_0_389_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_290_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0974_ _1160_/Q _1017_/A _0983_/B vssd1 vssd1 vccd1 vccd1 _0974_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0868__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_328_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_370_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1001__B1 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_291_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_272_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout584 hold105/X vssd1 vssd1 vccd1 vccd1 _0590_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout573 _1021_/A vssd1 vssd1 vccd1 vccd1 _0996_/A sky130_fd_sc_hd__buf_4
XFILLER_0_378_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout595 _0515_/Y vssd1 vssd1 vccd1 vccd1 _0516_/B sky130_fd_sc_hd__clkbuf_8
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0690_ _0690_/A1 _0746_/A2 _0746_/B1 _0690_/B2 vssd1 vssd1 vccd1 vccd1 _0693_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_267_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output455_A _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1242_ _1242_/A vssd1 vssd1 vccd1 vccd1 _1242_/X sky130_fd_sc_hd__buf_1
XFILLER_0_256_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1173_ _1180_/CLK _1173_/D vssd1 vssd1 vccd1 vccd1 _1173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_14 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_47 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_360_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_58 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0957_ _1082_/B _0957_/B vssd1 vssd1 vccd1 vccd1 _0957_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_69 hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_360_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0585__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0888_ _1085_/A _0888_/B vssd1 vssd1 vccd1 vccd1 _0888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_254_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold329_A _1102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_289_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_386_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 io_oeb_8x305[0] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
XFILLER_0_342_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output572_A hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0811_ _0811_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0811_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput45 io_oeb_scrapcpu[34] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
Xinput34 io_oeb_scrapcpu[24] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
X_0742_ _0742_/A1 _0746_/A2 _0746_/B1 _0742_/B2 vssd1 vssd1 vccd1 vccd1 _0745_/A sky130_fd_sc_hd__a22o_1
Xinput23 io_oeb_scrapcpu[14] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
XFILLER_0_181_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput78 io_oeb_vliw[31] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
Xinput67 io_oeb_vliw[21] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
Xinput56 io_oeb_vliw[11] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_1
Xinput89 io_oeb_vliw[9] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0673_ _0673_/A _0673_/B _0673_/C vssd1 vssd1 vccd1 vccd1 _0673_/X sky130_fd_sc_hd__or3_4
XFILLER_0_255_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_373_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1225_ _1225_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 _1225_/Q sky130_fd_sc_hd__dfxtp_1
X_1156_ _1167_/CLK _1156_/D vssd1 vssd1 vccd1 vccd1 _1156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1087_ _1205_/CLK _1087_/D vssd1 vssd1 vccd1 vccd1 _1087_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0963__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1233__A _1233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_372_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0791__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_371_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_324_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_292_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_292_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_379_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0685__C _0685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_394_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1010_ _0803_/A _1021_/A hold588/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _1010_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_282_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0788__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0725_ _0725_/A _0725_/B _0725_/C vssd1 vssd1 vccd1 vccd1 _0725_/X sky130_fd_sc_hd__or3_4
Xhold626 _1087_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 _0851_/X vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__buf_1
Xhold615 _0990_/X vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_330_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0656_ _0656_/A1 _0660_/A2 _0696_/B1 _0656_/B2 vssd1 vssd1 vccd1 vccd1 _0657_/C sky130_fd_sc_hd__a22o_1
Xhold648 _0518_/A vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _1082_/X vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 _1156_/Q vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
X_0587_ hold86/X _0587_/B hold99/A vssd1 vssd1 vccd1 vccd1 _0587_/X sky130_fd_sc_hd__or3b_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1208_ _1215_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 _1208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1139_ _1189_/CLK _1139_/D vssd1 vssd1 vccd1 vccd1 _1139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput202 io_out_as1802[13] vssd1 vssd1 vccd1 vccd1 _0659_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_219_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput224 io_out_as1802[33] vssd1 vssd1 vccd1 vccd1 _0739_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput213 io_out_as1802[23] vssd1 vssd1 vccd1 vccd1 _0699_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput235 io_out_scrapcpu[10] vssd1 vssd1 vccd1 vccd1 _0648_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_274_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput279 io_out_vliw[18] vssd1 vssd1 vccd1 vccd1 _0680_/B2 sky130_fd_sc_hd__buf_2
Xinput257 io_out_scrapcpu[30] vssd1 vssd1 vccd1 vccd1 _0728_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput246 io_out_scrapcpu[20] vssd1 vssd1 vccd1 vccd1 _0688_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput268 io_out_scrapcpu[8] vssd1 vssd1 vccd1 vccd1 _0640_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_376_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_312_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0510_ _0518_/A _0510_/B vssd1 vssd1 vccd1 vccd1 _0510_/X sky130_fd_sc_hd__and2_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output535_A _0518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_379_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0630__B2 _0630_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold401 hold787/X vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold412 hold745/X vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__buf_1
Xhold423 hold7/X vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold445 hold445/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dlygate4sd3_1
X_0708_ _0708_/A1 _0732_/A2 _0748_/B1 _0708_/B2 vssd1 vssd1 vccd1 vccd1 _0709_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_256_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold478 hold478/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 hold29/X vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
X_0639_ _0639_/A1 _0514_/B _0695_/B1 _0639_/B2 vssd1 vssd1 vccd1 vccd1 _0641_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold489 hold49/X vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_378_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_247_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0688__B2 _0688_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0990_ _0793_/A _0996_/A hold614/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0990_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_372_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output485_A _0737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0612__B2 _0612_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput517 _1232_/X vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_12
Xoutput506 hold84/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__buf_6
XFILLER_0_288_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput539 _0506_/X vssd1 vssd1 vccd1 vccd1 rst_z80 sky130_fd_sc_hd__buf_12
Xoutput528 _1233_/X vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_12
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0500__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0679__A1 _0679_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0679__B2 _0679_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_367_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0603__A1 _0603_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold220 hold382/X vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_198_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold231 _0951_/Y vssd1 vssd1 vccd1 vccd1 _1153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _0900_/Y vssd1 vssd1 vccd1 vccd1 _1136_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold253 _0855_/X vssd1 vssd1 vccd1 vccd1 _1123_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold286 hold749/X vssd1 vssd1 vccd1 vccd1 _1072_/A sky130_fd_sc_hd__buf_1
Xhold275 hold706/X vssd1 vssd1 vccd1 vccd1 _1105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _0888_/Y vssd1 vssd1 vccd1 vccd1 _1132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold411/X vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__clkbuf_2
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_364_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_104 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_115 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1241__A _1241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_126 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_148 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_137 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_380_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_159 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_307_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0693__C _0693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0973_ _0847_/A _0996_/A _0972_/Y _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0597__B1 hold95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0521__B1 _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_395_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1077__A1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_336_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_351_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1236__A _1236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0760__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 _1076_/B vssd1 vssd1 vccd1 vccd1 _1021_/A sky130_fd_sc_hd__buf_4
Xfanout585 _0505_/Y vssd1 vssd1 vccd1 vccd1 _0746_/A2 sky130_fd_sc_hd__buf_4
Xfanout596 _0593_/A vssd1 vssd1 vccd1 vccd1 _0514_/B sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_386_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_354_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_267_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output448_A hold96/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1241_ _1241_/A vssd1 vssd1 vccd1 vccd1 _1241_/X sky130_fd_sc_hd__buf_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1172_ _1180_/CLK _1172_/D vssd1 vssd1 vccd1 vccd1 _1172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1059__A1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_48 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_360_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_59 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0956_ _1082_/B _0957_/B vssd1 vssd1 vccd1 vccd1 _0956_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_360_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0887_ hold262/X _0880_/A _0886_/X vssd1 vssd1 vccd1 vccd1 _0887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_383_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_336_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0789__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_386_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_386_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_255_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output398_A _1103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 io_oeb_8x305[1] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_342_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0810_ hold308/X _0810_/A2 _0809_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0810_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 io_oeb_scrapcpu[35] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
Xinput35 io_oeb_scrapcpu[25] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
X_0741_ _0741_/A _0741_/B _0741_/C vssd1 vssd1 vccd1 vccd1 _0741_/X sky130_fd_sc_hd__or3_4
Xinput24 io_oeb_scrapcpu[15] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
XFILLER_0_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput79 io_oeb_vliw[32] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
Xinput68 io_oeb_vliw[22] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
Xinput57 io_oeb_vliw[12] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_1
XANTENNA_output565_A hold257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0672_ _0672_/A1 _0732_/A2 _0696_/B1 _0672_/B2 vssd1 vssd1 vccd1 vccd1 _0673_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_296_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_296_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1224_ _1224_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _1224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_315_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1155_ _1214_/CLK _1155_/D vssd1 vssd1 vccd1 vccd1 _1155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1086_ _1214_/CLK _1086_/D vssd1 vssd1 vccd1 vccd1 _1086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0939_ _1036_/A _0939_/B vssd1 vssd1 vccd1 vccd1 _0939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_286_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout596_A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0715__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_371_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_252_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_282_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_347_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0724_ _0724_/A1 _0732_/A2 _0748_/B1 _0724_/B2 vssd1 vssd1 vccd1 vccd1 _0725_/C sky130_fd_sc_hd__a22o_1
XANTENNA__0503__A hold76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold627 _0778_/X vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold605 hold605/A vssd1 vssd1 vccd1 vccd1 _0957_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 hold616/A vssd1 vssd1 vccd1 vccd1 _1164_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_268_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0655_ _0655_/A1 _0514_/B _0695_/B1 _0655_/B2 vssd1 vssd1 vccd1 vccd1 _0657_/B sky130_fd_sc_hd__a22o_1
Xhold649 hold74/X vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _1083_/X vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_283_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0586_ input37/X _0598_/A2 _0586_/B1 input73/X _0585_/X vssd1 vssd1 vccd1 vccd1 _1258_/A
+ sky130_fd_sc_hd__a221o_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_243_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1207_ _1215_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 _1207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1138_ _1189_/CLK _1138_/D vssd1 vssd1 vccd1 vccd1 _1138_/Q sky130_fd_sc_hd__dfxtp_1
X_1069_ _1072_/B hold554/X _1080_/B vssd1 vssd1 vccd1 vccd1 _1069_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0881__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_353_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_A _0507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput225 io_out_as1802[34] vssd1 vssd1 vccd1 vccd1 _0743_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput214 io_out_as1802[24] vssd1 vssd1 vccd1 vccd1 _0703_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput203 io_out_as1802[14] vssd1 vssd1 vccd1 vccd1 _0663_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput236 io_out_scrapcpu[11] vssd1 vssd1 vccd1 vccd1 _0652_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_274_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1244__A _1244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput258 io_out_scrapcpu[31] vssd1 vssd1 vccd1 vccd1 _0732_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput247 io_out_scrapcpu[21] vssd1 vssd1 vccd1 vccd1 _0692_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput269 io_out_scrapcpu[9] vssd1 vssd1 vccd1 vccd1 _0644_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_236_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_242_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output430_A _1246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_379_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__buf_1
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0863__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_390_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold402 hold735/X vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ _0707_/A1 _0747_/A2 _0516_/B _0707_/B2 vssd1 vssd1 vccd1 vccd1 _0709_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold424 hold424/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold748/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold435 hold15/X vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 hold37/X vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 hold457/A vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0638_ _0638_/A1 _0674_/A2 _0674_/B1 _0638_/B2 vssd1 vssd1 vccd1 vccd1 _0641_/A sky130_fd_sc_hd__a22o_1
Xhold479 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0569_ _0569_/A _0569_/B _0569_/C vssd1 vssd1 vccd1 vccd1 _1250_/A sky130_fd_sc_hd__or3_4
XFILLER_0_216_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_353_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_366_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1239__A _1239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0797__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_394_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_357_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output478_A _0713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput518 hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__buf_6
Xoutput507 _1249_/X vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_12
XFILLER_0_151_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1022__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput529 _1234_/X vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_12
XFILLER_0_238_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_261_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_348_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold210 _0917_/Y vssd1 vssd1 vccd1 vccd1 _0918_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_288_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold232 hold406/X vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__clkbuf_2
Xhold243 _1120_/Q vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _0859_/X vssd1 vssd1 vccd1 vccd1 _1124_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold287 hold750/X vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _1108_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold407/X vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__clkbuf_2
Xhold265 _1095_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold298 _0863_/X vssd1 vssd1 vccd1 vccd1 _1125_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_364_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_149 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_127 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_138 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_380_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_354_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_354_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_275_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_290_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ _0996_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_299_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0597__A1 _0597_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_336_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0824__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0588__B2 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0588__A1 _0588_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_375_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout575 _1076_/B vssd1 vssd1 vccd1 vccd1 _1080_/B sky130_fd_sc_hd__buf_4
Xfanout597 _0593_/A vssd1 vssd1 vccd1 vccd1 _0747_/A2 sky130_fd_sc_hd__buf_4
Xfanout586 _0882_/X vssd1 vssd1 vccd1 vccd1 _0952_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_225_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1252__A _1252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_386_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_386_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0579__A1 _0579_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1240_ _1240_/A vssd1 vssd1 vccd1 vccd1 _1240_/X sky130_fd_sc_hd__buf_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1171_ _1205_/CLK _1171_/D vssd1 vssd1 vccd1 vccd1 _1171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_290_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_263_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_304_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0806__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0506__A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_16 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold78_A hold78/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0955_ _0955_/A _0955_/B vssd1 vssd1 vccd1 vccd1 _0955_/X sky130_fd_sc_hd__and2_1
XFILLER_0_360_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0886_ hold166/X _0776_/A hold605/A _0992_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0886_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0742__A1 _0742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0742__B2 _0742_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_368_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_368_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1222__D hold6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_383_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_336_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1247__A _1247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_386_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_272_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_255_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 io_oeb_8x305[2] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_342_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0740_ _0740_/A1 _0508_/B _0748_/B1 _0740_/B2 vssd1 vssd1 vccd1 vccd1 _0741_/C sky130_fd_sc_hd__a22o_1
Xinput36 io_oeb_scrapcpu[26] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
Xinput25 io_oeb_scrapcpu[16] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 io_oeb_scrapcpu[3] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput69 io_oeb_vliw[23] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
Xinput58 io_oeb_vliw[13] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_1
XANTENNA_output460_A _0645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0671_ _0671_/A1 _0514_/B _0683_/B1 _0671_/B2 vssd1 vssd1 vccd1 vccd1 _0673_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_220_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0996__A _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0724__B2 _0724_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1223_ _1224_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _1223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_251_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1154_ _1154_/CLK _1154_/D vssd1 vssd1 vccd1 vccd1 _1154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1085_ _1085_/A _1085_/B vssd1 vssd1 vccd1 vccd1 _1085_/X sky130_fd_sc_hd__or2_1
XFILLER_0_365_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0938_ hold185/X _0953_/A2 _0937_/X vssd1 vssd1 vccd1 vccd1 _0938_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0869_ hold333/X _0776_/A hold605/A _0983_/A _0868_/X vssd1 vssd1 vccd1 vccd1 _0869_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_286_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0715__A1 _0715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0715__B2 _0715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_242_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_324_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0651__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_324_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0706__B2 _0706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_268_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0723_ _0723_/A1 _0747_/A2 _0516_/B _0723_/B2 vssd1 vssd1 vccd1 vccd1 _0725_/B sky130_fd_sc_hd__a22o_1
Xhold606 _0876_/X vssd1 vssd1 vccd1 vccd1 _0877_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 hold776/X vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__buf_1
XFILLER_0_311_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0654_ _0654_/A1 _0674_/A2 _0674_/B1 _0654_/B2 vssd1 vssd1 vccd1 vccd1 _0657_/A sky130_fd_sc_hd__a22o_1
Xhold628 hold777/X vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__buf_1
Xhold639 _1160_/Q vssd1 vssd1 vccd1 vccd1 _0983_/A sky130_fd_sc_hd__clkbuf_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0585_ _0585_/A1 _0506_/B _0683_/B1 _0526_/X vssd1 vssd1 vccd1 vccd1 _0585_/X sky130_fd_sc_hd__a211o_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1206_ _1215_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 _1206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1137_ _1189_/CLK _1137_/D vssd1 vssd1 vccd1 vccd1 _1137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1068_ _1071_/A _1071_/D _1071_/B vssd1 vssd1 vccd1 vccd1 _1068_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput226 io_out_as1802[35] vssd1 vssd1 vccd1 vccd1 _0747_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput215 io_out_as1802[25] vssd1 vssd1 vccd1 vccd1 _0707_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput204 io_out_as1802[15] vssd1 vssd1 vccd1 vccd1 _0667_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput259 io_out_scrapcpu[32] vssd1 vssd1 vccd1 vccd1 _0736_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput248 io_out_scrapcpu[22] vssd1 vssd1 vccd1 vccd1 _0696_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput237 io_out_scrapcpu[12] vssd1 vssd1 vccd1 vccd1 _0656_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_242_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_383_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output423_A _1239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_379_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0615__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_343_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0514__A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0706_ _0706_/A1 _0746_/A2 _0746_/B1 _0706_/B2 vssd1 vssd1 vccd1 vccd1 _0709_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_187_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 hold796/X vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 hold1/X vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold425 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 hold436/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 hold19/X vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold458 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dlygate4sd3_1
X_0637_ _0637_/A _0637_/B _0637_/C vssd1 vssd1 vccd1 vccd1 _0637_/X sky130_fd_sc_hd__or3_4
XFILLER_0_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0568_ _0568_/A1 _0605_/A2 _0604_/A2 input28/X vssd1 vssd1 vccd1 vccd1 _0569_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_271_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0499_ _0860_/A vssd1 vssd1 vccd1 vccd1 _0517_/B sky130_fd_sc_hd__inv_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1255__A _1255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_394_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_327_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_263_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_372_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_308_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput508 _1250_/X vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput519 _1260_/X vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0509__A hold99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_382_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold211 _0918_/Y vssd1 vssd1 vccd1 vccd1 _1142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 hold659/X vssd1 vssd1 vccd1 vccd1 _0967_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1205_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold244 hold98/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _0920_/Y vssd1 vssd1 vccd1 vccd1 _0921_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold408/X vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold277 hold708/X vssd1 vssd1 vccd1 vccd1 _1108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _0896_/Y vssd1 vssd1 vccd1 vccd1 _0897_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 hold688/X vssd1 vssd1 vccd1 vccd1 _1095_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold288 _1074_/X vssd1 vssd1 vccd1 vccd1 _1185_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _1104_/Q vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1225__D hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_128 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_117 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 hold47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_290_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_364_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_372_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0971_ _0983_/A _1017_/A vssd1 vssd1 vccd1 vccd1 _0971_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output490_A _0617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_372_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_285_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_334_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_304_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout598 _0513_/Y vssd1 vssd1 vccd1 vccd1 _0593_/A sky130_fd_sc_hd__buf_4
Xfanout587 _0882_/X vssd1 vssd1 vccd1 vccd1 _0934_/C1 sky130_fd_sc_hd__buf_2
Xfanout576 _0957_/X vssd1 vssd1 vccd1 vccd1 _1076_/B sky130_fd_sc_hd__buf_2
XFILLER_0_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_386_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_386_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_263_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1170_ _1205_/CLK _1170_/D vssd1 vssd1 vccd1 vccd1 _1170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_377_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_17 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0506__B _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0954_ _1085_/A _0954_/B vssd1 vssd1 vccd1 vccd1 _0954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_144_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0885_ _1085_/A _0885_/B vssd1 vssd1 vccd1 vccd1 _0885_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_103_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_360_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0990__A2 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0966__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_386_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1263__A hold89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_359_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 io_oeb_8x305[3] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_330_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 io_oeb_scrapcpu[27] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
Xinput26 io_oeb_scrapcpu[17] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_342_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput48 io_oeb_scrapcpu[4] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
X_0670_ _0670_/A1 _0674_/A2 _0674_/B1 _0670_/B2 vssd1 vssd1 vccd1 vccd1 _0673_/A sky130_fd_sc_hd__a22o_1
Xinput59 io_oeb_vliw[14] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_1
XANTENNA_output453_A _1233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1222_ _1224_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _1222_/Q sky130_fd_sc_hd__dfxtp_1
X_1153_ _1187_/CLK _1153_/D vssd1 vssd1 vccd1 vccd1 _1153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_254_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1084_ hold73/X hold374/X _1084_/S vssd1 vssd1 vccd1 vccd1 _1084_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_365_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0517__A hold99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0660__B2 _0660_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0937_ hold318/X _0952_/A2 _0952_/B1 _1060_/C _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0937_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0868_ _0868_/A _1082_/C vssd1 vssd1 vccd1 vccd1 _0868_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0799_ _0799_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0799_/X sky130_fd_sc_hd__or2_1
XFILLER_0_286_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0715__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_388_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0651__B2 _0651_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0651__A1 _0651_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1258__A _1258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_379_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0890__A1 hold291/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_355_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0642__B2 _0642_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_370_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output570_A hold316/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0722_ _0722_/A1 _0746_/A2 _0746_/B1 _0722_/B2 vssd1 vssd1 vccd1 vccd1 _0725_/A sky130_fd_sc_hd__a22o_1
Xhold607 _0877_/X vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _1003_/Y vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0653_ _0653_/A _0653_/B _0653_/C vssd1 vssd1 vccd1 vccd1 _0653_/X sky130_fd_sc_hd__or3_4
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold629 _0991_/Y vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_283_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0584_ input72/X _0586_/B1 _0574_/X _0583_/X vssd1 vssd1 vccd1 vccd1 _1257_/A sky130_fd_sc_hd__a211o_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_371_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1205_ _1205_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 _1205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1136_ _1189_/CLK _1136_/D vssd1 vssd1 vccd1 vccd1 _1136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1067_ _1071_/A _1071_/B _1071_/D vssd1 vssd1 vccd1 vccd1 _1072_/B sky130_fd_sc_hd__and3_1
XANTENNA__0881__A1 hold316/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_306_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_367_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput216 io_out_as1802[26] vssd1 vssd1 vccd1 vccd1 _0711_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput205 io_out_as1802[16] vssd1 vssd1 vccd1 vccd1 _0671_/B2 sky130_fd_sc_hd__buf_2
Xinput227 io_out_as1802[3] vssd1 vssd1 vccd1 vccd1 _0619_/B2 sky130_fd_sc_hd__buf_2
Xinput249 io_out_scrapcpu[23] vssd1 vssd1 vccd1 vccd1 _0700_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput238 io_out_scrapcpu[13] vssd1 vssd1 vccd1 vccd1 _0660_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_242_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_242_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_384_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_337_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0624__B2 _0624_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0560__B1 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_379_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0863__A1 hold297/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0615__A1 _0615_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0615__B2 _0615_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_390_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_343_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0514__B _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0705_ _0705_/A _0705_/B _0705_/C vssd1 vssd1 vccd1 vccd1 _0705_/X sky130_fd_sc_hd__or3_4
Xhold404 hold797/X vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold426 hold11/X vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold437 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 hold31/X vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 hold448/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0636_ _0636_/A1 _0660_/A2 _0696_/B1 _0636_/B2 vssd1 vssd1 vccd1 vccd1 _0637_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0567_ input64/X _0586_/B1 _0526_/A input16/X vssd1 vssd1 vccd1 vccd1 _0569_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_271_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _1175_/CLK _1119_/D vssd1 vssd1 vccd1 vccd1 _1119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_366_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_381_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0606__A1 _0606_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0606__B2 _0606_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_302_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout614_A _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput509 _1251_/X vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_12
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_390_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 _0958_/Y vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold234 _0921_/Y vssd1 vssd1 vccd1 vccd1 _1143_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _0914_/Y vssd1 vssd1 vccd1 vccd1 _0915_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold212 _1094_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold278 _1115_/Q vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold698/X vssd1 vssd1 vccd1 vccd1 _1073_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _0897_/Y vssd1 vssd1 vccd1 vccd1 _1135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold763/X vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__buf_1
X_0619_ _0619_/A1 _0514_/B _0695_/B1 _0619_/B2 vssd1 vssd1 vccd1 vccd1 _0621_/B sky130_fd_sc_hd__a22o_1
Xhold289 _1107_/Q vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_107 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_118 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_366_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_322_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1266__A _1266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold790 _1139_/Q vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_290_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_275_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_290_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_372_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0970_ _0845_/A _1021_/A hold537/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_372_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output483_A _0729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0754__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_304_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0993__B1 _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_359_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_375_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout599 hold82/X vssd1 vssd1 vccd1 vccd1 _0586_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout577 _0809_/B vssd1 vssd1 vccd1 vccd1 _0839_/B sky130_fd_sc_hd__clkbuf_4
Xfanout588 _0773_/Y vssd1 vssd1 vccd1 vccd1 _0880_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_359_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_324_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_282_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_285_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_318_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0953_ hold257/X _0953_/A2 _0952_/X vssd1 vssd1 vccd1 vccd1 _0953_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0884_ hold280/X _0880_/A _0883_/X vssd1 vssd1 vccd1 vccd1 _0884_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_258_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0727__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_254_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_345_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_383_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold105_A _0505_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_310_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0718__B1 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_272_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_359_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 io_oeb_8x305[4] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
Xinput27 io_oeb_scrapcpu[18] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
Xinput38 io_oeb_scrapcpu[28] vssd1 vssd1 vccd1 vccd1 _0587_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_268_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput49 io_oeb_scrapcpu[5] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_1
XFILLER_0_220_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_295_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output446_A _0592_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1221_ _1221_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 _1221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_251_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1152_ _1187_/CLK _1152_/D vssd1 vssd1 vccd1 vccd1 _1152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_245_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1083_ _0852_/A _1084_/S hold637/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _1083_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_365_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_373_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold83_A hold83/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0936_ _1036_/A _0936_/B vssd1 vssd1 vccd1 vccd1 _0936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0867_ hold250/X hold729/A hold602/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0867_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0798_ hold267/X _0810_/A2 _0797_/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0798_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_286_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_254_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0651__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0875__C1 _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_387_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_347_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_347_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output396_A _1101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0721_ _0721_/A _0721_/B _0721_/C vssd1 vssd1 vccd1 vccd1 _0721_/X sky130_fd_sc_hd__or3_4
Xhold608 hold773/X vssd1 vssd1 vccd1 vccd1 _1050_/A sky130_fd_sc_hd__buf_1
XANTENNA_output563_A hold297/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0652_ _0652_/A1 _0660_/A2 _0696_/B1 _0652_/B2 vssd1 vssd1 vccd1 vccd1 _0653_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_268_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold619 _1005_/Y vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_268_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0583_ _0583_/A1 _0590_/A2 _0604_/A2 input36/X _0516_/B vssd1 vssd1 vccd1 vccd1 _0583_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_228_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _1204_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _1204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_251_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1135_ _1189_/CLK _1135_/D vssd1 vssd1 vccd1 vccd1 _1135_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_378_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1066_ _0956_/Y hold215/X _1065_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1066_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_149_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0919_ hold289/X _0952_/A2 _0952_/B1 _1038_/A _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0919_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_302_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_367_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout594_A _0515_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput217 io_out_as1802[27] vssd1 vssd1 vccd1 vccd1 _0715_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput206 io_out_as1802[17] vssd1 vssd1 vccd1 vccd1 _0675_/B2 sky130_fd_sc_hd__buf_2
Xinput228 io_out_as1802[4] vssd1 vssd1 vccd1 vccd1 _0623_/B2 sky130_fd_sc_hd__buf_2
Xinput239 io_out_scrapcpu[14] vssd1 vssd1 vccd1 vccd1 _0664_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_236_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_384_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold604_A _0851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_297_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0560__B2 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_379_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_387_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0615__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0704_ _0704_/A1 _0732_/A2 _0748_/B1 _0704_/B2 vssd1 vssd1 vccd1 vccd1 _0705_/C sky130_fd_sc_hd__a22o_1
Xhold405 hold790/X vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold416 hold791/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dlygate4sd3_1
X_0635_ _0635_/A1 _0514_/B _0695_/B1 _0635_/B2 vssd1 vssd1 vccd1 vccd1 _0637_/B sky130_fd_sc_hd__a22o_1
Xhold438 hold13/X vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_311_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0566_ input11/X _0593_/A hold95/X vssd1 vssd1 vccd1 vccd1 _0569_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_110_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1118_ _1221_/CLK _1118_/D vssd1 vssd1 vccd1 vccd1 _1118_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1049_ _1050_/C _1049_/B vssd1 vssd1 vccd1 vccd1 _1049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_319_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_302_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_255_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0533__A1 _0533_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0509__C _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0836__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_390_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_371_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold202 hold552/X vssd1 vssd1 vccd1 vccd1 _1156_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold235 _1109_/Q vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _0915_/Y vssd1 vssd1 vccd1 vccd1 _1141_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold213 hold680/X vssd1 vssd1 vccd1 vccd1 _1094_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_348_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold246 _0835_/X vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold384/X vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold268 hold663/X vssd1 vssd1 vccd1 vccd1 _1097_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0618_ _0618_/A1 _0674_/A2 _0674_/B1 _0618_/B2 vssd1 vssd1 vccd1 vccd1 _0621_/A sky130_fd_sc_hd__a22o_1
Xhold279 hold701/X vssd1 vssd1 vccd1 vccd1 _1115_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0549_ input21/X _0604_/A2 _0586_/B1 input57/X vssd1 vssd1 vccd1 vccd1 _0549_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_237_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_108 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_366_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_322_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold780 _1148_/Q vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_274_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0818__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_372_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_353_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output476_A _0705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_348_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout589 _0773_/Y vssd1 vssd1 vccd1 vccd1 _0953_/A2 sky130_fd_sc_hd__buf_4
Xfanout578 _0827_/B vssd1 vssd1 vccd1 vccd1 _0809_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_308_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0736__B2 _0736_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_19 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0952_ hold525/X _0952_/A2 _0952_/B1 hold322/X _0952_/C1 vssd1 vssd1 vccd1 vccd1
+ _0952_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0803__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0883_ hold265/X _0776_/A hold605/A _0999_/A _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0883_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_341_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0727__A1 _0727_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0727__B2 _0727_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_266_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0663__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0966__A1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0718__B2 _0718_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 io_oeb_as1802 vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_330_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput28 io_oeb_scrapcpu[19] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput39 io_oeb_scrapcpu[29] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
XFILLER_0_220_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output439_A _1254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1220_ _1221_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 _1220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1151_ _1154_/CLK _1151_/D vssd1 vssd1 vccd1 vccd1 _1151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_251_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1082_ _1082_/A _1082_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _1082_/X sky130_fd_sc_hd__or3_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_373_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0935_ hold179/X _0953_/A2 _0934_/X vssd1 vssd1 vccd1 vccd1 _0935_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0866_ _0880_/A _0866_/B vssd1 vssd1 vccd1 vccd1 _0866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0797_ _0797_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_254_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0581__C1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_388_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput490 _0617_/X vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_12
XFILLER_0_233_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0627__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_362_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0720_ _0720_/A1 _0732_/A2 _0748_/B1 _0720_/B2 vssd1 vssd1 vccd1 vccd1 _0721_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output389_A _0765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 _1041_/Y vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0651_ _0651_/A1 _0593_/A _0695_/B1 _0651_/B2 vssd1 vssd1 vccd1 vccd1 _0653_/B sky130_fd_sc_hd__a22o_1
XANTENNA_output556_A hold173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0582_ input71/X _0586_/B1 _0574_/X _0581_/X vssd1 vssd1 vccd1 vccd1 _1256_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_283_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_326_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_256_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1203_ _1204_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _1203_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1134_ _1157_/CLK _1134_/D vssd1 vssd1 vccd1 vccd1 _1134_/Q sky130_fd_sc_hd__dfxtp_1
X_1065_ _1065_/A _1076_/B vssd1 vssd1 vccd1 vccd1 _1065_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0918_ _1036_/A _0918_/B vssd1 vssd1 vccd1 vccd1 _0918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_367_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0849_ _0849_/A _0849_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _0849_/X sky130_fd_sc_hd__or3_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput218 io_out_as1802[28] vssd1 vssd1 vccd1 vccd1 _0719_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput207 io_out_as1802[18] vssd1 vssd1 vccd1 vccd1 _0679_/B2 sky130_fd_sc_hd__buf_2
Xinput229 io_out_as1802[5] vssd1 vssd1 vccd1 vccd1 _0627_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_215_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_384_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_384_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0560__A2 hold100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__buf_1
XFILLER_0_387_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_242_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0703_ _0703_/A1 _0747_/A2 _0515_/Y _0703_/B2 vssd1 vssd1 vccd1 vccd1 _0705_/B sky130_fd_sc_hd__a22o_1
Xhold406 hold802/X vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0811__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold417 hold3/X vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0634_ _0634_/A1 _0674_/A2 _0674_/B1 _0634_/B2 vssd1 vssd1 vccd1 vccd1 _0637_/A sky130_fd_sc_hd__a22o_1
XANTENNA__0784__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold428 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 hold439/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0565_ _0565_/A _0565_/B _0565_/C vssd1 vssd1 vccd1 vccd1 _1249_/A sky130_fd_sc_hd__or3_4
XFILLER_0_110_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_366_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1117_ _1221_/CLK _1117_/D vssd1 vssd1 vccd1 vccd1 _1117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1048_ _0821_/A _1080_/B hold593/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_381_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0705__C _0705_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0790__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_255_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_369_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_384_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold9_A hold9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0533__A2 _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output421_A _1095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_316_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold214 hold769/X vssd1 vssd1 vccd1 vccd1 _1071_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold203 hold389/X vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__clkbuf_2
Xhold225 _1119_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold247 hold524/X vssd1 vssd1 vccd1 vccd1 _1116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _0953_/Y vssd1 vssd1 vccd1 vccd1 _0954_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold654/X vssd1 vssd1 vccd1 vccd1 _1109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold388/X vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0617_ _0617_/A _0617_/B _0617_/C vssd1 vssd1 vccd1 vccd1 _0617_/X sky130_fd_sc_hd__or3_4
XFILLER_0_284_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_284_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0548_ input92/X _0605_/A2 _0565_/A _0547_/X vssd1 vssd1 vccd1 vccd1 _1242_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_364_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_109 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_380_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold781 _1147_/Q vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold770 _1172_/Q vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold792 _1149_/Q vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_389_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_360_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output469_A _0609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0690__B2 _0690_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_351_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_304_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout579 _0810_/A2 vssd1 vssd1 vccd1 vccd1 _0840_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_308_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_324_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_354_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_290_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1215_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0672__B2 _0672_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0951_ _1036_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_333_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0882_ _0882_/A _0882_/B _0882_/C vssd1 vssd1 vccd1 vccd1 _0882_/X sky130_fd_sc_hd__and3_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_341_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_329_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0663__B2 _0663_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0663__A1 _0663_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0718__A2 _0505_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_255_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_272_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0654__B2 _0654_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_382_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 io_oeb_scrapcpu[0] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 io_oeb_scrapcpu[1] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1150_ _1187_/CLK _1150_/D vssd1 vssd1 vccd1 vccd1 _1150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_359_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1081_ _0956_/Y _1078_/X hold323/X _1080_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1081_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__0893__A1 hold303/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_318_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_306_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0934_ hold527/X _0775_/A _0851_/X hold725/X _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0934_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0865_ hold339/X _0776_/A hold605/A hold600/A _0864_/X vssd1 vssd1 vccd1 vccd1 _0865_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_341_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0796_ hold166/X _0810_/A2 _0795_/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0796_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_48_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_254_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0884__A1 hold280/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0636__B2 _0636_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_364_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_309_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_320_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput480 _0613_/X vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
Xoutput491 _0621_/X vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
XFILLER_0_233_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0875__A1 hold272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0627__B2 _0627_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0627__A1 _0627_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_370_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0650_ _0650_/A1 _0674_/A2 _0674_/B1 _0650_/B2 vssd1 vssd1 vccd1 vccd1 _0653_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0581_ _0581_/A1 _0590_/A2 _0604_/A2 input35/X _0516_/B vssd1 vssd1 vccd1 vccd1 _0581_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_output549_A hold206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output451_A _1265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_283_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0563__B1 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_291_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1202_ _1204_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 _1202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0809__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_378_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1133_ _1157_/CLK _1133_/D vssd1 vssd1 vccd1 vccd1 _1133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1064_ _1071_/A _1071_/D vssd1 vssd1 vccd1 vccd1 _1064_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_393_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0618__B2 _0618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0917_ hold209/X _0953_/A2 _0916_/X vssd1 vssd1 vccd1 vccd1 _0917_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0848_ _0868_/A hold739/X hold369/X _0955_/B vssd1 vssd1 vccd1 vccd1 _0848_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_367_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0779_ _0779_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput208 io_out_as1802[19] vssd1 vssd1 vccd1 vccd1 _0683_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_383_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput219 io_out_as1802[29] vssd1 vssd1 vccd1 vccd1 _0723_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_215_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_337_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_357_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0848__A1 _0868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_373_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_242_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0702_ _0702_/A1 _0746_/A2 _0746_/B1 _0702_/B2 vssd1 vssd1 vccd1 vccd1 _0705_/A sky130_fd_sc_hd__a22o_1
Xhold407 hold801/X vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 hold418/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0633_ _0633_/A _0633_/B _0633_/C vssd1 vssd1 vccd1 vccd1 _0633_/X sky130_fd_sc_hd__or3_4
XFILLER_0_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold429 hold23/X vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_337_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0564_ input99/X _0605_/A2 _0510_/B input63/X vssd1 vssd1 vccd1 vccd1 _0565_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1116_ _1221_/CLK _1116_/D vssd1 vssd1 vccd1 vccd1 _1116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_366_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1047_ hold592/X _1049_/B _1076_/B vssd1 vssd1 vccd1 vccd1 _1047_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_381_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_381_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1154_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_262_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0766__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_348_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_363_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 _1064_/X vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _0941_/Y vssd1 vssd1 vccd1 vccd1 _0942_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_348_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold248 hold717/X vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 _0954_/Y vssd1 vssd1 vccd1 vccd1 _1154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 hold404/X vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0616_ _0616_/A1 _0660_/A2 _0628_/B1 _0616_/B2 vssd1 vssd1 vccd1 vccd1 _0617_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0547_ input20/X _0604_/A2 _0586_/B1 input56/X vssd1 vssd1 vccd1 vccd1 _0547_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_244_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_366_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout612_A _0775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_258_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold782 _1151_/Q vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 _0892_/X vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _1096_/Q vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 _1133_/Q vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_389_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_353_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0739__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_266_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput380 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _0768_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0817__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold99_A hold99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_308_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_284_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_340_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_340_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 _1169_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_263_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_381_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_385_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0950_ hold229/X _0953_/A2 _0949_/X vssd1 vssd1 vccd1 vccd1 _0950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output481_A _0721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0881_ hold316/X hold729/A hold569/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0881_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_301_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_301_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0663__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_289_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_332_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_386_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_359_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 io_oeb_scrapcpu[10] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0590__A1 _0590_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_263_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0878__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1080_ _1080_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1080_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0933_ _1036_/A _0933_/B vssd1 vssd1 vccd1 vccd1 _0933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1070__A2 _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0864_ hold99/A _1082_/C vssd1 vssd1 vccd1 vccd1 _0864_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0795_ _0795_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0795_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0581__A1 _0581_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_254_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_242_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1061__A2 _1181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_320_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0572__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput470 _0681_/X vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
Xoutput492 _0625_/X vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
Xoutput481 _0721_/X vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_12
XFILLER_0_245_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0627__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_370_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0580_ input70/X _0586_/B1 _0574_/X _0579_/X vssd1 vssd1 vccd1 vccd1 _1255_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output444_A _1232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0563__B2 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_291_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1201_ _1204_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _1201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1132_ _1157_/CLK _1132_/D vssd1 vssd1 vccd1 vccd1 _1132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1063_ _0829_/A _1076_/B hold533/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _1063_/X sky130_fd_sc_hd__o211a_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0825__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0916_ hold320/X _0952_/A2 _0952_/B1 _1032_/B _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0916_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0847_ _0847_/A _1082_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _0847_/X sky130_fd_sc_hd__or3_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0778_ hold346/X _0810_/A2 _0777_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0778_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_302_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0554__A1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput209 io_out_as1802[1] vssd1 vssd1 vccd1 vccd1 _0611_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_267_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1019__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0751__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0545__A1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0629__C _0629_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__buf_1
XFILLER_0_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_383_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_242_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output394_A _1099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0701_ _0701_/A _0701_/B _0701_/C vssd1 vssd1 vccd1 vccd1 _0701_/X sky130_fd_sc_hd__or3_4
XFILLER_0_154_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output561_A hold188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 hold799/X vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0632_ _0632_/A1 _0660_/A2 _0696_/B1 _0632_/B2 vssd1 vssd1 vccd1 vccd1 _0633_/C sky130_fd_sc_hd__a22o_2
XFILLER_0_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold419 hold747/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0563_ input27/X hold100/X _0518_/B input15/X vssd1 vssd1 vccd1 vccd1 _0565_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_249_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1115_ _1184_/CLK _1115_/D vssd1 vssd1 vccd1 vccd1 _1115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_283_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1046_ _1177_/Q _1050_/B _1050_/D vssd1 vssd1 vccd1 vccd1 _1049_/B sky130_fd_sc_hd__and3_1
XFILLER_0_393_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_381_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_334_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_334_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout592_A _0526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_270_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_288_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0766__A1 _1095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output407_A _1111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold216 hold697/X vssd1 vssd1 vccd1 vccd1 _1183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _0942_/Y vssd1 vssd1 vccd1 vccd1 _1150_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold249 hold718/X vssd1 vssd1 vccd1 vccd1 _1110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold238 _0902_/Y vssd1 vssd1 vccd1 vccd1 _0903_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _1099_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_296_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0615_ _0615_/A1 _0514_/B _0695_/B1 _0615_/B2 vssd1 vssd1 vccd1 vccd1 _0617_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0546_ input17/X _0516_/B hold95/A vssd1 vssd1 vccd1 vccd1 _0565_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_364_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_252_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_366_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1029_ _1032_/A _1033_/A vssd1 vssd1 vccd1 vccd1 _1029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_A hold100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0748__B2 _0748_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold750 _1072_/X vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _1184_/Q vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold761 _1171_/Q vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold783 _1146_/Q vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _1131_/Q vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0920__A1 hold232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_357_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_370_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_313_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0739__B2 _0739_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0739__A1 _0739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0911__A1 hold206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput381 hold741/X vssd1 vssd1 vccd1 vccd1 _0774_/A sky130_fd_sc_hd__clkbuf_1
Xinput370 hold438/X vssd1 vssd1 vccd1 vccd1 hold439/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0675__B1 _0683_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_280_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0833__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0529_ input12/X _0518_/B hold95/A vssd1 vssd1 vccd1 vccd1 _0529_/X sky130_fd_sc_hd__a21o_4
XANTENNA__0902__A1 hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_324_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_342_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold580 _1051_/Y vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 hold778/X vssd1 vssd1 vccd1 vccd1 _1050_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_263_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_377_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0637__C _0637_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0880_ _0880_/A _0880_/B vssd1 vssd1 vccd1 vccd1 _0880_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output474_A _0697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_361_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_324_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_289_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0639__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_342_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_392_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1055__B1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ hold182/X _0953_/A2 _0931_/X vssd1 vssd1 vccd1 vccd1 _0932_/Y sky130_fd_sc_hd__a21oi_1
X_0863_ hold297/X hold729/A hold690/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0863_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0794_ hold265/X _0810_/A2 _0793_/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0794_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_392_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_282_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_372_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_250_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput460 _0645_/X vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
Xoutput471 _0685_/X vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_285_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput493 _0629_/X vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
Xoutput482 _0725_/X vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_346_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0563__A2 hold100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output437_A _1252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1200_ _1204_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _1200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_256_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ _1157_/CLK _1131_/D vssd1 vssd1 vccd1 vccd1 _1131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1062_ _1071_/D hold532/X _1080_/B vssd1 vssd1 vccd1 vccd1 _1062_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_378_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_319_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0915_ _1036_/A _0915_/B vssd1 vssd1 vccd1 vccd1 _0915_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_259_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0846_ hold99/X hold739/X hold353/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0777_ _1082_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0777_/X sky130_fd_sc_hd__or2_1
XFILLER_0_302_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_388_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_316_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0751__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0778__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_375_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0645__C _0645_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_390_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ _0700_/A1 _0732_/A2 _0748_/B1 _0700_/B2 vssd1 vssd1 vccd1 vccd1 _0701_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_111_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output387_A _0761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold409 hold795/X vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0784__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0631_ _0631_/A1 _0514_/B _0695_/B1 _0631_/B2 vssd1 vssd1 vccd1 vccd1 _0633_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_296_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_296_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0562_ _0565_/A _0562_/B _0562_/C vssd1 vssd1 vccd1 vccd1 _1248_/A sky130_fd_sc_hd__or3_4
XFILLER_0_267_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1114_ _1184_/CLK _1114_/D vssd1 vssd1 vccd1 vccd1 _1114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1045_ _1050_/B _1045_/B vssd1 vssd1 vccd1 vccd1 _1045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0829_ _0829_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0829_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout585_A _0505_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_270_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_372_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_363_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold217 hold390/X vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__clkbuf_2
Xhold206 hold393/X vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0614_ _0614_/A1 _0674_/A2 _0674_/B1 _0614_/B2 vssd1 vssd1 vccd1 vccd1 _0617_/A sky130_fd_sc_hd__a22o_1
Xhold239 _0903_/Y vssd1 vssd1 vccd1 vccd1 _1137_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold228 hold671/X vssd1 vssd1 vccd1 vccd1 _1099_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_278_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0545_ input91/X _0605_/A2 _0529_/X _0544_/X vssd1 vssd1 vccd1 vccd1 _1241_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_147_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1028_ _1032_/A _1037_/B _1037_/C vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__and3_1
XFILLER_0_366_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 _1186_/Q vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _1177_/Q vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 _1194_/Q vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold784 _1150_/Q vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 _1127_/Q vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0757__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_389_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0684__B2 _0684_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput371 hold516/X vssd1 vssd1 vccd1 vccd1 hold517/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput360 hold480/X vssd1 vssd1 vccd1 vccd1 hold481/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_395_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_264_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0675__A1 _0675_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0675__B2 _0675_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_318_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_359_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0528_ _0528_/A1 _0506_/B _0526_/X _0527_/X vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_379_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0666__B2 _0666_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold581 _1052_/X vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 hold770/X vssd1 vssd1 vccd1 vccd1 _1024_/A sky130_fd_sc_hd__buf_1
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold592 _1045_/Y vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_365_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_318_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0653__C _0653_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output467_A _0673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0896__A1 hold254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput190 io_out_8x305[35] vssd1 vssd1 vccd1 vccd1 _0746_/B2 sky130_fd_sc_hd__buf_2
XANTENNA__0648__B2 _0648_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_376_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0860__A _0860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_332_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_260_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0887__A1 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0639__B2 _0639_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0639__A1 _0639_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_367_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_291_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_248_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_263_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0878__A1 hold310/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_358_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ hold314/X _0952_/A2 _0952_/B1 _1060_/A _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0931_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0862_ _0880_/A _0862_/B vssd1 vssd1 vccd1 vccd1 _0862_/X sky130_fd_sc_hd__or2_1
XFILLER_0_314_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0793_ _0793_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0793_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0566__B1 hold95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_385_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0839__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_364_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1224_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_320_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0557__B1 _0518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_292_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput461 _0649_/X vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
Xoutput450 _0601_/X vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_0_245_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput494 _0633_/X vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
Xoutput472 _0689_/X vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
Xoutput483 _0729_/X vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_12
XFILLER_0_346_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0765__A _0767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1130_ _1157_/CLK _1130_/D vssd1 vssd1 vccd1 vccd1 _1130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_256_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_252_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1061_ _1060_/A _1181_/Q _1060_/D _1060_/C vssd1 vssd1 vccd1 vccd1 _1061_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_393_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_300_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0914_ hold222/X _0953_/A2 _0913_/X vssd1 vssd1 vccd1 vccd1 _0914_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0845_ _0845_/A _0849_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _0845_/X sky130_fd_sc_hd__or3_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_314_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0776_ _0776_/A _1082_/B vssd1 vssd1 vccd1 vccd1 _0827_/B sky130_fd_sc_hd__or2_1
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0711__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1259_ hold78/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_375_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_375_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_383_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0661__C _0661_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0630_ _0630_/A1 _0674_/A2 _0674_/B1 _0630_/B2 vssd1 vssd1 vccd1 vccd1 _0633_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0561_ input98/X _0605_/A2 _0510_/B input62/X vssd1 vssd1 vccd1 vccd1 _0562_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_249_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1113_ _1221_/CLK _1113_/D vssd1 vssd1 vccd1 vccd1 _1113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_378_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1044_ _0819_/A _1080_/B hold610/X _0955_/B vssd1 vssd1 vccd1 vccd1 _1044_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_393_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0852__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0828_ hold527/X _0840_/A2 hold169/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0828_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_302_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0759_ _0767_/A _0767_/B _0759_/C vssd1 vssd1 vccd1 vccd1 _0759_/X sky130_fd_sc_hd__and3_4
XFILLER_0_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_270_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_270_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_357_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_375_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold207 _0911_/Y vssd1 vssd1 vccd1 vccd1 _0912_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_296_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0613_ _0613_/A _0613_/B _0613_/C vssd1 vssd1 vccd1 vccd1 _0613_/X sky130_fd_sc_hd__or3_4
Xhold218 _0947_/Y vssd1 vssd1 vccd1 vccd1 _0948_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold394/X vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0544_ input19/X _0598_/A2 _0586_/B1 input55/X vssd1 vssd1 vccd1 vccd1 _0544_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_294_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_339_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ _0811_/A _1080_/B hold545/X _0955_/B vssd1 vssd1 vccd1 vccd1 _1027_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold730 _0871_/X vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold752 _1075_/X vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 wbs_we_i vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _1097_/Q vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold796 _1138_/Q vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _1132_/Q vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold774 _1166_/Q vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_290_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0757__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_313_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_274_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1187_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_234_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput372 hold504/X vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__clkbuf_1
Xinput350 hold441/X vssd1 vssd1 vccd1 vccd1 hold442/A sky130_fd_sc_hd__buf_1
Xinput361 hold492/X vssd1 vssd1 vccd1 vccd1 hold493/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_264_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0675__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_280_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_272_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0527_ input40/X _0598_/A2 _0586_/B1 input76/X vssd1 vssd1 vccd1 vccd1 _0527_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_339_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0593__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold571 _1020_/Y vssd1 vssd1 vccd1 vccd1 _1021_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _0981_/X vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_263_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold593 _1047_/Y vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 hold758/X vssd1 vssd1 vccd1 vccd1 _1016_/C sky130_fd_sc_hd__buf_1
XFILLER_0_256_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_381_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_326_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_254_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput180 io_out_8x305[26] vssd1 vssd1 vccd1 vccd1 _0710_/B2 sky130_fd_sc_hd__buf_2
Xinput191 io_out_8x305[3] vssd1 vssd1 vccd1 vccd1 _0618_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_291_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0820__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0860__B _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0639__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0575__A1 _0575_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold390 hold756/X vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_263_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_244_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ _1036_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0861_ hold337/X _0776_/A hold605/A _0967_/C _0860_/X vssd1 vssd1 vccd1 vccd1 _0862_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0802__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0792_ hold212/X _0810_/A2 _0791_/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0792_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_279_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0566__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_378_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0557__B2 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput462 _0653_/X vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
Xoutput440 _1255_/A vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__buf_12
Xoutput451 _1265_/A vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__buf_12
XFILLER_0_285_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_245_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput495 _0637_/X vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
Xoutput473 _0693_/X vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
Xoutput484 _0733_/X vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_12
XFILLER_0_346_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0765__B _0767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_362_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_362_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0548__A1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0720__B2 _0720_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1060_ _1060_/A _1181_/Q _1060_/C _1060_/D vssd1 vssd1 vccd1 vccd1 _1071_/D sky130_fd_sc_hd__and4_2
XFILLER_0_393_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0913_ hold274/X _0952_/A2 _0952_/B1 _1032_/A _0934_/C1 vssd1 vssd1 vccd1 vccd1 _0913_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0844_ _0860_/A hold739/X hold349/X _0966_/C1 vssd1 vssd1 vccd1 vccd1 _0844_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0539__A1 _0539_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0775_ _0775_/A _1082_/B vssd1 vssd1 vccd1 vccd1 _0775_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0711__B2 _0711_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0711__A1 _0711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1258_ _1258_/A vssd1 vssd1 vccd1 vccd1 _1258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_250_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1189_ _1189_/CLK _1189_/D vssd1 vssd1 vccd1 vccd1 _1189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_377_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0950__A1 hold229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0702__B2 _0702_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0560_ input26/X hold100/X _0518_/B input14/X vssd1 vssd1 vccd1 vccd1 _0562_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output442_A _1257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0941__A1 hold203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1112_ _1221_/CLK _1112_/D vssd1 vssd1 vccd1 vccd1 _1112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1043_ hold609/X _1045_/B _1080_/B vssd1 vssd1 vccd1 vccd1 _1043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_378_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_287_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ _1058_/A _0827_/B vssd1 vssd1 vccd1 vccd1 _0827_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0758_ input5/X _1091_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0759_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_394_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0689_ _0689_/A _0689_/B _0689_/C vssd1 vssd1 vccd1 vccd1 _0689_/X sky130_fd_sc_hd__or3_4
XANTENNA__0932__A1 hold182/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_369_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_368_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_261_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0687__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output392_A _1097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0611__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 _0912_/Y vssd1 vssd1 vccd1 vccd1 _1140_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0612_ _0612_/A1 _0660_/A2 _0628_/B1 _0612_/B2 vssd1 vssd1 vccd1 vccd1 _0613_/C sky130_fd_sc_hd__a22o_2
Xhold219 _0948_/Y vssd1 vssd1 vccd1 vccd1 _1152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_278_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0543_ _0543_/A1 _0605_/A2 _0529_/X _0542_/X vssd1 vssd1 vccd1 vccd1 _1240_/A sky130_fd_sc_hd__a211o_4
XANTENNA__0914__A1 hold222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0847__C _1082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1026_ hold544/X _1033_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1026_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_354_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0602__B1 _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold720 _0788_/X vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold764 _1153_/Q vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _0849_/B vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _1126_/Q vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _1195_/Q vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_275_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout590_A _0526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 _1145_/Q vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _1137_/Q vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 _1098_/Q vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_338_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_357_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_278_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput340 io_out_z80[8] vssd1 vssd1 vccd1 vccd1 _0638_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput362 hold501/X vssd1 vssd1 vccd1 vccd1 hold502/A sky130_fd_sc_hd__clkbuf_1
Xinput351 hold450/X vssd1 vssd1 vccd1 vccd1 hold451/A sky130_fd_sc_hd__buf_1
XFILLER_0_264_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_12
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_12
Xinput373 hold426/X vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_371_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0526_ _0526_/A hold95/A vssd1 vssd1 vccd1 vccd1 _0526_/X sky130_fd_sc_hd__or2_1
XFILLER_0_265_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_394_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1009_ hold587/X _1012_/B _1021_/A vssd1 vssd1 vccd1 vccd1 _1009_/Y sky130_fd_sc_hd__o21ai_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout603_A _0510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold572 _1021_/Y vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _1002_/X vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _1163_/Q vssd1 vssd1 vccd1 vccd1 _0983_/D sky130_fd_sc_hd__buf_1
Xhold594 _1048_/X vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _1012_/Y vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold648_A _0518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_318_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_360_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput181 io_out_8x305[27] vssd1 vssd1 vccd1 vccd1 _0714_/B2 sky130_fd_sc_hd__buf_2
Xinput170 io_out_8x305[17] vssd1 vssd1 vccd1 vccd1 _0674_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_262_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_262_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput192 io_out_8x305[4] vssd1 vssd1 vccd1 vccd1 _0622_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_376_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0509_ hold99/A hold86/X _0767_/A vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__and3_1
XFILLER_0_213_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_382_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_350_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold380 hold779/X vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold391 hold731/X vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_244_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0860_ _0860_/A _1082_/C vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output472_A _0689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0791_ _0791_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0791_/X sky130_fd_sc_hd__or2_1
XFILLER_0_314_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0566__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_364_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0989_ hold613/X _0992_/B _0996_/A vssd1 vssd1 vccd1 vccd1 _0989_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_332_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0557__A2 hold100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput430 _1246_/A vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput441 _1256_/A vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__buf_12
Xoutput452 _1266_/A vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_0_245_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput496 _1239_/X vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_12
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput463 _0657_/X vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
Xoutput474 _0697_/X vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
Xoutput485 _0737_/X vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__buf_12
XFILLER_0_245_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_387_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_395_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0781__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0796__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0972__A _0996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0912_ _1036_/A _0912_/B vssd1 vssd1 vccd1 vccd1 _0912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0843_ _0965_/A _0849_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _0843_/X sky130_fd_sc_hd__or3_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0774_ _0774_/A _0774_/B vssd1 vssd1 vccd1 vccd1 _0849_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_390_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0711__A2 _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1257_ _1257_/A vssd1 vssd1 vccd1 vccd1 _1257_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_384_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1188_ _1188_/CLK _1188_/D vssd1 vssd1 vccd1 vccd1 _1188_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0778__A2 _0810_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_375_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_383_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_311_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output435_A _1250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_362_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1111_ _1184_/CLK _1111_/D vssd1 vssd1 vccd1 vccd1 _1111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_366_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1042_ _1050_/A _1050_/D vssd1 vssd1 vccd1 vccd1 _1045_/B sky130_fd_sc_hd__and2_1
XFILLER_0_378_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0826_ hold314/X _0840_/A2 _0825_/X _0500_/Y vssd1 vssd1 vccd1 vccd1 _0826_/X sky130_fd_sc_hd__o211a_1
X_0757_ _0767_/A _0767_/B _0757_/C vssd1 vssd1 vccd1 vccd1 _0757_/X sky130_fd_sc_hd__and3_4
XFILLER_0_302_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0688_ _0688_/A1 _0732_/A2 _0696_/B1 _0688_/B2 vssd1 vssd1 vccd1 vccd1 _0689_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0696__B2 _0696_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_369_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_380_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0620__B2 _0620_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_368_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0687__B2 _0687_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0687__A1 _0687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output385_A _0757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0611__B2 _0611_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0611__A1 _0611_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0611_ _0611_/A1 _0514_/B _0695_/B1 _0611_/B2 vssd1 vssd1 vccd1 vccd1 _0613_/B sky130_fd_sc_hd__a22o_1
Xhold209 hold400/X vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output552_A hold220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0542_ input53/X _0598_/A2 _0598_/B1 input89/X vssd1 vssd1 vccd1 vccd1 _0542_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0678__B2 _0678_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_339_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1025_ _1037_/B _1037_/C vssd1 vssd1 vccd1 vccd1 _1033_/A sky130_fd_sc_hd__and2_1
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_362_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0850__A1 hold116/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_362_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0602__A1 input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold710 _0830_/X vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _1175_/Q vssd1 vssd1 vccd1 vccd1 _1032_/B sky130_fd_sc_hd__dlygate4sd3_1
X_0809_ _0809_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0809_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 _1123_/Q vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _0977_/X vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold743 _1193_/Q vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold765 _1180_/Q vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _1134_/Q vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 _1168_/Q vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_290_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold798 _1142_/Q vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput330 io_out_z80[31] vssd1 vssd1 vccd1 vccd1 _0730_/A1 sky130_fd_sc_hd__buf_1
Xinput341 io_out_z80[9] vssd1 vssd1 vccd1 vccd1 _0642_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput363 hold489/X vssd1 vssd1 vccd1 vccd1 hold490/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput352 hold432/X vssd1 vssd1 vccd1 vccd1 hold433/A sky130_fd_sc_hd__buf_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__clkbuf_2
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__clkbuf_4
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput374 hold459/X vssd1 vssd1 vccd1 vccd1 hold460/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_388_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_344_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0525_ _0525_/A1 _0506_/B hold95/X _0524_/X vssd1 vssd1 vccd1 vccd1 _1232_/A sky130_fd_sc_hd__a211o_4
XANTENNA__0899__A1 hold240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_394_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_394_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1008_ _1168_/Q _1016_/B _1008_/C vssd1 vssd1 vccd1 vccd1 _1012_/B sky130_fd_sc_hd__and3_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold540 _1038_/X vssd1 vssd1 vccd1 vccd1 _1039_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _0982_/Y vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold551 hold636/X vssd1 vssd1 vccd1 vccd1 _1082_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_275_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold573 _1022_/X vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _1013_/Y vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold761/X vssd1 vssd1 vccd1 vccd1 _1016_/D sky130_fd_sc_hd__buf_1
XFILLER_0_290_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0750__A0 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput171 io_out_8x305[18] vssd1 vssd1 vccd1 vccd1 _0678_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_268_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output515_A _1257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput160 io_out_6502[8] vssd1 vssd1 vccd1 vccd1 _0639_/A1 sky130_fd_sc_hd__buf_2
Xinput182 io_out_8x305[28] vssd1 vssd1 vccd1 vccd1 _0718_/B2 sky130_fd_sc_hd__buf_2
Xinput193 io_out_8x305[5] vssd1 vssd1 vccd1 vccd1 _0626_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_376_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_300_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0508_ _0518_/A _0508_/B vssd1 vssd1 vccd1 vccd1 _0508_/X sky130_fd_sc_hd__and2_2
XFILLER_0_272_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0885__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0779__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold381 hold780/X vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _0848_/X vssd1 vssd1 vccd1 vccd1 _1121_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0980__B1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold392 hold732/X vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_376_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_392_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_358_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_358_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_326_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0790_ hold331/X _0810_/A2 _0789_/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0790_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output465_A _0665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0723__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0988_ _0999_/A _1017_/A _1017_/B vssd1 vssd1 vccd1 vccd1 _0992_/B sky130_fd_sc_hd__and3_1
XFILLER_0_332_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput420 _1094_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[7] sky130_fd_sc_hd__buf_12
XFILLER_0_131_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0962__B1 _0956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput453 _1233_/A vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput431 _1247_/A vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput442 _1257_/A vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_0_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput464 _0661_/X vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
Xoutput475 _0701_/X vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_12
Xoutput486 _0741_/X vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__buf_12
XFILLER_0_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput497 _1240_/X vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_260_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_362_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_395_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_308_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_291_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0911_ hold206/X _0953_/A2 _0910_/X vssd1 vssd1 vccd1 vccd1 _0911_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0842_ _1082_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _1084_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_314_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0773_ _0882_/A _0882_/B vssd1 vssd1 vccd1 vccd1 _0773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_242_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_369_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1256_ _1256_/A vssd1 vssd1 vccd1 vccd1 _1256_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_250_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1187_ _1187_/CLK _1187_/D vssd1 vssd1 vccd1 vccd1 _1187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_250_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_392_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_357_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1234__A _1234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_387_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0871__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_383_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1110_ _1184_/CLK _1110_/D vssd1 vssd1 vccd1 vccd1 _1110_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output428_A _1244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1041_ _1050_/A _1050_/D vssd1 vssd1 vccd1 vccd1 _1041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1204_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_232_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_374_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0825_ _0825_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0825_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0756_ input4/X _1090_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0757_/C sky130_fd_sc_hd__mux2_1
X_0687_ _0687_/A1 _0747_/A2 _0695_/B1 _0687_/B2 vssd1 vssd1 vccd1 vccd1 _0689_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_255_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1239_ _1239_/A vssd1 vssd1 vccd1 vccd1 _1239_/X sky130_fd_sc_hd__buf_1
XFILLER_0_343_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_333_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_246_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0787__B _0839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_384_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_375_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0844__C1 _0966_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0611__A2 _0514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0610_ _0610_/A1 _0674_/A2 _0674_/B1 _0610_/B2 vssd1 vssd1 vccd1 vccd1 _0613_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_284_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0541_ _0541_/A1 _0605_/A2 _0529_/X _0540_/X vssd1 vssd1 vccd1 vccd1 _1239_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output545_A hold240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_294_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1024_ _1024_/A _1024_/B vssd1 vssd1 vccd1 vccd1 _1037_/C sky130_fd_sc_hd__and2_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_347_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_362_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_362_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold700 _1218_/Q vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
X_0808_ hold329/X _0810_/A2 _0807_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0808_/X sky130_fd_sc_hd__o211a_1
Xhold711 _1207_/Q vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold755 _1176_/Q vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 _1125_/Q vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0888__A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 hold740/X vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _1191_/Q vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
X_0739_ _0739_/A1 _0747_/A2 _0516_/B _0739_/B2 vssd1 vssd1 vccd1 vccd1 _0741_/B sky130_fd_sc_hd__a22o_1
Xhold788 _1140_/Q vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 _1188_/Q vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _1165_/Q vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold799 _1141_/Q vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_283_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_338_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0826__C1 _0500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_370_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_395_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_274_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput320 io_out_z80[22] vssd1 vssd1 vccd1 vccd1 _0694_/A1 sky130_fd_sc_hd__buf_1
Xinput331 io_out_z80[32] vssd1 vssd1 vccd1 vccd1 _0734_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput342 wb_rst_i vssd1 vssd1 vccd1 vccd1 input342/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput353 hold447/X vssd1 vssd1 vccd1 vccd1 hold448/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__buf_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput364 hold498/X vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__clkbuf_1
Xinput375 hold456/X vssd1 vssd1 vccd1 vccd1 hold457/A sky130_fd_sc_hd__clkbuf_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_329_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0832__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output495_A _0637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0596__A1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_2 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_257_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0524_ input29/X _0598_/A2 _0586_/B1 input65/X vssd1 vssd1 vccd1 vccd1 _0524_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_280_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_324_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_394_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_339_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0808__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1007_ _1016_/B _1007_/B vssd1 vssd1 vccd1 vccd1 _1007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_394_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold530 _0838_/X vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_275_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold541 _1039_/Y vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _0959_/X vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _0985_/Y vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 hold746/X vssd1 vssd1 vccd1 vccd1 _1032_/A sky130_fd_sc_hd__buf_1
Xhold596 _1015_/Y vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _1014_/X vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_365_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_283_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1242__A _1242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0814__A2 _0840_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_239_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_275_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput172 io_out_8x305[19] vssd1 vssd1 vccd1 vccd1 _0682_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_262_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput150 io_out_6502[31] vssd1 vssd1 vccd1 vccd1 _0731_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput161 io_out_6502[9] vssd1 vssd1 vccd1 vccd1 _0643_/A1 sky130_fd_sc_hd__buf_2
Xinput183 io_out_8x305[29] vssd1 vssd1 vccd1 vccd1 _0722_/B2 sky130_fd_sc_hd__buf_2
Xinput194 io_out_8x305[6] vssd1 vssd1 vccd1 vccd1 _0630_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0507_ hold99/X _0517_/B _0767_/A vssd1 vssd1 vccd1 vccd1 _0507_/X sky130_fd_sc_hd__and3_2
XFILLER_0_265_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1189_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_331_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1237__A _1237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 hold766/X vssd1 vssd1 vccd1 vccd1 _0852_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold360 hold373/X vssd1 vssd1 vccd1 vccd1 _0779_/A sky130_fd_sc_hd__buf_1
XFILLER_0_376_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold393 hold788/X vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 hold737/X vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0732__B2 _0732_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0795__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0689__C _0689_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output458_A _1238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0723__A1 _0723_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0723__B2 _0723_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_389_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0987_ _0999_/A _0987_/B vssd1 vssd1 vccd1 vccd1 _0987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_313_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput410 _1114_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[27] sky130_fd_sc_hd__buf_12
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput421 _1095_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[8] sky130_fd_sc_hd__buf_12
XANTENNA__1057__A _1181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput432 _1248_/A vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__buf_12
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput443 _1258_/A vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_0_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput454 _1234_/A vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__buf_12
Xoutput465 _0665_/X vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
Xoutput476 _0705_/X vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_12
Xoutput487 _0745_/X vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__buf_12
XANTENNA__0714__B2 _0714_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput498 _1241_/X vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_226_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_311_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_276_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0953__A1 hold257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold190 _0945_/Y vssd1 vssd1 vccd1 vccd1 _1151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_244_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0910_ hold299/X _0952_/A2 _0952_/B1 _1024_/B _0952_/C1 vssd1 vssd1 vccd1 vccd1 _0910_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_299_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0841_ _0851_/A _0841_/B hold738/X vssd1 vssd1 vccd1 vccd1 _0882_/C sky130_fd_sc_hd__or3b_2
XFILLER_0_314_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ _0772_/A _0882_/B vssd1 vssd1 vccd1 vccd1 _0772_/X sky130_fd_sc_hd__and2_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0944__A1 hold188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_369_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1255_ _1255_/A vssd1 vssd1 vccd1 vccd1 _1255_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_384_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1186_ _1187_/CLK _1186_/D vssd1 vssd1 vccd1 vccd1 _1186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_377_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_301_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0699__B1 _0515_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_387_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_373_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_242_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1250__A _1250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0623__B1 _0695_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_311_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0926__A1 hold269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1040_ _0817_/A _1080_/B hold541/X _0955_/B vssd1 vssd1 vccd1 vccd1 _1040_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0504__A hold76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0824_ hold248/X _0840_/A2 _0823_/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0824_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0755_ _0767_/A _0767_/B _0755_/C vssd1 vssd1 vccd1 vccd1 _0755_/X sky130_fd_sc_hd__and3_4
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0686_ _0686_/A1 _0746_/A2 _0746_/B1 _0686_/B2 vssd1 vssd1 vccd1 vccd1 _0689_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1238_ _1238_/A vssd1 vssd1 vccd1 vccd1 _1238_/X sky130_fd_sc_hd__buf_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1169_ _1205_/CLK _1169_/D vssd1 vssd1 vccd1 vccd1 _1169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A _1085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0908__A1 hold197/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_368_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1245__A _1245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_384_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_388_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_261_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_390_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_383_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_312_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0540_ input52/X _0598_/A2 _0598_/B1 input88/X vssd1 vssd1 vccd1 vccd1 _0540_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output440_A _1255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output538_A _0510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0697__C _0697_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0780__C1 _1083_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1023_ _1172_/Q _1037_/B _1024_/B vssd1 vssd1 vccd1 vccd1 _1023_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_366_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_339_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_362_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_362_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold701 _0834_/X vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 _0812_/X vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
X_0807_ _0807_/A _0809_/B vssd1 vssd1 vccd1 vccd1 _0807_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0738_ _0738_/A1 _0746_/A2 _0746_/B1 _0738_/B2 vssd1 vssd1 vccd1 vccd1 _0741_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold734 _1128_/Q vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _1155_/Q vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold723 hold768/X vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_268_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold756 _1152_/Q vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _1178_/Q vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold767 _1164_/Q vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
X_0669_ _0669_/A _0669_/B _0669_/C vssd1 vssd1 vccd1 vccd1 _0669_/X sky130_fd_sc_hd__or3_4
Xhold789 _1154_/Q vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_283_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_243_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_372_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_380_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_395_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput321 io_out_z80[23] vssd1 vssd1 vccd1 vccd1 _0698_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_219_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput310 io_out_z80[13] vssd1 vssd1 vccd1 vccd1 _0658_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput332 io_out_z80[33] vssd1 vssd1 vccd1 vccd1 _0738_/A1 sky130_fd_sc_hd__buf_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput343 hold423/X vssd1 vssd1 vccd1 vccd1 hold424/A sky130_fd_sc_hd__clkbuf_1
Xinput354 hold462/X vssd1 vssd1 vccd1 vccd1 hold463/A sky130_fd_sc_hd__buf_1
XFILLER_0_199_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput365 hold483/X vssd1 vssd1 vccd1 vccd1 hold484/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput376 hold486/X vssd1 vssd1 vccd1 vccd1 hold487/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_388_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_348_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_325_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output390_A _0767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output488_A _0749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_289_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_312_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0523_ input54/X hold82/X _0522_/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__a21o_4
XFILLER_0_158_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_394_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1006_ _0801_/A _1021_/A hold619/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_394_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold520 hold520/A vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_349_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold553 hold772/X vssd1 vssd1 vccd1 vccd1 _1071_/B sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold531 _1182_/Q vssd1 vssd1 vccd1 vccd1 _1060_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _1040_/X vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold575 _1029_/Y vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _1018_/Y vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 hold757/X vssd1 vssd1 vccd1 vccd1 _1016_/B sky130_fd_sc_hd__buf_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold564 _0986_/X vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_256_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_283_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_262_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput162 io_out_8x305[0] vssd1 vssd1 vccd1 vccd1 _0606_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput151 io_out_6502[32] vssd1 vssd1 vccd1 vccd1 _0735_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput140 io_out_6502[22] vssd1 vssd1 vccd1 vccd1 _0695_/A1 sky130_fd_sc_hd__buf_2
Xinput195 io_out_8x305[7] vssd1 vssd1 vccd1 vccd1 _0634_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput184 io_out_8x305[2] vssd1 vssd1 vccd1 vccd1 _0614_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput173 io_out_8x305[1] vssd1 vssd1 vccd1 vccd1 _0610_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_291_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_376_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_391_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_257_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0512__A hold76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_257_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_300_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0506_ _0518_/A _0506_/B vssd1 vssd1 vccd1 vccd1 _0506_/X sky130_fd_sc_hd__and2_1
XFILLER_0_185_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_265_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_367_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold350 _0844_/X vssd1 vssd1 vccd1 vccd1 _1119_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _0963_/X vssd1 vssd1 vccd1 vccd1 _1157_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_376_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold394 hold764/X vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold781/X vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold638/X vssd1 vssd1 vccd1 vccd1 _1188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_244_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1253__A _1253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_325_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_381_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_341_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_294_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_294_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_262_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_321_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0507__A hold99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0986_ _0791_/A _0996_/A hold563/X _1006_/C1 vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_320_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput411 _1115_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[28] sky130_fd_sc_hd__buf_12
Xoutput400 _1105_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[18] sky130_fd_sc_hd__buf_12
Xoutput422 _1096_/Q vssd1 vssd1 vccd1 vccd1 custom_settings[9] sky130_fd_sc_hd__buf_12
Xoutput433 hold83/A vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput444 _1232_/A vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__buf_12
Xoutput455 _1235_/A vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__buf_12
Xoutput466 _0669_/X vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput477 _0709_/X vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_12
XANTENNA__0714__A2 _0505_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput499 _1242_/X vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_12
Xoutput488 _0749_/X vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__buf_12
XFILLER_0_226_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_387_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1223__D hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_395_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold227_A _1099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0650__B2 _0650_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1248__A _1248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold180 _0935_/Y vssd1 vssd1 vccd1 vccd1 _0936_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold191 hold403/X vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold763_A _1097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_378_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ hold525/X _0840_/A2 hold295/X _1081_/C1 vssd1 vssd1 vccd1 vccd1 _0840_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_302_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0771_ hold412/X _0771_/B _0955_/A vssd1 vssd1 vccd1 vccd1 _0882_/B sky130_fd_sc_hd__and3b_1
XANTENNA_output568_A hold272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output470_A _0681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1254_ _1254_/A vssd1 vssd1 vccd1 vccd1 _1254_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_369_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1185_ _1187_/CLK _1185_/D vssd1 vssd1 vccd1 vccd1 _1185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_377_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_392_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0632__B2 _0632_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_360_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0969_ _1017_/A hold536/X _1021_/A vssd1 vssd1 vccd1 vccd1 _0969_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout599_A hold82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0699__A1 _0699_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0699__B2 _0699_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_242_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0871__A1 hold301/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0623__A1 _0623_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0623__B2 _0623_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_311_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_374_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_374_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_302_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0614__B2 _0614_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0823_ _0823_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0823_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0754_ input3/X _1089_/Q _1188_/Q vssd1 vssd1 vccd1 vccd1 _0755_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_295_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0685_ _0685_/A _0685_/B _0685_/C vssd1 vssd1 vccd1 vccd1 _0685_/X sky130_fd_sc_hd__or3_4
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0520__A hold99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_369_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1237_ _1237_/A vssd1 vssd1 vccd1 vccd1 _1237_/X sky130_fd_sc_hd__buf_1
XFILLER_0_211_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1168_ _1205_/CLK _1168_/D vssd1 vssd1 vccd1 vccd1 _1168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_377_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1099_ _1205_/CLK _1099_/D vssd1 vssd1 vccd1 vccd1 _1099_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_392_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0605__A1 _0605_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1261__A _1261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0844__A1 _0860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_356_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output433_A hold83/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1022_ _0809_/A _1021_/A hold572/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_359_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_374_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_362_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold702 _1111_/Q vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
X_0806_ hold306/X _0810_/A2 _0805_/X _1083_/C1 vssd1 vssd1 vccd1 vccd1 _0806_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0737_ _0737_/A _0737_/B _0737_/C vssd1 vssd1 vccd1 vccd1 _0737_/X sky130_fd_sc_hd__or3_4
Xhold746 _1174_/Q vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold713 _1210_/Q vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 _1130_/Q vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold724 hold753/X vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _1144_/Q vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 _1169_/Q vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold768 _1192_/Q vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
X_0668_ _0668_/A1 _0732_/A2 _0696_/B1 _0668_/B2 vssd1 vssd1 vccd1 vccd1 _0669_/C sky130_fd_sc_hd__a22o_1
XANTENNA__1065__B _1076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0599_ _0599_/A1 _0605_/A2 hold95/A _0598_/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__a211o_4
XANTENNA__0523__B1 _0522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_385_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_338_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_380_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_380_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_379_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_248_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1256__A _1256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_395_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_248_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0762__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput300 io_out_vliw[4] vssd1 vssd1 vccd1 vccd1 _0624_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput311 io_out_z80[14] vssd1 vssd1 vccd1 vccd1 _0662_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput333 io_out_z80[34] vssd1 vssd1 vccd1 vccd1 _0742_/A1 sky130_fd_sc_hd__buf_1
Xinput322 io_out_z80[24] vssd1 vssd1 vccd1 vccd1 _0702_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_117_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput344 hold420/X vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__clkbuf_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_388_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__buf_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput366 hold507/X vssd1 vssd1 vccd1 vccd1 hold508/A sky130_fd_sc_hd__clkbuf_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput377 hold495/X vssd1 vssd1 vccd1 vccd1 hold496/A sky130_fd_sc_hd__clkbuf_1
Xinput355 hold477/X vssd1 vssd1 vccd1 vccd1 hold478/A sky130_fd_sc_hd__buf_1
XFILLER_0_388_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__buf_2
XFILLER_0_199_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__buf_1
XFILLER_0_187_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_344_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output383_A _0753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output550_A hold222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_4 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0522_ input90/X _0506_/B _0598_/A2 input18/X hold95/A vssd1 vssd1 vccd1 vccd1 _0522_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_367_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_351_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1005_ hold618/X _1007_/B _1021_/A vssd1 vssd1 vccd1 vccd1 _1005_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_362_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_248_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold510 hold67/X vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold521 _1114_/Q vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _1068_/Y vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _1061_/Y vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _1173_/Q vssd1 vssd1 vccd1 vccd1 _1024_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold576 _1030_/Y vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 _1007_/Y vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/A vssd1 vssd1 vccd1 vccd1 _1163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_290_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout581_A _0506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 _1019_/X vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_365_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_385_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_338_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_341_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0735__B1 _0516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_275_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput163 io_out_8x305[10] vssd1 vssd1 vccd1 vccd1 _0646_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_262_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput152 io_out_6502[33] vssd1 vssd1 vccd1 vccd1 _0739_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput141 io_out_6502[23] vssd1 vssd1 vccd1 vccd1 _0699_/A1 sky130_fd_sc_hd__buf_2
Xinput130 io_out_6502[13] vssd1 vssd1 vccd1 vccd1 _0659_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_349_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput185 io_out_8x305[30] vssd1 vssd1 vccd1 vccd1 _0726_/B2 sky130_fd_sc_hd__buf_2
Xinput174 io_out_8x305[20] vssd1 vssd1 vccd1 vccd1 _0686_/B2 sky130_fd_sc_hd__buf_2
Xinput196 io_out_8x305[8] vssd1 vssd1 vccd1 vccd1 _0638_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_262_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_391_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0512__B hold99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0505_ _0505_/A hold77/X vssd1 vssd1 vccd1 vccd1 _0505_/Y sky130_fd_sc_hd__nor2_4
XANTENNA_hold33_A hold33/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
.ends

